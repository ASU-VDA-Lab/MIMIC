module fake_jpeg_77_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_61),
.Y(n_71)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_0),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_52),
.B1(n_48),
.B2(n_50),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_66),
.B1(n_56),
.B2(n_2),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_43),
.B1(n_52),
.B2(n_48),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_70),
.B1(n_3),
.B2(n_4),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_45),
.B1(n_42),
.B2(n_54),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_54),
.B1(n_45),
.B2(n_42),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_44),
.B(n_56),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_53),
.B1(n_51),
.B2(n_46),
.Y(n_70)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_78),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_44),
.B(n_2),
.C(n_3),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_4),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_82),
.Y(n_98)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_20),
.Y(n_93)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_22),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_24),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_5),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_74),
.B1(n_6),
.B2(n_7),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_104),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_40),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_10),
.C(n_11),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_111),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_26),
.B1(n_36),
.B2(n_35),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_16),
.B1(n_34),
.B2(n_33),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_114),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_116),
.B(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_8),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_9),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_90),
.B1(n_92),
.B2(n_95),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_118),
.B1(n_109),
.B2(n_111),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_100),
.B(n_89),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_133),
.C(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_9),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_124),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_134),
.B(n_137),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_139),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_123),
.C(n_132),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_112),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_143),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_127),
.C(n_126),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_122),
.B1(n_137),
.B2(n_129),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_141),
.C(n_11),
.Y(n_146)
);

OAI221xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.C(n_18),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

NOR2xp67_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_144),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_28),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_31),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_39),
.Y(n_153)
);


endmodule