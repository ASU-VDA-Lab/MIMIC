module fake_netlist_1_924_n_774 (n_117, n_44, n_133, n_149, n_81, n_69, n_204, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_96, n_39, n_774);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_204;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_96;
input n_39;
output n_774;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_383;
wire n_288;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_227;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_732;
wire n_752;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_580;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g209 ( .A(n_122), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_203), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_79), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_139), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_105), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_167), .Y(n_214) );
NOR2xp67_ASAP7_75t_L g215 ( .A(n_117), .B(n_164), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_155), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_84), .B(n_131), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_75), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_84), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_112), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_65), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_132), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_143), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_179), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_18), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_146), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_160), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_91), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_176), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_128), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_76), .Y(n_232) );
INVxp67_ASAP7_75t_L g233 ( .A(n_60), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_52), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_82), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_106), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_130), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_188), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_71), .Y(n_239) );
INVxp33_ASAP7_75t_SL g240 ( .A(n_37), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_180), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_173), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_142), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_88), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_140), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_24), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_73), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_89), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_78), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_96), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_16), .Y(n_251) );
INVxp33_ASAP7_75t_L g252 ( .A(n_25), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_202), .Y(n_253) );
INVxp33_ASAP7_75t_L g254 ( .A(n_104), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_147), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_172), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_64), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_152), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_108), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_178), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_2), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_61), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_17), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_70), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_177), .Y(n_265) );
INVxp67_ASAP7_75t_L g266 ( .A(n_208), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_175), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_121), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_77), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_26), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_97), .Y(n_271) );
INVxp33_ASAP7_75t_SL g272 ( .A(n_187), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_67), .Y(n_273) );
INVxp33_ASAP7_75t_L g274 ( .A(n_25), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_199), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_23), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_14), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_103), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_101), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_77), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_157), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_156), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_50), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_116), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_83), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_118), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_70), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_141), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_200), .Y(n_289) );
BUFx5_ASAP7_75t_L g290 ( .A(n_19), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_67), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_113), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_72), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_43), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_66), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_135), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_138), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_154), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_93), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_144), .Y(n_300) );
CKINVDCx14_ASAP7_75t_R g301 ( .A(n_86), .Y(n_301) );
INVxp67_ASAP7_75t_SL g302 ( .A(n_196), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_3), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_74), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_166), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_158), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_62), .Y(n_307) );
OA21x2_ASAP7_75t_L g308 ( .A1(n_212), .A2(n_0), .B(n_1), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_290), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_255), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_290), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_290), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_255), .Y(n_313) );
OA21x2_ASAP7_75t_L g314 ( .A1(n_212), .A2(n_2), .B(n_3), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_290), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_222), .A2(n_99), .B(n_98), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_237), .Y(n_317) );
AND2x6_ASAP7_75t_L g318 ( .A(n_241), .B(n_100), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_290), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_290), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_255), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_255), .Y(n_323) );
OAI22xp5_ASAP7_75t_SL g324 ( .A1(n_218), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_247), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_247), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_273), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_254), .B(n_7), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_254), .B(n_7), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_265), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_249), .B(n_8), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_252), .B(n_8), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_265), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_265), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_273), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_301), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_274), .B(n_9), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_265), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_301), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_274), .B(n_9), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_276), .B(n_10), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_240), .A2(n_13), .B1(n_11), .B2(n_12), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_241), .Y(n_343) );
INVx6_ASAP7_75t_L g344 ( .A(n_242), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_276), .B(n_13), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_278), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_323), .Y(n_347) );
INVx4_ASAP7_75t_L g348 ( .A(n_318), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_323), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_311), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_341), .A2(n_211), .B1(n_225), .B2(n_219), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_340), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_311), .B(n_245), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_323), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_317), .B(n_297), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_311), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_336), .Y(n_358) );
INVx6_ASAP7_75t_L g359 ( .A(n_318), .Y(n_359) );
INVx5_ASAP7_75t_L g360 ( .A(n_318), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_315), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_336), .B(n_271), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_341), .A2(n_232), .B1(n_235), .B2(n_234), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_315), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_315), .Y(n_365) );
AO21x2_ASAP7_75t_L g366 ( .A1(n_329), .A2(n_216), .B(n_210), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_319), .Y(n_367) );
NAND2xp33_ASAP7_75t_L g368 ( .A(n_318), .B(n_278), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_319), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_343), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_317), .B(n_266), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_339), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_319), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_319), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_341), .A2(n_239), .B1(n_246), .B2(n_244), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_341), .A2(n_248), .B1(n_251), .B2(n_250), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_366), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_353), .B(n_332), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_353), .A2(n_332), .B1(n_337), .B2(n_328), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_358), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_354), .Y(n_381) );
AND2x6_ASAP7_75t_L g382 ( .A(n_362), .B(n_345), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_370), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g384 ( .A(n_372), .B(n_345), .Y(n_384) );
BUFx5_ASAP7_75t_L g385 ( .A(n_370), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_370), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_366), .Y(n_387) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_351), .B(n_331), .C(n_342), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_348), .B(n_213), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_348), .B(n_243), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_348), .B(n_345), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_362), .Y(n_392) );
NOR2xp33_ASAP7_75t_SL g393 ( .A(n_348), .B(n_229), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_371), .B(n_345), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_372), .B(n_345), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_356), .B(n_331), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_348), .B(n_312), .Y(n_397) );
AND3x2_ASAP7_75t_SL g398 ( .A(n_363), .B(n_324), .C(n_221), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_375), .B(n_227), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_369), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_376), .A2(n_308), .B1(n_314), .B2(n_312), .Y(n_401) );
NAND2xp33_ASAP7_75t_L g402 ( .A(n_360), .B(n_318), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_366), .B(n_238), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_368), .A2(n_314), .B1(n_308), .B2(n_320), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_369), .B(n_209), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_360), .B(n_320), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_369), .B(n_296), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_373), .B(n_272), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_373), .B(n_326), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_350), .B(n_322), .Y(n_412) );
O2A1O1Ixp33_ASAP7_75t_L g413 ( .A1(n_368), .A2(n_233), .B(n_228), .C(n_309), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_359), .A2(n_314), .B1(n_308), .B2(n_322), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_381), .B(n_374), .Y(n_415) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_405), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_380), .B(n_306), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_397), .A2(n_357), .B(n_352), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_382), .B(n_374), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_382), .B(n_396), .Y(n_420) );
BUFx12f_ASAP7_75t_L g421 ( .A(n_382), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_400), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_391), .A2(n_364), .B(n_361), .Y(n_423) );
INVx5_ASAP7_75t_L g424 ( .A(n_382), .Y(n_424) );
NOR2xp67_ASAP7_75t_L g425 ( .A(n_388), .B(n_295), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g426 ( .A1(n_410), .A2(n_316), .B(n_309), .C(n_365), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_379), .B(n_299), .Y(n_427) );
OAI21x1_ASAP7_75t_L g428 ( .A1(n_414), .A2(n_316), .B(n_365), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_395), .B(n_367), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_414), .A2(n_316), .B(n_314), .Y(n_430) );
AOI22x1_ASAP7_75t_L g431 ( .A1(n_377), .A2(n_310), .B1(n_321), .B2(n_313), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_393), .B(n_214), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_384), .B(n_308), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_411), .Y(n_434) );
INVx4_ASAP7_75t_L g435 ( .A(n_385), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_383), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_403), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_394), .B(n_359), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_386), .Y(n_439) );
INVx5_ASAP7_75t_L g440 ( .A(n_405), .Y(n_440) );
O2A1O1Ixp5_ASAP7_75t_L g441 ( .A1(n_389), .A2(n_302), .B(n_217), .C(n_282), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_399), .Y(n_442) );
INVx8_ASAP7_75t_L g443 ( .A(n_405), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_412), .A2(n_387), .B(n_377), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_412), .A2(n_349), .B(n_347), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_390), .A2(n_261), .B(n_262), .C(n_257), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_406), .Y(n_447) );
O2A1O1Ixp5_ASAP7_75t_L g448 ( .A1(n_409), .A2(n_282), .B(n_292), .C(n_267), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_408), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_401), .A2(n_335), .B1(n_325), .B2(n_264), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_401), .A2(n_269), .B(n_270), .C(n_263), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_385), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_413), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_385), .B(n_280), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_398), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_405), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g457 ( .A1(n_404), .A2(n_307), .B(n_291), .Y(n_457) );
OAI21x1_ASAP7_75t_L g458 ( .A1(n_404), .A2(n_349), .B(n_347), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_402), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_407), .A2(n_285), .B(n_287), .C(n_283), .Y(n_460) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_405), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_381), .B(n_359), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_397), .A2(n_355), .B(n_223), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_397), .A2(n_355), .B(n_224), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_397), .A2(n_226), .B(n_220), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_381), .A2(n_335), .B1(n_325), .B2(n_293), .Y(n_466) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_405), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_400), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_405), .Y(n_469) );
AOI33xp33_ASAP7_75t_L g470 ( .A1(n_392), .A2(n_327), .A3(n_303), .B1(n_304), .B2(n_294), .B3(n_236), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_378), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_397), .A2(n_231), .B(n_230), .Y(n_472) );
AO31x2_ASAP7_75t_L g473 ( .A1(n_426), .A2(n_310), .A3(n_321), .B(n_313), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g474 ( .A1(n_451), .A2(n_256), .B(n_259), .C(n_258), .Y(n_474) );
AOI31xp67_ASAP7_75t_L g475 ( .A1(n_433), .A2(n_313), .A3(n_321), .B(n_310), .Y(n_475) );
OAI21x1_ASAP7_75t_L g476 ( .A1(n_458), .A2(n_292), .B(n_268), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_444), .A2(n_279), .B(n_275), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_430), .A2(n_284), .B(n_281), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_436), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_433), .A2(n_318), .B(n_289), .Y(n_480) );
AO31x2_ASAP7_75t_L g481 ( .A1(n_450), .A2(n_313), .A3(n_321), .B(n_310), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_439), .Y(n_482) );
NAND3xp33_ASAP7_75t_SL g483 ( .A(n_455), .B(n_300), .C(n_253), .Y(n_483) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_430), .A2(n_305), .B(n_298), .Y(n_484) );
OAI21x1_ASAP7_75t_L g485 ( .A1(n_428), .A2(n_215), .B(n_330), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g486 ( .A(n_424), .B(n_277), .Y(n_486) );
AOI21x1_ASAP7_75t_L g487 ( .A1(n_450), .A2(n_425), .B(n_432), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_448), .A2(n_318), .B(n_330), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_446), .A2(n_260), .B(n_288), .C(n_286), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_471), .Y(n_490) );
OAI21x1_ASAP7_75t_L g491 ( .A1(n_431), .A2(n_338), .B(n_334), .Y(n_491) );
INVx4_ASAP7_75t_L g492 ( .A(n_424), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_424), .B(n_15), .Y(n_493) );
OR2x6_ASAP7_75t_L g494 ( .A(n_421), .B(n_278), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_437), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_442), .A2(n_338), .B(n_334), .C(n_278), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_434), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_420), .A2(n_333), .B(n_323), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_453), .A2(n_333), .B(n_346), .C(n_323), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_447), .B(n_323), .Y(n_500) );
AO31x2_ASAP7_75t_L g501 ( .A1(n_466), .A2(n_346), .A3(n_333), .B(n_344), .Y(n_501) );
AO31x2_ASAP7_75t_L g502 ( .A1(n_460), .A2(n_346), .A3(n_333), .B(n_21), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_470), .B(n_20), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_441), .A2(n_346), .B(n_333), .C(n_22), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_438), .A2(n_346), .B(n_102), .Y(n_505) );
AO31x2_ASAP7_75t_L g506 ( .A1(n_435), .A2(n_29), .A3(n_27), .B(n_28), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_415), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_423), .A2(n_109), .B(n_107), .Y(n_508) );
INVx4_ASAP7_75t_L g509 ( .A(n_443), .Y(n_509) );
AO31x2_ASAP7_75t_L g510 ( .A1(n_435), .A2(n_32), .A3(n_30), .B(n_31), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_427), .B(n_33), .Y(n_511) );
AO21x1_ASAP7_75t_L g512 ( .A1(n_454), .A2(n_111), .B(n_110), .Y(n_512) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_416), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_422), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_418), .A2(n_115), .B(n_114), .Y(n_515) );
AO31x2_ASAP7_75t_L g516 ( .A1(n_452), .A2(n_36), .A3(n_34), .B(n_35), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_417), .Y(n_517) );
AO32x2_ASAP7_75t_L g518 ( .A1(n_457), .A2(n_38), .A3(n_39), .B1(n_40), .B2(n_41), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_449), .Y(n_519) );
OAI21x1_ASAP7_75t_L g520 ( .A1(n_445), .A2(n_120), .B(n_119), .Y(n_520) );
INVx5_ASAP7_75t_L g521 ( .A(n_443), .Y(n_521) );
AO31x2_ASAP7_75t_L g522 ( .A1(n_465), .A2(n_45), .A3(n_42), .B(n_44), .Y(n_522) );
AO31x2_ASAP7_75t_L g523 ( .A1(n_472), .A2(n_46), .A3(n_44), .B(n_45), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_462), .A2(n_124), .B(n_123), .Y(n_524) );
OAI21x1_ASAP7_75t_SL g525 ( .A1(n_429), .A2(n_46), .B(n_47), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_443), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_440), .B(n_48), .Y(n_527) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_419), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_468), .Y(n_529) );
AOI221xp5_ASAP7_75t_SL g530 ( .A1(n_463), .A2(n_49), .B1(n_51), .B2(n_53), .C(n_54), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_464), .Y(n_531) );
AO31x2_ASAP7_75t_L g532 ( .A1(n_459), .A2(n_56), .A3(n_53), .B(n_55), .Y(n_532) );
INVx8_ASAP7_75t_L g533 ( .A(n_416), .Y(n_533) );
CKINVDCx11_ASAP7_75t_R g534 ( .A(n_461), .Y(n_534) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_456), .A2(n_126), .B(n_125), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_461), .A2(n_129), .B(n_127), .Y(n_536) );
AO31x2_ASAP7_75t_L g537 ( .A1(n_461), .A2(n_57), .A3(n_58), .B(n_59), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_467), .A2(n_134), .B(n_133), .Y(n_538) );
INVx3_ASAP7_75t_L g539 ( .A(n_469), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_490), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_497), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_519), .B(n_63), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_503), .Y(n_543) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_534), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_478), .A2(n_65), .B(n_66), .Y(n_545) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_485), .A2(n_137), .B(n_136), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_514), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g548 ( .A(n_521), .B(n_68), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_493), .A2(n_69), .B1(n_71), .B2(n_73), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_499), .A2(n_80), .B(n_81), .Y(n_550) );
OAI21x1_ASAP7_75t_L g551 ( .A1(n_476), .A2(n_168), .B(n_207), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_529), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_479), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_482), .Y(n_554) );
AO31x2_ASAP7_75t_L g555 ( .A1(n_512), .A2(n_85), .A3(n_87), .B(n_88), .Y(n_555) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_505), .A2(n_171), .B(n_206), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_498), .A2(n_170), .B(n_205), .Y(n_557) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_491), .A2(n_169), .B(n_204), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_525), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_522), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_507), .B(n_90), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_522), .Y(n_562) );
INVx3_ASAP7_75t_L g563 ( .A(n_509), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_501), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_526), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_527), .A2(n_92), .B1(n_94), .B2(n_95), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_522), .Y(n_567) );
INVx4_ASAP7_75t_L g568 ( .A(n_494), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_523), .Y(n_569) );
OR2x6_ASAP7_75t_L g570 ( .A(n_494), .B(n_94), .Y(n_570) );
OAI21x1_ASAP7_75t_L g571 ( .A1(n_520), .A2(n_174), .B(n_201), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_501), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_475), .Y(n_573) );
INVx3_ASAP7_75t_SL g574 ( .A(n_533), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_495), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_523), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_492), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_492), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_481), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g580 ( .A1(n_480), .A2(n_145), .B(n_148), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_517), .B(n_149), .Y(n_581) );
AO31x2_ASAP7_75t_L g582 ( .A1(n_504), .A2(n_150), .A3(n_151), .B(n_153), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_523), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_511), .B(n_159), .Y(n_584) );
OA21x2_ASAP7_75t_L g585 ( .A1(n_488), .A2(n_161), .B(n_162), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_481), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_531), .A2(n_163), .B(n_165), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_506), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_506), .Y(n_589) );
OA21x2_ASAP7_75t_L g590 ( .A1(n_530), .A2(n_181), .B(n_182), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_483), .B(n_183), .Y(n_591) );
OA21x2_ASAP7_75t_L g592 ( .A1(n_508), .A2(n_184), .B(n_185), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_528), .B(n_186), .Y(n_593) );
AO21x2_ASAP7_75t_L g594 ( .A1(n_524), .A2(n_189), .B(n_191), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_484), .A2(n_192), .B(n_193), .Y(n_595) );
OA21x2_ASAP7_75t_L g596 ( .A1(n_496), .A2(n_194), .B(n_195), .Y(n_596) );
AOI21xp33_ASAP7_75t_L g597 ( .A1(n_484), .A2(n_197), .B(n_198), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_510), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_502), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_510), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_510), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_532), .Y(n_602) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_487), .A2(n_477), .B(n_489), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_532), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_532), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_513), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_518), .B(n_516), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_516), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_486), .A2(n_535), .B1(n_500), .B2(n_538), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_474), .B(n_473), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_539), .B(n_536), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_502), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_473), .B(n_539), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_518), .B(n_516), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_473), .B(n_502), .Y(n_615) );
OR2x6_ASAP7_75t_L g616 ( .A(n_570), .B(n_515), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_552), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_543), .B(n_537), .Y(n_618) );
INVx8_ASAP7_75t_L g619 ( .A(n_570), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_572), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_579), .Y(n_621) );
AO21x2_ASAP7_75t_L g622 ( .A1(n_615), .A2(n_610), .B(n_589), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_553), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_554), .Y(n_624) );
AO21x2_ASAP7_75t_L g625 ( .A1(n_588), .A2(n_600), .B(n_598), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_561), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_586), .Y(n_627) );
OA21x2_ASAP7_75t_L g628 ( .A1(n_599), .A2(n_612), .B(n_562), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_613), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_563), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_565), .B(n_542), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_577), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_565), .B(n_575), .Y(n_633) );
OA21x2_ASAP7_75t_L g634 ( .A1(n_560), .A2(n_576), .B(n_569), .Y(n_634) );
BUFx2_ASAP7_75t_L g635 ( .A(n_574), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_548), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_545), .B(n_567), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_548), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_613), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_583), .B(n_566), .Y(n_640) );
AO21x2_ASAP7_75t_L g641 ( .A1(n_601), .A2(n_604), .B(n_605), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_549), .Y(n_642) );
OR2x6_ASAP7_75t_L g643 ( .A(n_568), .B(n_581), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_609), .A2(n_593), .B(n_584), .Y(n_644) );
AOI21x1_ASAP7_75t_L g645 ( .A1(n_602), .A2(n_608), .B(n_559), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_581), .Y(n_646) );
OA21x2_ASAP7_75t_L g647 ( .A1(n_607), .A2(n_614), .B(n_597), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_591), .Y(n_648) );
AO21x2_ASAP7_75t_L g649 ( .A1(n_550), .A2(n_603), .B(n_595), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_590), .Y(n_650) );
AO21x2_ASAP7_75t_L g651 ( .A1(n_603), .A2(n_580), .B(n_546), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_555), .Y(n_652) );
OR2x6_ASAP7_75t_L g653 ( .A(n_544), .B(n_578), .Y(n_653) );
AOI21x1_ASAP7_75t_L g654 ( .A1(n_556), .A2(n_611), .B(n_592), .Y(n_654) );
AO21x2_ASAP7_75t_L g655 ( .A1(n_580), .A2(n_546), .B(n_551), .Y(n_655) );
OR2x6_ASAP7_75t_L g656 ( .A(n_577), .B(n_578), .Y(n_656) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_571), .Y(n_657) );
BUFx3_ASAP7_75t_L g658 ( .A(n_582), .Y(n_658) );
OR2x6_ASAP7_75t_L g659 ( .A(n_587), .B(n_557), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_558), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_582), .B(n_594), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_585), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_596), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_541), .B(n_547), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_541), .B(n_547), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_563), .Y(n_666) );
OA21x2_ASAP7_75t_L g667 ( .A1(n_615), .A2(n_485), .B(n_599), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_564), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_540), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_573), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_606), .Y(n_671) );
AOI21xp5_ASAP7_75t_SL g672 ( .A1(n_570), .A2(n_609), .B(n_592), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_629), .B(n_639), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_645), .Y(n_674) );
CKINVDCx5p33_ASAP7_75t_R g675 ( .A(n_635), .Y(n_675) );
INVx5_ASAP7_75t_L g676 ( .A(n_643), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_637), .B(n_640), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_637), .B(n_640), .Y(n_678) );
INVx3_ASAP7_75t_L g679 ( .A(n_632), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_664), .B(n_665), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_642), .B(n_620), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_633), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_634), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_621), .B(n_627), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_668), .B(n_652), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_641), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_618), .B(n_631), .Y(n_687) );
INVx2_ASAP7_75t_SL g688 ( .A(n_632), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_643), .Y(n_689) );
AND2x4_ASAP7_75t_L g690 ( .A(n_625), .B(n_670), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_669), .B(n_617), .Y(n_691) );
INVx2_ASAP7_75t_SL g692 ( .A(n_656), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_628), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_628), .Y(n_694) );
INVx4_ASAP7_75t_L g695 ( .A(n_619), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_623), .B(n_624), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_622), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_647), .B(n_648), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_647), .B(n_626), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_667), .B(n_646), .Y(n_700) );
BUFx2_ASAP7_75t_L g701 ( .A(n_636), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_658), .B(n_649), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_658), .B(n_649), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_661), .B(n_672), .Y(n_704) );
BUFx2_ASAP7_75t_L g705 ( .A(n_638), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_651), .B(n_630), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_666), .B(n_644), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_693), .Y(n_708) );
INVx1_ASAP7_75t_SL g709 ( .A(n_675), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_700), .B(n_616), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_691), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_687), .B(n_671), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_673), .B(n_653), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_673), .B(n_653), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_677), .B(n_663), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_678), .B(n_662), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_680), .B(n_666), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_694), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_699), .B(n_660), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_698), .B(n_650), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_696), .Y(n_721) );
INVx4_ASAP7_75t_L g722 ( .A(n_676), .Y(n_722) );
BUFx3_ASAP7_75t_L g723 ( .A(n_701), .Y(n_723) );
BUFx3_ASAP7_75t_L g724 ( .A(n_705), .Y(n_724) );
BUFx3_ASAP7_75t_L g725 ( .A(n_705), .Y(n_725) );
OR2x6_ASAP7_75t_L g726 ( .A(n_689), .B(n_657), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_684), .B(n_655), .Y(n_727) );
AND2x4_ASAP7_75t_L g728 ( .A(n_704), .B(n_657), .Y(n_728) );
INVx3_ASAP7_75t_L g729 ( .A(n_690), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_682), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_685), .B(n_654), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_681), .B(n_659), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_685), .B(n_657), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_683), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_730), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_708), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_711), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_712), .Y(n_738) );
OR2x6_ASAP7_75t_L g739 ( .A(n_723), .B(n_689), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_721), .Y(n_740) );
NAND2xp33_ASAP7_75t_SL g741 ( .A(n_722), .B(n_695), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_712), .Y(n_742) );
INVxp67_ASAP7_75t_L g743 ( .A(n_723), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_716), .B(n_706), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_716), .B(n_706), .Y(n_745) );
INVx2_ASAP7_75t_SL g746 ( .A(n_724), .Y(n_746) );
OR2x2_ASAP7_75t_L g747 ( .A(n_715), .B(n_686), .Y(n_747) );
OR2x6_ASAP7_75t_L g748 ( .A(n_725), .B(n_707), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_718), .Y(n_749) );
INVx1_ASAP7_75t_SL g750 ( .A(n_709), .Y(n_750) );
INVx1_ASAP7_75t_SL g751 ( .A(n_750), .Y(n_751) );
INVx1_ASAP7_75t_SL g752 ( .A(n_741), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_736), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_742), .A2(n_710), .B1(n_732), .B2(n_717), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_738), .B(n_713), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_743), .B(n_732), .C(n_734), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_736), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_751), .B(n_735), .Y(n_758) );
NAND2x1p5_ASAP7_75t_L g759 ( .A(n_752), .B(n_746), .Y(n_759) );
INVxp67_ASAP7_75t_L g760 ( .A(n_756), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_760), .A2(n_755), .B1(n_754), .B2(n_740), .C(n_737), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_759), .B(n_753), .Y(n_762) );
AOI21xp33_ASAP7_75t_L g763 ( .A1(n_758), .A2(n_692), .B(n_713), .Y(n_763) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_759), .A2(n_748), .B1(n_739), .B2(n_747), .C(n_714), .Y(n_764) );
AOI322xp5_ASAP7_75t_L g765 ( .A1(n_761), .A2(n_744), .A3(n_745), .B1(n_731), .B2(n_757), .C1(n_727), .C2(n_719), .Y(n_765) );
OAI211xp5_ASAP7_75t_SL g766 ( .A1(n_765), .A2(n_764), .B(n_762), .C(n_763), .Y(n_766) );
OR5x1_ASAP7_75t_L g767 ( .A(n_766), .B(n_726), .C(n_728), .D(n_729), .E(n_688), .Y(n_767) );
XNOR2x1_ASAP7_75t_L g768 ( .A(n_767), .B(n_659), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_768), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_769), .A2(n_674), .B(n_697), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_770), .B(n_749), .Y(n_771) );
OR2x6_ASAP7_75t_L g772 ( .A(n_771), .B(n_679), .Y(n_772) );
OAI21xp5_ASAP7_75t_SL g773 ( .A1(n_772), .A2(n_733), .B(n_720), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_773), .A2(n_733), .B1(n_702), .B2(n_703), .Y(n_774) );
endmodule