module fake_jpeg_19578_n_176 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx5_ASAP7_75t_SL g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_27),
.B1(n_21),
.B2(n_15),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_46),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_27),
.B1(n_15),
.B2(n_26),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_38),
.B1(n_30),
.B2(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_22),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_23),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_21),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_57),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_26),
.B(n_22),
.C(n_17),
.Y(n_58)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_50),
.B(n_46),
.C(n_39),
.D(n_16),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_60),
.B(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_68),
.Y(n_75)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_39),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_44),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_44),
.B1(n_49),
.B2(n_45),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_73),
.B(n_74),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_43),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_78),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_43),
.B1(n_40),
.B2(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_32),
.C(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_59),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_45),
.A3(n_49),
.B1(n_31),
.B2(n_32),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_44),
.B(n_49),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_88),
.B(n_62),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_67),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_69),
.C(n_39),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_44),
.Y(n_93)
);

OAI31xp33_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_63),
.A3(n_61),
.B(n_59),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_70),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_104),
.C(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_100),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_107),
.B1(n_85),
.B2(n_79),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_58),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_77),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_60),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_119),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_80),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_118),
.A2(n_115),
.B(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_102),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_78),
.B1(n_93),
.B2(n_83),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_94),
.B1(n_98),
.B2(n_90),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_82),
.C(n_77),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_97),
.C(n_91),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_30),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_76),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_134),
.C(n_118),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_100),
.B(n_105),
.C(n_94),
.D(n_88),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_135),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_80),
.C(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_138),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_1),
.B(n_2),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_115),
.B(n_116),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_137),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_10),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_143),
.A2(n_4),
.B(n_5),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_147),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_120),
.C(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_4),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_120),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_117),
.B1(n_126),
.B2(n_125),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_133),
.B(n_128),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_151),
.A2(n_9),
.B(n_11),
.Y(n_163)
);

NOR4xp25_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_125),
.C(n_134),
.D(n_112),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_141),
.B(n_142),
.C(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_112),
.C(n_67),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_24),
.C(n_16),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_157),
.B(n_6),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_142),
.B(n_7),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_162),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_160),
.C(n_161),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_153),
.B(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_13),
.B(n_6),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_174),
.C(n_172),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_166),
.B(n_6),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_175),
.B(n_7),
.Y(n_176)
);


endmodule