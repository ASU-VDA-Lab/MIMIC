module fake_netlist_1_7111_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g10 ( .A(n_2), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_5), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_12), .B(n_0), .Y(n_17) );
BUFx4f_ASAP7_75t_L g18 ( .A(n_10), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_13), .B(n_0), .Y(n_20) );
OAI21xp33_ASAP7_75t_L g21 ( .A1(n_10), .A2(n_0), .B(n_9), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
NAND2xp5_ASAP7_75t_SL g23 ( .A(n_18), .B(n_12), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_20), .A2(n_11), .B1(n_15), .B2(n_14), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_18), .A2(n_16), .B1(n_2), .B2(n_3), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_20), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_24), .A2(n_18), .B1(n_17), .B2(n_21), .Y(n_28) );
AOI22xp33_ASAP7_75t_L g29 ( .A1(n_23), .A2(n_22), .B1(n_19), .B2(n_7), .Y(n_29) );
AND2x4_ASAP7_75t_L g30 ( .A(n_27), .B(n_26), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g31 ( .A(n_27), .B(n_22), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_28), .B(n_19), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_30), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_30), .B(n_29), .Y(n_35) );
OAI211xp5_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_32), .B(n_4), .C(n_7), .Y(n_36) );
AOI21xp5_ASAP7_75t_L g37 ( .A1(n_33), .A2(n_1), .B(n_9), .Y(n_37) );
BUFx2_ASAP7_75t_L g38 ( .A(n_34), .Y(n_38) );
A2O1A1Ixp33_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_35), .B(n_37), .C(n_38), .Y(n_39) );
INVx1_ASAP7_75t_SL g40 ( .A(n_38), .Y(n_40) );
NAND2xp33_ASAP7_75t_L g41 ( .A(n_40), .B(n_39), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_41), .Y(n_42) );
endmodule