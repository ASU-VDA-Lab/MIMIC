module fake_ariane_336_n_1599 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_1599);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_1599;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_334;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_552;
wire n_348;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_1552;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1587;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1477;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1571;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_275;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g230 ( 
.A(n_115),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_113),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_37),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_193),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_81),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_63),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_145),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_29),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_92),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_127),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_152),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_5),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_17),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_62),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_229),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_97),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_151),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_1),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_76),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_41),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_44),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_100),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_136),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_41),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_56),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_130),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_202),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_162),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_144),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_175),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_158),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_80),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_124),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_111),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_131),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_45),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_13),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_208),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_103),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_38),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_108),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_122),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_86),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_51),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_201),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_101),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_116),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_18),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_29),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_57),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_39),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_82),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_196),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_77),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_226),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_93),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_166),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_191),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_179),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_120),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_39),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g294 ( 
.A(n_227),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_155),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_56),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_34),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_164),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_110),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_200),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_74),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_96),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_40),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_194),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_95),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_52),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_62),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_85),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_171),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_223),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_105),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_55),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_11),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_224),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_206),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_43),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_173),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_135),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_172),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_73),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_118),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_54),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_47),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_114),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_104),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_33),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_38),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_94),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_184),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_51),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_24),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_21),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_148),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_125),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_7),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_46),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_119),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_75),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_91),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_71),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_50),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_212),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_112),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_99),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_205),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_13),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_174),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_102),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_28),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_187),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_167),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_153),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_64),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_117),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_72),
.Y(n_355)
);

BUFx8_ASAP7_75t_SL g356 ( 
.A(n_220),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_16),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_209),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_176),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_22),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_128),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_67),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_225),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_47),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_181),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_165),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_142),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_14),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_20),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_356),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_236),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_236),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_236),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_236),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_303),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_356),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_242),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_245),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_245),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_242),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_268),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_303),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_303),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_285),
.B(n_0),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_299),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_323),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_320),
.B(n_0),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_323),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_293),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_248),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_230),
.B(n_231),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_232),
.B(n_1),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_263),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_296),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_261),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_248),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_238),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_281),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_299),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_307),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_281),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_306),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_367),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_315),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_R g408 ( 
.A(n_241),
.B(n_68),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_306),
.B(n_2),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_254),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_312),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_312),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_330),
.B(n_2),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_315),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_235),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_313),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_239),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_235),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_316),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_261),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_278),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_326),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_278),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_327),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_336),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_353),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_347),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_301),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_247),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_368),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_347),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_301),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_337),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_330),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_343),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_254),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_343),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_243),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_252),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_346),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_341),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_257),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_354),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_250),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_346),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_341),
.B(n_3),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_364),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_354),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_349),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_244),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_251),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_364),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_255),
.B(n_3),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_264),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_406),
.B(n_249),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_398),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_379),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_398),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_419),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_370),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_442),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_SL g467 ( 
.A(n_447),
.B(n_244),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_453),
.A2(n_267),
.B1(n_282),
.B2(n_276),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_398),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_419),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_422),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_422),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_406),
.B(n_266),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_424),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_449),
.B(n_271),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_424),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_411),
.B(n_418),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_398),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_455),
.Y(n_480)
);

NOR2x1_ASAP7_75t_L g481 ( 
.A(n_429),
.B(n_240),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_411),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_421),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_429),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_418),
.B(n_274),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_430),
.B(n_290),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_421),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_421),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_430),
.B(n_295),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_433),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_421),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_421),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_259),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_449),
.B(n_283),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_441),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_371),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_441),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_433),
.Y(n_498)
);

OA21x2_ASAP7_75t_L g499 ( 
.A1(n_434),
.A2(n_305),
.B(n_300),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_434),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_371),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_436),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_436),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_372),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_381),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_410),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_437),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_372),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_444),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_444),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_396),
.B(n_241),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_385),
.B(n_233),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_373),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_438),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_439),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_439),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_373),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_374),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_380),
.A2(n_282),
.B1(n_267),
.B2(n_280),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_374),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_375),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_375),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_376),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_376),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_383),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_382),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_378),
.B(n_262),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_389),
.B1(n_395),
.B2(n_456),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_513),
.B(n_392),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_513),
.B(n_397),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_481),
.B(n_435),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_514),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_458),
.B(n_457),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_481),
.B(n_443),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_480),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_518),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_461),
.Y(n_538)
);

NAND3x1_ASAP7_75t_L g539 ( 
.A(n_476),
.B(n_448),
.C(n_414),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_458),
.B(n_403),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_518),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_467),
.A2(n_408),
.B1(n_322),
.B2(n_357),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_496),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_482),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_514),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_514),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_514),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_482),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_512),
.B(n_417),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_519),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_499),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_519),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_466),
.B(n_420),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_515),
.B(n_423),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_501),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_522),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_493),
.B(n_456),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_480),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_493),
.B(n_425),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_466),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_522),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_524),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_482),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_515),
.B(n_426),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_524),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_526),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_499),
.A2(n_394),
.B1(n_446),
.B2(n_400),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_527),
.B(n_427),
.Y(n_568)
);

AND2x2_ASAP7_75t_SL g569 ( 
.A(n_499),
.B(n_261),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_501),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_465),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_478),
.B(n_409),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_526),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_501),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_496),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_493),
.B(n_431),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_493),
.B(n_440),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_475),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_460),
.Y(n_579)
);

CKINVDCx14_ASAP7_75t_R g580 ( 
.A(n_465),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_504),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_460),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_505),
.B(n_450),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_505),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_462),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_520),
.B(n_377),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_462),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_495),
.B(n_383),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_464),
.B(n_261),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_499),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_495),
.B(n_440),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_476),
.B(n_451),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_537),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_537),
.Y(n_595)
);

OAI221xp5_ASAP7_75t_L g596 ( 
.A1(n_529),
.A2(n_360),
.B1(n_335),
.B2(n_332),
.C(n_369),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_L g597 ( 
.A(n_554),
.B(n_506),
.C(n_520),
.Y(n_597)
);

OAI221xp5_ASAP7_75t_L g598 ( 
.A1(n_542),
.A2(n_331),
.B1(n_297),
.B2(n_489),
.C(n_486),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_541),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_577),
.B(n_494),
.Y(n_600)
);

BUFx8_ASAP7_75t_L g601 ( 
.A(n_560),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_539),
.A2(n_506),
.B1(n_494),
.B2(n_497),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_543),
.Y(n_603)
);

OR2x2_ASAP7_75t_SL g604 ( 
.A(n_583),
.B(n_386),
.Y(n_604)
);

BUFx8_ASAP7_75t_L g605 ( 
.A(n_560),
.Y(n_605)
);

NAND2x1p5_ASAP7_75t_L g606 ( 
.A(n_571),
.B(n_495),
.Y(n_606)
);

AO22x2_ASAP7_75t_L g607 ( 
.A1(n_583),
.A2(n_468),
.B1(n_407),
.B2(n_415),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_536),
.B(n_495),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_580),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_541),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_550),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_540),
.B(n_402),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_550),
.Y(n_613)
);

NAND2x1p5_ASAP7_75t_L g614 ( 
.A(n_536),
.B(n_497),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_552),
.Y(n_615)
);

AO22x2_ASAP7_75t_L g616 ( 
.A1(n_530),
.A2(n_468),
.B1(n_432),
.B2(n_445),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_539),
.A2(n_509),
.B1(n_510),
.B2(n_497),
.Y(n_617)
);

AO22x2_ASAP7_75t_L g618 ( 
.A1(n_531),
.A2(n_428),
.B1(n_486),
.B2(n_485),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_532),
.B(n_497),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_564),
.B(n_452),
.Y(n_620)
);

AO22x2_ASAP7_75t_L g621 ( 
.A1(n_557),
.A2(n_489),
.B1(n_485),
.B2(n_478),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_532),
.B(n_509),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_532),
.B(n_509),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_586),
.B(n_246),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_532),
.B(n_509),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_552),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_556),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_556),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_561),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_577),
.B(n_454),
.Y(n_630)
);

BUFx8_ASAP7_75t_L g631 ( 
.A(n_584),
.Y(n_631)
);

OAI221xp5_ASAP7_75t_L g632 ( 
.A1(n_542),
.A2(n_473),
.B1(n_454),
.B2(n_500),
.C(n_517),
.Y(n_632)
);

AO22x2_ASAP7_75t_L g633 ( 
.A1(n_557),
.A2(n_584),
.B1(n_558),
.B2(n_535),
.Y(n_633)
);

OAI221xp5_ASAP7_75t_L g634 ( 
.A1(n_567),
.A2(n_473),
.B1(n_500),
.B2(n_477),
.C(n_517),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_535),
.A2(n_572),
.B1(n_569),
.B2(n_557),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_555),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_558),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_561),
.Y(n_638)
);

INVxp33_ASAP7_75t_L g639 ( 
.A(n_568),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_562),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_562),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_565),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_555),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_535),
.B(n_510),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_538),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_565),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_566),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_538),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_566),
.Y(n_649)
);

AO22x2_ASAP7_75t_L g650 ( 
.A1(n_557),
.A2(n_471),
.B1(n_472),
.B2(n_470),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_577),
.B(n_510),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_573),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_573),
.Y(n_653)
);

AO22x2_ASAP7_75t_L g654 ( 
.A1(n_535),
.A2(n_592),
.B1(n_553),
.B2(n_576),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_534),
.B(n_577),
.Y(n_655)
);

BUFx8_ASAP7_75t_L g656 ( 
.A(n_591),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_570),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_591),
.B(n_510),
.Y(n_658)
);

AO22x2_ASAP7_75t_L g659 ( 
.A1(n_559),
.A2(n_471),
.B1(n_472),
.B2(n_470),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_549),
.A2(n_477),
.B1(n_484),
.B2(n_474),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_579),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_579),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_544),
.B(n_474),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_582),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_582),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_585),
.Y(n_666)
);

OR2x6_ASAP7_75t_L g667 ( 
.A(n_572),
.B(n_484),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_585),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_570),
.Y(n_669)
);

OAI221xp5_ASAP7_75t_L g670 ( 
.A1(n_587),
.A2(n_593),
.B1(n_498),
.B2(n_507),
.C(n_502),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_572),
.B(n_490),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_587),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_593),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_588),
.Y(n_674)
);

AO22x2_ASAP7_75t_L g675 ( 
.A1(n_551),
.A2(n_498),
.B1(n_502),
.B2(n_490),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_572),
.A2(n_507),
.B1(n_511),
.B2(n_503),
.Y(n_676)
);

AO22x2_ASAP7_75t_L g677 ( 
.A1(n_551),
.A2(n_511),
.B1(n_516),
.B2(n_503),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_572),
.B(n_516),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_544),
.B(n_393),
.Y(n_679)
);

AO22x2_ASAP7_75t_L g680 ( 
.A1(n_551),
.A2(n_399),
.B1(n_401),
.B2(n_393),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_630),
.B(n_548),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_630),
.B(n_548),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_600),
.B(n_399),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_600),
.B(n_401),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_SL g685 ( 
.A(n_639),
.B(n_578),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_637),
.B(n_563),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_655),
.B(n_563),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_631),
.B(n_578),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_631),
.B(n_578),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_635),
.B(n_578),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_678),
.B(n_543),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_678),
.B(n_543),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_624),
.B(n_543),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_612),
.B(n_679),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_679),
.B(n_543),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_608),
.B(n_575),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_614),
.B(n_575),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_651),
.B(n_569),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_676),
.B(n_575),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_606),
.B(n_575),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_602),
.B(n_575),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_620),
.B(n_594),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_597),
.B(n_404),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_594),
.B(n_533),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_595),
.B(n_533),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_595),
.B(n_545),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_671),
.B(n_660),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_663),
.B(n_545),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_633),
.B(n_569),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_599),
.B(n_546),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_633),
.B(n_619),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_SL g712 ( 
.A(n_609),
.B(n_546),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_622),
.B(n_547),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_610),
.B(n_547),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_611),
.B(n_551),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_613),
.B(n_590),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_615),
.B(n_590),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_626),
.B(n_590),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_627),
.B(n_590),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_SL g720 ( 
.A(n_628),
.B(n_246),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_629),
.B(n_253),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_638),
.B(n_640),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_641),
.B(n_253),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_SL g724 ( 
.A(n_642),
.B(n_256),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_646),
.B(n_256),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_647),
.B(n_258),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_623),
.B(n_574),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_649),
.B(n_258),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_652),
.B(n_340),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_603),
.B(n_574),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_653),
.B(n_340),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_SL g732 ( 
.A(n_661),
.B(n_342),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_SL g733 ( 
.A(n_662),
.B(n_342),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_664),
.B(n_344),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_665),
.B(n_666),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_668),
.B(n_344),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_672),
.B(n_348),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_625),
.B(n_581),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_673),
.B(n_656),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_SL g740 ( 
.A(n_603),
.B(n_348),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_656),
.B(n_350),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_601),
.B(n_350),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_601),
.B(n_351),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_644),
.B(n_581),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_605),
.B(n_351),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_605),
.B(n_352),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_617),
.B(n_352),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_667),
.B(n_404),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_SL g749 ( 
.A(n_603),
.B(n_658),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_SL g750 ( 
.A(n_674),
.B(n_234),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_645),
.B(n_648),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_636),
.B(n_237),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_643),
.B(n_265),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_657),
.B(n_269),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_669),
.B(n_273),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_632),
.B(n_499),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_650),
.B(n_277),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_650),
.B(n_279),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_654),
.B(n_284),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_654),
.B(n_286),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_667),
.B(n_287),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_621),
.B(n_288),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_621),
.B(n_289),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_659),
.B(n_291),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_659),
.B(n_292),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_SL g766 ( 
.A(n_596),
.B(n_302),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_680),
.B(n_304),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_598),
.B(n_504),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_680),
.B(n_308),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_675),
.B(n_317),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_675),
.B(n_405),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_677),
.B(n_318),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_618),
.B(n_504),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_677),
.B(n_319),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_670),
.B(n_321),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_618),
.B(n_523),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_604),
.B(n_309),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_634),
.B(n_475),
.Y(n_778)
);

OAI21x1_ASAP7_75t_L g779 ( 
.A1(n_730),
.A2(n_523),
.B(n_463),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_715),
.A2(n_260),
.B(n_259),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_681),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_685),
.A2(n_270),
.B(n_260),
.Y(n_782)
);

NOR2xp67_ASAP7_75t_L g783 ( 
.A(n_694),
.B(n_405),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_722),
.Y(n_784)
);

OA21x2_ASAP7_75t_L g785 ( 
.A1(n_773),
.A2(n_523),
.B(n_463),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_707),
.B(n_616),
.Y(n_786)
);

AO31x2_ASAP7_75t_L g787 ( 
.A1(n_776),
.A2(n_412),
.A3(n_413),
.B(n_387),
.Y(n_787)
);

OAI21x1_ASAP7_75t_L g788 ( 
.A1(n_730),
.A2(n_463),
.B(n_459),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_716),
.A2(n_311),
.B(n_310),
.Y(n_789)
);

AO21x2_ASAP7_75t_L g790 ( 
.A1(n_762),
.A2(n_324),
.B(n_314),
.Y(n_790)
);

OAI21x1_ASAP7_75t_L g791 ( 
.A1(n_717),
.A2(n_469),
.B(n_459),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_718),
.A2(n_275),
.B(n_270),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_735),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_719),
.A2(n_275),
.B(n_459),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_699),
.A2(n_487),
.B(n_469),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_710),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_727),
.A2(n_487),
.B(n_469),
.Y(n_797)
);

AO21x1_ASAP7_75t_L g798 ( 
.A1(n_693),
.A2(n_701),
.B(n_771),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_681),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_683),
.B(n_412),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_681),
.B(n_748),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_766),
.A2(n_366),
.B(n_358),
.C(n_359),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_684),
.Y(n_803)
);

OA21x2_ASAP7_75t_L g804 ( 
.A1(n_763),
.A2(n_491),
.B(n_487),
.Y(n_804)
);

AO31x2_ASAP7_75t_L g805 ( 
.A1(n_709),
.A2(n_413),
.A3(n_391),
.B(n_387),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_748),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_698),
.B(n_616),
.Y(n_807)
);

OA21x2_ASAP7_75t_L g808 ( 
.A1(n_756),
.A2(n_491),
.B(n_334),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_SL g809 ( 
.A1(n_771),
.A2(n_345),
.B(n_329),
.Y(n_809)
);

OAI21x1_ASAP7_75t_L g810 ( 
.A1(n_738),
.A2(n_744),
.B(n_705),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_702),
.B(n_713),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_748),
.B(n_607),
.Y(n_812)
);

OAI21x1_ASAP7_75t_SL g813 ( 
.A1(n_682),
.A2(n_363),
.B(n_362),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_751),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_687),
.A2(n_328),
.B(n_325),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_739),
.B(n_384),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_688),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_720),
.B(n_732),
.C(n_724),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_704),
.A2(n_491),
.B(n_388),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_706),
.A2(n_488),
.B(n_475),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_750),
.A2(n_388),
.B(n_390),
.C(n_391),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_714),
.A2(n_488),
.B(n_475),
.Y(n_822)
);

AO31x2_ASAP7_75t_L g823 ( 
.A1(n_711),
.A2(n_777),
.A3(n_768),
.B(n_765),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_733),
.B(n_333),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_771),
.A2(n_607),
.B1(n_384),
.B2(n_390),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_690),
.A2(n_496),
.B(n_525),
.C(n_521),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_778),
.A2(n_294),
.B(n_589),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_SL g828 ( 
.A(n_689),
.B(n_338),
.Y(n_828)
);

BUFx4f_ASAP7_75t_L g829 ( 
.A(n_703),
.Y(n_829)
);

OAI21x1_ASAP7_75t_L g830 ( 
.A1(n_778),
.A2(n_294),
.B(n_589),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_695),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_708),
.A2(n_355),
.B(n_339),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_691),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_696),
.A2(n_488),
.B(n_589),
.C(n_521),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_712),
.B(n_365),
.Y(n_835)
);

OAI22x1_ASAP7_75t_L g836 ( 
.A1(n_761),
.A2(n_488),
.B1(n_5),
.B2(n_6),
.Y(n_836)
);

OA21x2_ASAP7_75t_L g837 ( 
.A1(n_764),
.A2(n_294),
.B(n_496),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_692),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_697),
.A2(n_298),
.B(n_272),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_700),
.A2(n_294),
.B(n_589),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_721),
.B(n_4),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_770),
.A2(n_294),
.B(n_589),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_772),
.A2(n_294),
.B(n_589),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_723),
.B(n_4),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_686),
.Y(n_845)
);

BUFx6f_ASAP7_75t_SL g846 ( 
.A(n_741),
.Y(n_846)
);

AND2x6_ASAP7_75t_L g847 ( 
.A(n_749),
.B(n_272),
.Y(n_847)
);

AO31x2_ASAP7_75t_L g848 ( 
.A1(n_759),
.A2(n_589),
.A3(n_525),
.B(n_521),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_742),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_747),
.B(n_496),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_767),
.A2(n_525),
.B(n_521),
.C(n_508),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_760),
.B(n_496),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_769),
.Y(n_853)
);

AOI21xp33_ASAP7_75t_L g854 ( 
.A1(n_774),
.A2(n_508),
.B(n_496),
.Y(n_854)
);

AOI221x1_ASAP7_75t_L g855 ( 
.A1(n_740),
.A2(n_525),
.B1(n_521),
.B2(n_508),
.C(n_492),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_743),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_745),
.B(n_508),
.Y(n_857)
);

CKINVDCx6p67_ASAP7_75t_R g858 ( 
.A(n_746),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_775),
.A2(n_483),
.B(n_479),
.Y(n_859)
);

INVx8_ASAP7_75t_L g860 ( 
.A(n_757),
.Y(n_860)
);

OAI21x1_ASAP7_75t_L g861 ( 
.A1(n_758),
.A2(n_294),
.B(n_508),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_725),
.A2(n_521),
.B(n_508),
.Y(n_862)
);

AOI221x1_ASAP7_75t_L g863 ( 
.A1(n_726),
.A2(n_525),
.B1(n_521),
.B2(n_508),
.C(n_492),
.Y(n_863)
);

BUFx10_ASAP7_75t_L g864 ( 
.A(n_728),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_729),
.A2(n_492),
.B(n_483),
.Y(n_865)
);

AO31x2_ASAP7_75t_L g866 ( 
.A1(n_731),
.A2(n_525),
.A3(n_492),
.B(n_483),
.Y(n_866)
);

AOI21xp33_ASAP7_75t_L g867 ( 
.A1(n_734),
.A2(n_737),
.B(n_736),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_752),
.B(n_753),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_754),
.B(n_525),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_755),
.A2(n_272),
.B1(n_298),
.B2(n_361),
.Y(n_870)
);

OAI21x1_ASAP7_75t_L g871 ( 
.A1(n_730),
.A2(n_106),
.B(n_228),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_681),
.B(n_272),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_803),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_800),
.B(n_6),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_797),
.A2(n_492),
.B(n_483),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_795),
.A2(n_492),
.B(n_483),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_799),
.B(n_7),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_814),
.A2(n_361),
.B1(n_298),
.B2(n_479),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_827),
.A2(n_830),
.B(n_861),
.Y(n_879)
);

BUFx12f_ASAP7_75t_L g880 ( 
.A(n_856),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_841),
.A2(n_298),
.B(n_361),
.C(n_10),
.Y(n_881)
);

OA21x2_ASAP7_75t_L g882 ( 
.A1(n_863),
.A2(n_492),
.B(n_483),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_788),
.A2(n_483),
.B(n_479),
.Y(n_883)
);

NAND3xp33_ASAP7_75t_L g884 ( 
.A(n_802),
.B(n_361),
.C(n_479),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_781),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_859),
.A2(n_479),
.B(n_89),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_784),
.Y(n_887)
);

OA21x2_ASAP7_75t_L g888 ( 
.A1(n_810),
.A2(n_479),
.B(n_90),
.Y(n_888)
);

OAI21x1_ASAP7_75t_SL g889 ( 
.A1(n_811),
.A2(n_8),
.B(n_9),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_806),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_859),
.A2(n_479),
.B(n_88),
.Y(n_891)
);

OAI21x1_ASAP7_75t_L g892 ( 
.A1(n_791),
.A2(n_87),
.B(n_221),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_825),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_818),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_779),
.A2(n_109),
.B(n_219),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_801),
.B(n_12),
.Y(n_896)
);

CKINVDCx11_ASAP7_75t_R g897 ( 
.A(n_858),
.Y(n_897)
);

AO21x2_ASAP7_75t_L g898 ( 
.A1(n_852),
.A2(n_107),
.B(n_217),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_793),
.Y(n_899)
);

AO21x1_ASAP7_75t_L g900 ( 
.A1(n_844),
.A2(n_15),
.B(n_16),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_801),
.B(n_15),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_842),
.A2(n_843),
.B(n_840),
.Y(n_902)
);

OAI21xp33_ASAP7_75t_SL g903 ( 
.A1(n_811),
.A2(n_17),
.B(n_18),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_799),
.B(n_19),
.Y(n_904)
);

OAI21x1_ASAP7_75t_L g905 ( 
.A1(n_871),
.A2(n_123),
.B(n_215),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_783),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_812),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_845),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_829),
.B(n_19),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_867),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_833),
.Y(n_911)
);

AOI21x1_ASAP7_75t_L g912 ( 
.A1(n_855),
.A2(n_852),
.B(n_808),
.Y(n_912)
);

OR2x6_ASAP7_75t_L g913 ( 
.A(n_860),
.B(n_23),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_818),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_781),
.B(n_25),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_785),
.Y(n_916)
);

OA21x2_ASAP7_75t_L g917 ( 
.A1(n_826),
.A2(n_133),
.B(n_214),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_831),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_829),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_787),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_787),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_787),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_785),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_796),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_846),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_808),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_794),
.A2(n_132),
.B(n_211),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_782),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_786),
.Y(n_929)
);

AO21x2_ASAP7_75t_L g930 ( 
.A1(n_798),
.A2(n_129),
.B(n_210),
.Y(n_930)
);

OAI21x1_ASAP7_75t_SL g931 ( 
.A1(n_813),
.A2(n_26),
.B(n_27),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_786),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_794),
.A2(n_134),
.B(n_207),
.Y(n_933)
);

AO21x1_ASAP7_75t_L g934 ( 
.A1(n_870),
.A2(n_854),
.B(n_780),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_865),
.A2(n_126),
.B(n_204),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_789),
.A2(n_30),
.B(n_31),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_865),
.A2(n_121),
.B(n_203),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_825),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_938)
);

INVxp67_ASAP7_75t_SL g939 ( 
.A(n_872),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_807),
.B(n_32),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_807),
.B(n_33),
.Y(n_941)
);

OAI221xp5_ASAP7_75t_L g942 ( 
.A1(n_853),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.C(n_37),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_839),
.A2(n_139),
.B(n_199),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_854),
.B(n_35),
.C(n_36),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_823),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_819),
.A2(n_140),
.B(n_198),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_789),
.A2(n_40),
.B(n_42),
.Y(n_947)
);

NAND2x1p5_ASAP7_75t_L g948 ( 
.A(n_838),
.B(n_141),
.Y(n_948)
);

OAI21x1_ASAP7_75t_L g949 ( 
.A1(n_804),
.A2(n_138),
.B(n_197),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_849),
.B(n_42),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_817),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_856),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_823),
.B(n_43),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_860),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_864),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_804),
.A2(n_147),
.B(n_195),
.Y(n_956)
);

NOR2xp67_ASAP7_75t_SL g957 ( 
.A(n_809),
.B(n_48),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_780),
.A2(n_851),
.B(n_862),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_823),
.Y(n_959)
);

AO21x2_ASAP7_75t_L g960 ( 
.A1(n_862),
.A2(n_146),
.B(n_192),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_846),
.Y(n_961)
);

OAI21x1_ASAP7_75t_L g962 ( 
.A1(n_837),
.A2(n_143),
.B(n_190),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_860),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_864),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_816),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_837),
.A2(n_137),
.B(n_189),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_834),
.A2(n_98),
.B(n_188),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_866),
.Y(n_968)
);

AO21x2_ASAP7_75t_L g969 ( 
.A1(n_792),
.A2(n_84),
.B(n_186),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_866),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_790),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_816),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_838),
.B(n_49),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_850),
.A2(n_149),
.B(n_185),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_857),
.B(n_52),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_868),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_R g977 ( 
.A1(n_836),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_977)
);

OAI21x1_ASAP7_75t_SL g978 ( 
.A1(n_867),
.A2(n_53),
.B(n_57),
.Y(n_978)
);

OR2x6_ASAP7_75t_L g979 ( 
.A(n_835),
.B(n_58),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_850),
.A2(n_156),
.B(n_183),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_824),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_SL g982 ( 
.A(n_847),
.B(n_154),
.Y(n_982)
);

CKINVDCx11_ASAP7_75t_R g983 ( 
.A(n_870),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_916),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_975),
.B(n_805),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_920),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_921),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_916),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_877),
.B(n_790),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_975),
.B(n_805),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_953),
.B(n_805),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_922),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_885),
.B(n_848),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_875),
.A2(n_869),
.B(n_820),
.Y(n_994)
);

AO21x2_ASAP7_75t_L g995 ( 
.A1(n_912),
.A2(n_926),
.B(n_945),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_959),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_897),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_923),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_926),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_968),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_911),
.B(n_848),
.Y(n_1001)
);

NAND2x1_ASAP7_75t_L g1002 ( 
.A(n_888),
.B(n_847),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_968),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_970),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_970),
.Y(n_1005)
);

OA21x2_ASAP7_75t_L g1006 ( 
.A1(n_875),
.A2(n_869),
.B(n_820),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_929),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_932),
.B(n_848),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_877),
.B(n_828),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_918),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_919),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_908),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_924),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_887),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_952),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_899),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_930),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_919),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_891),
.A2(n_822),
.B(n_815),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_888),
.Y(n_1020)
);

INVxp33_ASAP7_75t_L g1021 ( 
.A(n_897),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_930),
.Y(n_1022)
);

OR2x6_ASAP7_75t_L g1023 ( 
.A(n_976),
.B(n_822),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_888),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_890),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_898),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_885),
.B(n_976),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_898),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_898),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_948),
.B(n_821),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_885),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_873),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_940),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_891),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_881),
.A2(n_832),
.B(n_847),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_949),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_952),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_974),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_893),
.A2(n_847),
.B1(n_60),
.B2(n_61),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_949),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_956),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_951),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_974),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_956),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_902),
.A2(n_866),
.B(n_159),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_980),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_980),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_948),
.Y(n_1048)
);

AO21x2_ASAP7_75t_L g1049 ( 
.A1(n_958),
.A2(n_157),
.B(n_182),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_963),
.Y(n_1050)
);

OR2x6_ASAP7_75t_L g1051 ( 
.A(n_913),
.B(n_150),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_882),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_962),
.Y(n_1053)
);

OA21x2_ASAP7_75t_L g1054 ( 
.A1(n_883),
.A2(n_59),
.B(n_61),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_896),
.B(n_63),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_882),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_907),
.B(n_64),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_960),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_874),
.B(n_65),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_909),
.B(n_65),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_960),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_882),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_964),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_951),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_902),
.A2(n_163),
.B(n_69),
.Y(n_1065)
);

CKINVDCx12_ASAP7_75t_R g1066 ( 
.A(n_913),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_935),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_935),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_937),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_963),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_962),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_966),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_SL g1073 ( 
.A1(n_881),
.A2(n_168),
.B(n_70),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_937),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_904),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_1015),
.B(n_964),
.Y(n_1076)
);

XNOR2xp5_ASAP7_75t_L g1077 ( 
.A(n_1063),
.B(n_925),
.Y(n_1077)
);

XNOR2xp5_ASAP7_75t_L g1078 ( 
.A(n_997),
.B(n_925),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_R g1079 ( 
.A(n_1051),
.B(n_913),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_1025),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_R g1081 ( 
.A(n_1051),
.B(n_913),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_1064),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1032),
.B(n_941),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_1064),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_1075),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1013),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_1027),
.B(n_965),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1007),
.B(n_973),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_1027),
.B(n_896),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_1037),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1007),
.B(n_973),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1027),
.B(n_961),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_1027),
.B(n_906),
.Y(n_1093)
);

BUFx10_ASAP7_75t_L g1094 ( 
.A(n_1060),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_1018),
.Y(n_1095)
);

NAND2xp33_ASAP7_75t_R g1096 ( 
.A(n_1051),
.B(n_950),
.Y(n_1096)
);

NAND2xp33_ASAP7_75t_R g1097 ( 
.A(n_1051),
.B(n_979),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1013),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_1059),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1010),
.Y(n_1100)
);

BUFx10_ASAP7_75t_L g1101 ( 
.A(n_1051),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_R g1102 ( 
.A(n_1009),
.B(n_979),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1033),
.B(n_915),
.Y(n_1103)
);

NAND2xp33_ASAP7_75t_R g1104 ( 
.A(n_1033),
.B(n_979),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1012),
.B(n_1010),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_SL g1106 ( 
.A(n_1018),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1012),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_1057),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_989),
.B(n_915),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1055),
.B(n_901),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1055),
.B(n_979),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_R g1112 ( 
.A(n_1066),
.B(n_955),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_R g1113 ( 
.A(n_1066),
.B(n_955),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1014),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_R g1115 ( 
.A(n_1011),
.B(n_880),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_1050),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1014),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1031),
.B(n_939),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_1057),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1016),
.Y(n_1120)
);

NAND2xp33_ASAP7_75t_R g1121 ( 
.A(n_1048),
.B(n_917),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1031),
.B(n_944),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_1001),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_1073),
.B(n_972),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1001),
.Y(n_1125)
);

NAND2xp33_ASAP7_75t_R g1126 ( 
.A(n_1048),
.B(n_917),
.Y(n_1126)
);

XOR2xp5_ASAP7_75t_L g1127 ( 
.A(n_1021),
.B(n_914),
.Y(n_1127)
);

INVx8_ASAP7_75t_L g1128 ( 
.A(n_1023),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1042),
.B(n_900),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_985),
.B(n_936),
.Y(n_1130)
);

OR2x2_ASAP7_75t_L g1131 ( 
.A(n_1016),
.B(n_985),
.Y(n_1131)
);

NAND2xp33_ASAP7_75t_R g1132 ( 
.A(n_1054),
.B(n_917),
.Y(n_1132)
);

OR2x6_ASAP7_75t_L g1133 ( 
.A(n_1073),
.B(n_972),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_990),
.B(n_880),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_R g1135 ( 
.A(n_1054),
.B(n_947),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_1050),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_R g1137 ( 
.A(n_1011),
.B(n_982),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1023),
.B(n_927),
.Y(n_1138)
);

XOR2xp5_ASAP7_75t_L g1139 ( 
.A(n_1070),
.B(n_894),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_R g1140 ( 
.A(n_1070),
.B(n_983),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_990),
.B(n_1031),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1107),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1141),
.B(n_991),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1105),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1080),
.Y(n_1145)
);

OR2x6_ASAP7_75t_SL g1146 ( 
.A(n_1109),
.B(n_986),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1105),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1114),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1117),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1120),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1086),
.Y(n_1151)
);

NOR2x1_ASAP7_75t_L g1152 ( 
.A(n_1103),
.B(n_1023),
.Y(n_1152)
);

OR2x2_ASAP7_75t_SL g1153 ( 
.A(n_1109),
.B(n_1054),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1124),
.A2(n_983),
.B1(n_977),
.B2(n_991),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_1082),
.B(n_1058),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1100),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1131),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1124),
.A2(n_977),
.B1(n_1039),
.B2(n_1035),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1138),
.B(n_993),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1123),
.B(n_993),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1138),
.B(n_993),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_1121),
.Y(n_1162)
);

NAND2xp33_ASAP7_75t_SL g1163 ( 
.A(n_1140),
.B(n_1031),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1098),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1106),
.B(n_66),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1138),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1094),
.B(n_66),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1125),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1128),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1095),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1110),
.B(n_993),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1128),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1083),
.B(n_986),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1128),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1085),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1088),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1103),
.B(n_987),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1088),
.B(n_987),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1130),
.A2(n_1061),
.B1(n_1049),
.B2(n_942),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1124),
.A2(n_1061),
.B1(n_971),
.B2(n_957),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1084),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1091),
.Y(n_1182)
);

BUFx3_ASAP7_75t_R g1183 ( 
.A(n_1079),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1111),
.B(n_1052),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1139),
.A2(n_938),
.B1(n_928),
.B2(n_954),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1091),
.B(n_992),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1087),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1129),
.B(n_1052),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1130),
.A2(n_1049),
.B1(n_1054),
.B2(n_1058),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1087),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1093),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1093),
.B(n_1023),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1089),
.B(n_1056),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1158),
.A2(n_1133),
.B1(n_1094),
.B2(n_1127),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1170),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1151),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1144),
.Y(n_1197)
);

AOI221x1_ASAP7_75t_SL g1198 ( 
.A1(n_1167),
.A2(n_1076),
.B1(n_1092),
.B2(n_1122),
.C(n_1089),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1168),
.B(n_1108),
.Y(n_1199)
);

NAND5xp2_ASAP7_75t_SL g1200 ( 
.A(n_1154),
.B(n_910),
.C(n_1077),
.D(n_981),
.E(n_928),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1181),
.Y(n_1201)
);

INVx5_ASAP7_75t_SL g1202 ( 
.A(n_1192),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1170),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1143),
.B(n_1134),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1168),
.B(n_1119),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1181),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1144),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1170),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1145),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1182),
.B(n_1099),
.Y(n_1210)
);

OAI31xp33_ASAP7_75t_L g1211 ( 
.A1(n_1185),
.A2(n_1162),
.A3(n_1180),
.B(n_1165),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1147),
.Y(n_1212)
);

NOR2xp67_ASAP7_75t_L g1213 ( 
.A(n_1162),
.B(n_1090),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1143),
.B(n_1116),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1151),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1184),
.B(n_1136),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1184),
.B(n_1092),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1193),
.B(n_1118),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1192),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1182),
.Y(n_1220)
);

AOI221xp5_ASAP7_75t_L g1221 ( 
.A1(n_1185),
.A2(n_903),
.B1(n_978),
.B2(n_889),
.C(n_931),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1176),
.B(n_1118),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1151),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1147),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1142),
.Y(n_1225)
);

AOI33xp33_ASAP7_75t_L g1226 ( 
.A1(n_1179),
.A2(n_1122),
.A3(n_1102),
.B1(n_1135),
.B2(n_1047),
.B3(n_1046),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1193),
.B(n_1056),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1142),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1157),
.B(n_995),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1175),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1192),
.Y(n_1231)
);

BUFx5_ASAP7_75t_L g1232 ( 
.A(n_1159),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1159),
.B(n_1133),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1179),
.A2(n_1133),
.B1(n_1049),
.B2(n_1101),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1159),
.B(n_1023),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1188),
.B(n_1062),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1157),
.B(n_995),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1148),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1176),
.B(n_992),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1188),
.B(n_1062),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1176),
.B(n_996),
.Y(n_1241)
);

AOI211xp5_ASAP7_75t_L g1242 ( 
.A1(n_1186),
.A2(n_1097),
.B(n_1137),
.C(n_1115),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1171),
.B(n_1038),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1148),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1145),
.B(n_996),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1149),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1146),
.A2(n_1030),
.B1(n_1081),
.B2(n_1078),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1173),
.B(n_995),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_SL g1249 ( 
.A1(n_1153),
.A2(n_1030),
.B1(n_1104),
.B2(n_1113),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1220),
.B(n_1153),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1236),
.B(n_1146),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1209),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1229),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1197),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1236),
.B(n_1146),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1240),
.B(n_1171),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1240),
.B(n_1160),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1229),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1237),
.Y(n_1259)
);

AOI21xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1206),
.A2(n_1096),
.B(n_1173),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1207),
.B(n_1178),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1237),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1248),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1230),
.B(n_1186),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1196),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1248),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1232),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1227),
.B(n_1160),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1212),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1224),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1219),
.B(n_1159),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1233),
.B(n_1152),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1232),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1199),
.B(n_1210),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1225),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1245),
.B(n_1178),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1227),
.B(n_1152),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1204),
.B(n_1166),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1196),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1204),
.B(n_1166),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1243),
.B(n_1166),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1232),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1252),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1276),
.B(n_1228),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1271),
.B(n_1213),
.Y(n_1285)
);

AO221x2_ASAP7_75t_L g1286 ( 
.A1(n_1267),
.A2(n_1247),
.B1(n_1249),
.B2(n_1198),
.C(n_1206),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1252),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1276),
.B(n_1230),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1250),
.A2(n_1194),
.B1(n_1234),
.B2(n_1242),
.Y(n_1289)
);

NAND2xp33_ASAP7_75t_SL g1290 ( 
.A(n_1250),
.B(n_1195),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1251),
.A2(n_1126),
.B1(n_1221),
.B2(n_1132),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1274),
.B(n_1199),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1264),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1264),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1274),
.B(n_1205),
.Y(n_1295)
);

AO221x2_ASAP7_75t_L g1296 ( 
.A1(n_1267),
.A2(n_1211),
.B1(n_1201),
.B2(n_1226),
.C(n_1183),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1274),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1251),
.A2(n_1233),
.B1(n_1235),
.B2(n_1177),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1250),
.Y(n_1299)
);

AO221x2_ASAP7_75t_L g1300 ( 
.A1(n_1267),
.A2(n_1226),
.B1(n_1200),
.B2(n_1163),
.C(n_1195),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1254),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1260),
.A2(n_1222),
.B1(n_1190),
.B2(n_1177),
.Y(n_1302)
);

AO221x2_ASAP7_75t_L g1303 ( 
.A1(n_1267),
.A2(n_1195),
.B1(n_1208),
.B2(n_1232),
.C(n_1203),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1251),
.B(n_1214),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1255),
.B(n_1214),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1254),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_1261),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1261),
.B(n_1243),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1255),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1255),
.B(n_1216),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1256),
.B(n_1218),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1271),
.B(n_1219),
.Y(n_1312)
);

INVxp33_ASAP7_75t_SL g1313 ( 
.A(n_1256),
.Y(n_1313)
);

AO221x2_ASAP7_75t_L g1314 ( 
.A1(n_1282),
.A2(n_1232),
.B1(n_1203),
.B2(n_1191),
.C(n_1101),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1293),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1309),
.B(n_1271),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1303),
.B(n_1256),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1303),
.B(n_1268),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1306),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1297),
.B(n_1269),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1293),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1294),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1303),
.B(n_1268),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1304),
.B(n_1268),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1306),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1292),
.B(n_1269),
.Y(n_1326)
);

NOR2x1_ASAP7_75t_L g1327 ( 
.A(n_1294),
.B(n_1270),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1307),
.B(n_1270),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1305),
.B(n_1257),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1287),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1288),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1311),
.B(n_1257),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1313),
.B(n_1277),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1284),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1295),
.B(n_1275),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1314),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1285),
.B(n_1257),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1299),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1300),
.B(n_1275),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1296),
.A2(n_1189),
.B1(n_1258),
.B2(n_1253),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1285),
.B(n_1273),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1299),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1283),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1313),
.B(n_1283),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1308),
.B(n_1263),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1300),
.B(n_1277),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1301),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1301),
.Y(n_1348)
);

AOI222xp33_ASAP7_75t_L g1349 ( 
.A1(n_1340),
.A2(n_1289),
.B1(n_1296),
.B2(n_1302),
.C1(n_1286),
.C2(n_1300),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1338),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1315),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1315),
.B(n_1312),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1321),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1338),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1346),
.A2(n_1296),
.B1(n_1286),
.B2(n_1291),
.Y(n_1355)
);

AOI322xp5_ASAP7_75t_L g1356 ( 
.A1(n_1339),
.A2(n_1302),
.A3(n_1317),
.B1(n_1318),
.B2(n_1323),
.C1(n_1322),
.C2(n_1327),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1336),
.A2(n_1286),
.B1(n_1331),
.B2(n_1333),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_SL g1358 ( 
.A(n_1330),
.B(n_1290),
.C(n_1260),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1316),
.Y(n_1359)
);

AOI332xp33_ASAP7_75t_L g1360 ( 
.A1(n_1342),
.A2(n_1285),
.A3(n_1312),
.B1(n_1298),
.B2(n_1310),
.B3(n_1263),
.C1(n_1266),
.C2(n_1259),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1342),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1319),
.Y(n_1362)
);

OAI221xp5_ASAP7_75t_L g1363 ( 
.A1(n_1336),
.A2(n_1290),
.B1(n_1259),
.B2(n_1262),
.C(n_1189),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1327),
.A2(n_1277),
.B(n_1030),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_SL g1365 ( 
.A(n_1330),
.B(n_1282),
.C(n_1112),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1334),
.B(n_1278),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1336),
.A2(n_1314),
.B1(n_1262),
.B2(n_1266),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1324),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1336),
.A2(n_1312),
.B1(n_1273),
.B2(n_1271),
.Y(n_1369)
);

OAI21xp33_ASAP7_75t_L g1370 ( 
.A1(n_1317),
.A2(n_1273),
.B(n_1282),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1347),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1318),
.A2(n_1271),
.B1(n_1272),
.B2(n_1219),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1335),
.B(n_1314),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1323),
.A2(n_1253),
.B1(n_1258),
.B2(n_1272),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1319),
.A2(n_1282),
.B(n_1253),
.C(n_1258),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1335),
.A2(n_1272),
.B1(n_1231),
.B2(n_1191),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1325),
.Y(n_1377)
);

NOR2xp67_ASAP7_75t_L g1378 ( 
.A(n_1316),
.B(n_1343),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1324),
.B(n_1218),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1325),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1362),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1349),
.A2(n_1334),
.B1(n_1337),
.B2(n_1316),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1352),
.B(n_1329),
.Y(n_1383)
);

NAND2x1_ASAP7_75t_SL g1384 ( 
.A(n_1357),
.B(n_1355),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1353),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1377),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1380),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1351),
.B(n_1329),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1359),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1350),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1371),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1379),
.B(n_1337),
.Y(n_1392)
);

AOI222xp33_ASAP7_75t_L g1393 ( 
.A1(n_1363),
.A2(n_1328),
.B1(n_1320),
.B2(n_1344),
.C1(n_1348),
.C2(n_1343),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1371),
.B(n_1348),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1368),
.B(n_1332),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1354),
.B(n_1332),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1361),
.B(n_1326),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1356),
.B(n_1326),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1349),
.B(n_1316),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1373),
.B(n_1343),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1367),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1366),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1378),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1375),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1374),
.B(n_1343),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1364),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1364),
.B(n_1345),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1369),
.B(n_1341),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1358),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1372),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1365),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_L g1412 ( 
.A(n_1370),
.B(n_1341),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1391),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1385),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1384),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1381),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1381),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1386),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1385),
.B(n_1345),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1386),
.Y(n_1420)
);

CKINVDCx6p67_ASAP7_75t_R g1421 ( 
.A(n_1394),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1387),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1384),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1387),
.Y(n_1424)
);

CKINVDCx6p67_ASAP7_75t_R g1425 ( 
.A(n_1400),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1390),
.Y(n_1426)
);

CKINVDCx16_ASAP7_75t_R g1427 ( 
.A(n_1409),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1383),
.B(n_1376),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1409),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1399),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1383),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1390),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1389),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1389),
.Y(n_1434)
);

INVxp33_ASAP7_75t_SL g1435 ( 
.A(n_1401),
.Y(n_1435)
);

INVxp33_ASAP7_75t_SL g1436 ( 
.A(n_1401),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1388),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1396),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1397),
.Y(n_1439)
);

INVxp67_ASAP7_75t_SL g1440 ( 
.A(n_1411),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1395),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1392),
.B(n_1216),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1395),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1402),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1405),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1398),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1404),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1392),
.Y(n_1448)
);

INVxp33_ASAP7_75t_SL g1449 ( 
.A(n_1382),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1404),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1415),
.B(n_1393),
.C(n_1403),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1427),
.B(n_1410),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1421),
.B(n_1410),
.Y(n_1453)
);

NAND5xp2_ASAP7_75t_L g1454 ( 
.A(n_1448),
.B(n_1405),
.C(n_1360),
.D(n_1408),
.E(n_1406),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1415),
.B(n_1406),
.C(n_1407),
.Y(n_1455)
);

AOI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1446),
.A2(n_1412),
.B1(n_1408),
.B2(n_1281),
.C(n_1238),
.Y(n_1456)
);

OAI21xp33_ASAP7_75t_L g1457 ( 
.A1(n_1440),
.A2(n_1281),
.B(n_1280),
.Y(n_1457)
);

O2A1O1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1423),
.A2(n_1030),
.B(n_1280),
.C(n_1278),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1443),
.Y(n_1459)
);

NOR3xp33_ASAP7_75t_L g1460 ( 
.A(n_1423),
.B(n_1239),
.C(n_1241),
.Y(n_1460)
);

NOR2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1431),
.B(n_1233),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1443),
.Y(n_1462)
);

NOR3xp33_ASAP7_75t_L g1463 ( 
.A(n_1429),
.B(n_1065),
.C(n_1244),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1430),
.B(n_1030),
.C(n_1155),
.Y(n_1464)
);

OAI211xp5_ASAP7_75t_L g1465 ( 
.A1(n_1414),
.A2(n_1155),
.B(n_878),
.C(n_1278),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1429),
.B(n_1232),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1431),
.B(n_1280),
.Y(n_1467)
);

NAND4xp25_ASAP7_75t_SL g1468 ( 
.A(n_1428),
.B(n_1281),
.C(n_1217),
.D(n_1190),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1450),
.B(n_1246),
.C(n_1046),
.Y(n_1469)
);

NAND3x1_ASAP7_75t_L g1470 ( 
.A(n_1413),
.B(n_1217),
.C(n_1172),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1434),
.B(n_1232),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1434),
.B(n_1265),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1433),
.Y(n_1473)
);

NAND2x1_ASAP7_75t_L g1474 ( 
.A(n_1433),
.B(n_1231),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1441),
.Y(n_1475)
);

OAI211xp5_ASAP7_75t_L g1476 ( 
.A1(n_1444),
.A2(n_1002),
.B(n_1231),
.C(n_1047),
.Y(n_1476)
);

NAND3xp33_ASAP7_75t_SL g1477 ( 
.A(n_1447),
.B(n_1450),
.C(n_1419),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1447),
.B(n_1043),
.C(n_1038),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1420),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1445),
.B(n_1043),
.C(n_1235),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1421),
.B(n_1265),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_SL g1482 ( 
.A(n_1439),
.B(n_1272),
.C(n_1002),
.Y(n_1482)
);

NOR4xp25_ASAP7_75t_L g1483 ( 
.A(n_1420),
.B(n_1279),
.C(n_1265),
.D(n_884),
.Y(n_1483)
);

AOI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1449),
.A2(n_1279),
.B1(n_1058),
.B2(n_1028),
.C(n_1026),
.Y(n_1484)
);

NOR3xp33_ASAP7_75t_L g1485 ( 
.A(n_1445),
.B(n_1065),
.C(n_927),
.Y(n_1485)
);

NAND5xp2_ASAP7_75t_L g1486 ( 
.A(n_1449),
.B(n_1435),
.C(n_1436),
.D(n_1438),
.E(n_1426),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1486),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1473),
.Y(n_1488)
);

NAND4xp25_ASAP7_75t_SL g1489 ( 
.A(n_1456),
.B(n_1422),
.C(n_1424),
.D(n_1418),
.Y(n_1489)
);

AOI221xp5_ASAP7_75t_SL g1490 ( 
.A1(n_1454),
.A2(n_1435),
.B1(n_1436),
.B2(n_1416),
.C(n_1432),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1455),
.B(n_1437),
.C(n_1422),
.Y(n_1491)
);

NOR3xp33_ASAP7_75t_L g1492 ( 
.A(n_1486),
.B(n_1417),
.C(n_1424),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1451),
.A2(n_1425),
.B1(n_1442),
.B2(n_1202),
.Y(n_1493)
);

AOI32xp33_ASAP7_75t_L g1494 ( 
.A1(n_1453),
.A2(n_1442),
.A3(n_1425),
.B1(n_1068),
.B2(n_1067),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1477),
.A2(n_1279),
.B1(n_1235),
.B2(n_1192),
.Y(n_1495)
);

AND4x2_ASAP7_75t_L g1496 ( 
.A(n_1470),
.B(n_886),
.C(n_1202),
.D(n_1231),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1452),
.A2(n_1026),
.B1(n_1028),
.B2(n_1022),
.C(n_1017),
.Y(n_1497)
);

NOR3xp33_ASAP7_75t_L g1498 ( 
.A(n_1459),
.B(n_933),
.C(n_905),
.Y(n_1498)
);

AOI21xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1462),
.A2(n_1172),
.B(n_969),
.Y(n_1499)
);

OAI321xp33_ASAP7_75t_L g1500 ( 
.A1(n_1475),
.A2(n_1017),
.A3(n_1022),
.B1(n_1169),
.B2(n_1174),
.C(n_1149),
.Y(n_1500)
);

AOI222xp33_ASAP7_75t_L g1501 ( 
.A1(n_1484),
.A2(n_1029),
.B1(n_1024),
.B2(n_1150),
.C1(n_1020),
.C2(n_1223),
.Y(n_1501)
);

AOI311xp33_ASAP7_75t_L g1502 ( 
.A1(n_1479),
.A2(n_1068),
.A3(n_1074),
.B(n_1069),
.C(n_1067),
.Y(n_1502)
);

OAI211xp5_ASAP7_75t_L g1503 ( 
.A1(n_1466),
.A2(n_1069),
.B(n_1074),
.C(n_1172),
.Y(n_1503)
);

OAI211xp5_ASAP7_75t_SL g1504 ( 
.A1(n_1481),
.A2(n_1034),
.B(n_1172),
.C(n_1187),
.Y(n_1504)
);

OAI211xp5_ASAP7_75t_SL g1505 ( 
.A1(n_1471),
.A2(n_1034),
.B(n_1187),
.C(n_1169),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1467),
.B(n_1187),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1472),
.A2(n_969),
.B(n_1161),
.Y(n_1507)
);

AOI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1463),
.A2(n_1024),
.B1(n_1029),
.B2(n_1150),
.C(n_1034),
.Y(n_1508)
);

OAI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1474),
.A2(n_1223),
.B1(n_1215),
.B2(n_1156),
.C(n_1164),
.Y(n_1509)
);

AOI222xp33_ASAP7_75t_L g1510 ( 
.A1(n_1469),
.A2(n_1020),
.B1(n_1215),
.B2(n_1164),
.C1(n_1156),
.C2(n_1071),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1457),
.A2(n_1202),
.B1(n_1161),
.B2(n_1169),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1461),
.B(n_1202),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1468),
.B(n_1161),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_R g1514 ( 
.A(n_1482),
.B(n_78),
.Y(n_1514)
);

NOR3xp33_ASAP7_75t_L g1515 ( 
.A(n_1464),
.B(n_933),
.C(n_905),
.Y(n_1515)
);

OAI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1483),
.A2(n_1174),
.B1(n_1008),
.B2(n_1034),
.C(n_1036),
.Y(n_1516)
);

AOI221x1_ASAP7_75t_L g1517 ( 
.A1(n_1460),
.A2(n_1478),
.B1(n_1480),
.B2(n_1485),
.C(n_1465),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1487),
.B(n_1492),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1488),
.Y(n_1519)
);

NAND4xp75_ASAP7_75t_L g1520 ( 
.A(n_1490),
.B(n_1458),
.C(n_1476),
.D(n_934),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1506),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1491),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1489),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1512),
.B(n_1161),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1494),
.B(n_969),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1493),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1495),
.A2(n_1513),
.B1(n_1508),
.B2(n_1515),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1517),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_L g1529 ( 
.A(n_1503),
.B(n_1174),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1496),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1502),
.B(n_1019),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1516),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1504),
.B(n_79),
.Y(n_1533)
);

XNOR2xp5_ASAP7_75t_L g1534 ( 
.A(n_1511),
.B(n_1497),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1507),
.A2(n_1036),
.B1(n_1040),
.B2(n_1041),
.Y(n_1535)
);

NOR2x1_ASAP7_75t_L g1536 ( 
.A(n_1505),
.B(n_83),
.Y(n_1536)
);

NAND4xp75_ASAP7_75t_L g1537 ( 
.A(n_1514),
.B(n_1006),
.C(n_1072),
.D(n_1053),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1499),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1509),
.B(n_1019),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1510),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1497),
.B(n_160),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1501),
.A2(n_1040),
.B1(n_1041),
.B2(n_1044),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1498),
.Y(n_1543)
);

AND4x1_ASAP7_75t_L g1544 ( 
.A(n_1518),
.B(n_1500),
.C(n_169),
.D(n_170),
.Y(n_1544)
);

NOR3xp33_ASAP7_75t_SL g1545 ( 
.A(n_1523),
.B(n_161),
.C(n_177),
.Y(n_1545)
);

NAND2xp33_ASAP7_75t_SL g1546 ( 
.A(n_1522),
.B(n_1530),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_SL g1547 ( 
.A(n_1519),
.B(n_1008),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_R g1548 ( 
.A(n_1526),
.B(n_1528),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1521),
.B(n_178),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1538),
.B(n_1045),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1543),
.B(n_180),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1532),
.B(n_222),
.Y(n_1552)
);

NAND2xp33_ASAP7_75t_SL g1553 ( 
.A(n_1534),
.B(n_1531),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1533),
.B(n_1045),
.Y(n_1554)
);

AND3x1_ASAP7_75t_L g1555 ( 
.A(n_1527),
.B(n_1540),
.C(n_1536),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_R g1556 ( 
.A(n_1541),
.B(n_946),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1536),
.B(n_1072),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_R g1558 ( 
.A(n_1524),
.B(n_946),
.Y(n_1558)
);

NAND2xp33_ASAP7_75t_SL g1559 ( 
.A(n_1525),
.B(n_1071),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_R g1560 ( 
.A(n_1524),
.B(n_895),
.Y(n_1560)
);

XNOR2xp5_ASAP7_75t_L g1561 ( 
.A(n_1520),
.B(n_943),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_R g1562 ( 
.A(n_1539),
.B(n_895),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1529),
.B(n_1006),
.C(n_1053),
.Y(n_1563)
);

NAND2xp33_ASAP7_75t_SL g1564 ( 
.A(n_1537),
.B(n_1529),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1535),
.B(n_1006),
.C(n_1044),
.Y(n_1565)
);

NOR3xp33_ASAP7_75t_SL g1566 ( 
.A(n_1542),
.B(n_967),
.C(n_892),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1564),
.A2(n_1006),
.B1(n_967),
.B2(n_943),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1553),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1555),
.A2(n_966),
.B1(n_892),
.B2(n_994),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1548),
.Y(n_1570)
);

AOI32xp33_ASAP7_75t_L g1571 ( 
.A1(n_1546),
.A2(n_994),
.A3(n_879),
.B1(n_1005),
.B2(n_1003),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1545),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1551),
.B(n_1005),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1552),
.B(n_879),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1544),
.B(n_883),
.Y(n_1575)
);

NOR3xp33_ASAP7_75t_SL g1576 ( 
.A(n_1550),
.B(n_1004),
.C(n_1003),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1554),
.A2(n_998),
.B(n_1004),
.C(n_1000),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_R g1578 ( 
.A(n_1556),
.B(n_876),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1570),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1568),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1572),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1573),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1577),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1574),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1579),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1579),
.A2(n_1571),
.B1(n_1561),
.B2(n_1563),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_SL g1587 ( 
.A1(n_1580),
.A2(n_1549),
.B1(n_1574),
.B2(n_1575),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1581),
.A2(n_1557),
.B1(n_1576),
.B2(n_1565),
.Y(n_1588)
);

AOI31xp33_ASAP7_75t_L g1589 ( 
.A1(n_1587),
.A2(n_1584),
.A3(n_1582),
.B(n_1583),
.Y(n_1589)
);

AOI31xp33_ASAP7_75t_L g1590 ( 
.A1(n_1586),
.A2(n_1578),
.A3(n_1559),
.B(n_1569),
.Y(n_1590)
);

AOI31xp33_ASAP7_75t_L g1591 ( 
.A1(n_1585),
.A2(n_1547),
.A3(n_1562),
.B(n_1567),
.Y(n_1591)
);

AOI31xp33_ASAP7_75t_L g1592 ( 
.A1(n_1588),
.A2(n_1558),
.A3(n_1560),
.B(n_1566),
.Y(n_1592)
);

O2A1O1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1589),
.A2(n_998),
.B(n_1000),
.C(n_988),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1592),
.B(n_984),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1593),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1594),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1596),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1597),
.A2(n_1590),
.B1(n_1595),
.B2(n_1591),
.C(n_999),
.Y(n_1598)
);

AOI211xp5_ASAP7_75t_L g1599 ( 
.A1(n_1598),
.A2(n_876),
.B(n_999),
.C(n_988),
.Y(n_1599)
);


endmodule