module fake_jpeg_1839_n_69 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_69);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

BUFx10_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_8),
.B(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_10),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_11),
.A2(n_0),
.B1(n_5),
.B2(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_26),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_16),
.B1(n_14),
.B2(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_34),
.B1(n_35),
.B2(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_17),
.B1(n_19),
.B2(n_9),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_9),
.B1(n_25),
.B2(n_20),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_23),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_20),
.C(n_26),
.Y(n_39)
);

AND2x6_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_22),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_9),
.B(n_28),
.C(n_24),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_43),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_31),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_24),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_30),
.B(n_34),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_32),
.B1(n_49),
.B2(n_50),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_53),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_32),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_32),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_61),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_54),
.C(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_57),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_65),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);


endmodule