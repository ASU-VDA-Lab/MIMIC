module fake_aes_3926_n_362 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_362);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_362;
wire n_117;
wire n_361;
wire n_185;
wire n_284;
wire n_278;
wire n_114;
wire n_125;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_296;
wire n_157;
wire n_202;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_163;
wire n_227;
wire n_231;
wire n_298;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_150;
wire n_301;
wire n_222;
wire n_234;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_167;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_241;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_247;
wire n_304;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_235;
wire n_243;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_153;
wire n_259;
wire n_308;
wire n_140;
wire n_207;
wire n_224;
wire n_219;
wire n_133;
wire n_149;
wire n_214;
wire n_204;
wire n_254;
wire n_262;
wire n_239;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_342;
wire n_217;
wire n_139;
wire n_193;
wire n_273;
wire n_120;
wire n_245;
wire n_357;
wire n_260;
wire n_197;
wire n_201;
wire n_317;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_179;
wire n_315;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_344;
wire n_136;
wire n_283;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_168;
wire n_134;
wire n_233;
wire n_173;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_115;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_359;
wire n_346;
wire n_180;
wire n_335;
wire n_272;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_188;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_138;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_355;
wire n_226;
wire n_159;
wire n_337;
wire n_176;
wire n_123;
wire n_223;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_332;
wire n_350;
wire n_164;
wire n_175;
wire n_145;
wire n_290;
wire n_280;
wire n_109;
wire n_132;
wire n_151;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_12), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_82), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_50), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_17), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_16), .Y(n_112) );
BUFx5_ASAP7_75t_L g113 ( .A(n_93), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_62), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_11), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_88), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_23), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_54), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_85), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_91), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_57), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_60), .Y(n_122) );
BUFx5_ASAP7_75t_L g123 ( .A(n_97), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_106), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_87), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_76), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_72), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_1), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_92), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_19), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_46), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_104), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_35), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_105), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_33), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_29), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_53), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_43), .Y(n_142) );
BUFx10_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_15), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_95), .Y(n_145) );
CKINVDCx14_ASAP7_75t_R g146 ( .A(n_74), .Y(n_146) );
BUFx2_ASAP7_75t_L g147 ( .A(n_98), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_3), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_75), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_55), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_48), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_103), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_38), .Y(n_154) );
CKINVDCx14_ASAP7_75t_R g155 ( .A(n_100), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_2), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_8), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_80), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_21), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_58), .Y(n_160) );
INVxp33_ASAP7_75t_L g161 ( .A(n_52), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_69), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_78), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_90), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_77), .Y(n_166) );
BUFx5_ASAP7_75t_L g167 ( .A(n_101), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_25), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_51), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_30), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_59), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_32), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_40), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_102), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_94), .Y(n_175) );
NOR2xp67_ASAP7_75t_L g176 ( .A(n_34), .B(n_6), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_9), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_107), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_96), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_109), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_147), .B(n_0), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_134), .B(n_0), .Y(n_182) );
OAI22xp5_ASAP7_75t_SL g183 ( .A1(n_128), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_113), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_116), .B(n_4), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_117), .B(n_4), .Y(n_187) );
INVx5_ASAP7_75t_L g188 ( .A(n_143), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_148), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_108), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_110), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_113), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_112), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_132), .B(n_5), .Y(n_194) );
INVx5_ASAP7_75t_L g195 ( .A(n_119), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_114), .Y(n_196) );
OAI22xp5_ASAP7_75t_SL g197 ( .A1(n_115), .A2(n_7), .B1(n_10), .B2(n_13), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_161), .B(n_14), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_184), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_188), .B(n_146), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_192), .Y(n_201) );
BUFx6f_ASAP7_75t_SL g202 ( .A(n_181), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_196), .B(n_155), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_180), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_180), .Y(n_205) );
NAND2xp33_ASAP7_75t_SL g206 ( .A(n_198), .B(n_120), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_191), .B(n_111), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_185), .B(n_162), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_186), .Y(n_209) );
AND2x6_ASAP7_75t_L g210 ( .A(n_182), .B(n_118), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_209), .B(n_187), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_200), .B(n_189), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_199), .Y(n_213) );
INVx8_ASAP7_75t_L g214 ( .A(n_202), .Y(n_214) );
OAI221xp5_ASAP7_75t_L g215 ( .A1(n_204), .A2(n_194), .B1(n_183), .B2(n_197), .C(n_176), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_205), .B(n_124), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_207), .B(n_126), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_201), .Y(n_218) );
NOR3xp33_ASAP7_75t_L g219 ( .A(n_206), .B(n_193), .C(n_122), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_210), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_203), .B(n_127), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_210), .B(n_129), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_208), .Y(n_223) );
INVx1_ASAP7_75t_SL g224 ( .A(n_214), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_218), .A2(n_223), .B(n_213), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_216), .A2(n_217), .B(n_221), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_220), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_212), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_214), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_212), .A2(n_190), .B1(n_153), .B2(n_152), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_222), .A2(n_125), .B(n_121), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_219), .B(n_130), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_215), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_211), .A2(n_133), .B(n_131), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_211), .A2(n_137), .B(n_136), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_224), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_228), .B(n_138), .Y(n_237) );
O2A1O1Ixp5_ASAP7_75t_L g238 ( .A1(n_231), .A2(n_170), .B(n_175), .C(n_144), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_229), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_226), .A2(n_145), .B(n_142), .Y(n_240) );
INVxp67_ASAP7_75t_L g241 ( .A(n_230), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_232), .B(n_135), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_227), .Y(n_243) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_225), .A2(n_150), .B(n_149), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_234), .Y(n_245) );
AO31x2_ASAP7_75t_L g246 ( .A1(n_235), .A2(n_166), .A3(n_179), .B(n_178), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_233), .B(n_157), .Y(n_247) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_227), .A2(n_165), .A3(n_177), .B(n_173), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_239), .Y(n_249) );
AOI21x1_ASAP7_75t_L g250 ( .A1(n_244), .A2(n_160), .B(n_159), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_243), .Y(n_251) );
AOI21x1_ASAP7_75t_L g252 ( .A1(n_240), .A2(n_164), .B(n_163), .Y(n_252) );
BUFx4_ASAP7_75t_SL g253 ( .A(n_236), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_242), .B(n_139), .Y(n_254) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_238), .A2(n_172), .B(n_168), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_237), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_237), .B(n_141), .Y(n_257) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_247), .A2(n_167), .B(n_123), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_248), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_246), .B(n_140), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_248), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_246), .Y(n_262) );
INVxp67_ASAP7_75t_SL g263 ( .A(n_236), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_245), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_241), .B(n_151), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_SL g266 ( .A1(n_240), .A2(n_18), .B(n_20), .C(n_22), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_245), .Y(n_267) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_261), .A2(n_24), .A3(n_26), .B(n_27), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_263), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_259), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_264), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_267), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_267), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_262), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_256), .B(n_154), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_257), .Y(n_276) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_258), .A2(n_169), .B(n_158), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_254), .Y(n_278) );
OAI21x1_ASAP7_75t_SL g279 ( .A1(n_252), .A2(n_28), .B(n_31), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_260), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_265), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_250), .Y(n_282) );
AOI21x1_ASAP7_75t_L g283 ( .A1(n_255), .A2(n_195), .B(n_36), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_266), .Y(n_284) );
INVx2_ASAP7_75t_SL g285 ( .A(n_253), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_251), .Y(n_286) );
AO31x2_ASAP7_75t_L g287 ( .A1(n_261), .A2(n_37), .A3(n_39), .B(n_41), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_249), .B(n_42), .Y(n_288) );
OA21x2_ASAP7_75t_L g289 ( .A1(n_261), .A2(n_174), .B(n_171), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_251), .Y(n_290) );
BUFx12f_ASAP7_75t_L g291 ( .A(n_256), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_251), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_259), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_269), .B(n_44), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_281), .B(n_45), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_272), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_286), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_278), .B(n_47), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_271), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_280), .B(n_273), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_285), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_290), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_292), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_288), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_276), .B(n_49), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_291), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_288), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_270), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_274), .B(n_56), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_293), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_268), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_268), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_289), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_275), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_287), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_283), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_300), .B(n_277), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_296), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_303), .B(n_297), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_301), .B(n_61), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_302), .B(n_284), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_306), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_311), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_311), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_304), .B(n_63), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_307), .B(n_64), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_315), .B(n_65), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_295), .B(n_66), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_308), .Y(n_332) );
INVx5_ASAP7_75t_L g333 ( .A(n_309), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_325), .B(n_310), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_321), .B(n_317), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_320), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_326), .B(n_314), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_324), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_327), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_332), .B(n_294), .Y(n_340) );
AND2x4_ASAP7_75t_SL g341 ( .A(n_338), .B(n_330), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_335), .B(n_319), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_336), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_341), .Y(n_344) );
AOI322xp5_ASAP7_75t_L g345 ( .A1(n_342), .A2(n_340), .A3(n_339), .B1(n_337), .B2(n_334), .C1(n_322), .C2(n_305), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_343), .B(n_337), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_346), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_344), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_347), .B(n_345), .Y(n_349) );
OAI211xp5_ASAP7_75t_L g350 ( .A1(n_348), .A2(n_333), .B(n_331), .C(n_298), .Y(n_350) );
NOR3xp33_ASAP7_75t_L g351 ( .A(n_349), .B(n_350), .C(n_328), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_351), .B(n_323), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_352), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_353), .Y(n_354) );
XNOR2xp5_ASAP7_75t_L g355 ( .A(n_354), .B(n_329), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_355), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_356), .Y(n_357) );
OAI22xp33_ASAP7_75t_SL g358 ( .A1(n_357), .A2(n_316), .B1(n_313), .B2(n_312), .Y(n_358) );
AO21x2_ASAP7_75t_L g359 ( .A1(n_358), .A2(n_318), .B(n_68), .Y(n_359) );
AO21x2_ASAP7_75t_L g360 ( .A1(n_359), .A2(n_67), .B(n_70), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_360), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_361), .A2(n_71), .B(n_73), .Y(n_362) );
endmodule