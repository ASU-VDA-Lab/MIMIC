module fake_netlist_6_2386_n_2055 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2055);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2055;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_527;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_18),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_68),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_66),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_127),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_183),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_128),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_66),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_26),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_39),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_34),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_56),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_59),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_13),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_65),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_90),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_123),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_180),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_85),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_176),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_135),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_16),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_73),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_7),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_57),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_48),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_25),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_100),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_167),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_151),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_124),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_134),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_163),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_62),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_26),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_103),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_114),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_88),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_155),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_70),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_98),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_24),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_121),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_14),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_156),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_149),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_105),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_185),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_8),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_13),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_173),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_12),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_111),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_148),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_1),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_143),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_129),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_19),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_83),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_174),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_166),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_43),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_56),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_57),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_33),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_48),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_95),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_104),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_186),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_164),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_81),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_35),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_197),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_53),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_3),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_73),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_182),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_31),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_15),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_15),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_29),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_31),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_21),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_122),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_147),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_21),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_136),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_177),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_133),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_106),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_50),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_68),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_50),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_30),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_161),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_132),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_158),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_51),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_22),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_196),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_6),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_87),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_94),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_86),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_140),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_102),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_113),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_71),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_71),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_4),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_63),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_198),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_65),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_33),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_58),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_92),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_52),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_131),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_96),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_144),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_54),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_34),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_60),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_77),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_44),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_54),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_125),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_62),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_190),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_175),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_42),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_142),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_168),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_72),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_160),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_51),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_138),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_72),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_116),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_43),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_38),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_32),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_39),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_64),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_35),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_141),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_82),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_47),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_3),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_145),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_14),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_6),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_170),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_76),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_172),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_40),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_59),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_41),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_184),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_195),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_9),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_109),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_99),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_165),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_23),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_146),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_150),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_194),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_58),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_70),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_37),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_154),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_20),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_25),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_47),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_18),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_171),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_192),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_38),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_130),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_157),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_4),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_46),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_11),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_55),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_28),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_41),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_74),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_79),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_75),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_307),
.B(n_0),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_260),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_209),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_327),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_199),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_200),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_219),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_260),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_327),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_231),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_311),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_327),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_201),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_202),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_207),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_208),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_217),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_211),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_202),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_223),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_223),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_256),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_223),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_282),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_223),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_223),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_270),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_270),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_270),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_212),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_279),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_239),
.B(n_0),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_216),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_279),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_213),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_216),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_301),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_224),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_234),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_234),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_227),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_241),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_228),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_302),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_241),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_270),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_239),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_238),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_244),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_245),
.Y(n_452)
);

BUFx6f_ASAP7_75t_SL g453 ( 
.A(n_366),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_257),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_310),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_245),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_361),
.B(n_1),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_267),
.Y(n_458)
);

BUFx6f_ASAP7_75t_SL g459 ( 
.A(n_366),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_312),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_247),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_269),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_247),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_259),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_259),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_361),
.Y(n_466)
);

INVxp33_ASAP7_75t_L g467 ( 
.A(n_206),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_339),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_203),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_275),
.Y(n_470)
);

BUFx10_ASAP7_75t_L g471 ( 
.A(n_270),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_204),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_205),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_233),
.B(n_2),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_275),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_276),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_215),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_218),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_395),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_280),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_281),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_283),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_271),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_284),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_271),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_271),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_271),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_233),
.B(n_2),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_271),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_221),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_222),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_287),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_276),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_230),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_206),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_297),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_309),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_243),
.B(n_5),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_210),
.B(n_5),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_422),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_400),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_422),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_423),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_425),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_430),
.B(n_395),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_479),
.B(n_344),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_401),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_425),
.B(n_243),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_466),
.B(n_434),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_405),
.Y(n_513)
);

INVx6_ASAP7_75t_L g514 ( 
.A(n_471),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_474),
.B(n_344),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_407),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_427),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_428),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_409),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_435),
.B(n_344),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_403),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_438),
.B(n_344),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_471),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_429),
.B(n_226),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_471),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_403),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_433),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_457),
.B(n_277),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_431),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_412),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_431),
.B(n_226),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_488),
.B(n_344),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_448),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_412),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_441),
.B(n_442),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_448),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_483),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_404),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_483),
.B(n_289),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_498),
.B(n_232),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_414),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_485),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_485),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_411),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_414),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_486),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_486),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_487),
.B(n_235),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_487),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_489),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_489),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_444),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_447),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_452),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_456),
.B(n_309),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_461),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_463),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_464),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_465),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_470),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_475),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_476),
.B(n_313),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_493),
.Y(n_566)
);

INVx6_ASAP7_75t_L g567 ( 
.A(n_399),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_497),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_499),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_499),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_416),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_433),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_469),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_436),
.Y(n_574)
);

BUFx8_ASAP7_75t_L g575 ( 
.A(n_453),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_421),
.Y(n_576)
);

OA21x2_ASAP7_75t_L g577 ( 
.A1(n_495),
.A2(n_331),
.B(n_315),
.Y(n_577)
);

BUFx8_ASAP7_75t_L g578 ( 
.A(n_453),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_404),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_555),
.Y(n_580)
);

NOR2x1p5_ASAP7_75t_L g581 ( 
.A(n_572),
.B(n_449),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_569),
.B(n_419),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_507),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_531),
.A2(n_254),
.B1(n_263),
.B2(n_248),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_508),
.B(n_413),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_572),
.B(n_445),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_537),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_508),
.B(n_415),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_502),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_502),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_537),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_555),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_555),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_537),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_514),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_531),
.A2(n_398),
.B1(n_408),
.B2(n_397),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_530),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_L g598 ( 
.A1(n_572),
.A2(n_376),
.B1(n_381),
.B2(n_340),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_530),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_569),
.A2(n_331),
.B1(n_315),
.B2(n_214),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_557),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_502),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_569),
.A2(n_214),
.B1(n_225),
.B2(n_210),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_507),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_572),
.B(n_574),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_502),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_557),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_507),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_512),
.A2(n_317),
.B1(n_304),
.B2(n_305),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_557),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g611 ( 
.A(n_529),
.B(n_472),
.Y(n_611)
);

NOR2x1p5_ASAP7_75t_L g612 ( 
.A(n_572),
.B(n_225),
.Y(n_612)
);

BUFx4f_ASAP7_75t_L g613 ( 
.A(n_577),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_566),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_566),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_573),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_566),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_508),
.B(n_415),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_568),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_572),
.B(n_473),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_514),
.Y(n_621)
);

AND3x2_ASAP7_75t_L g622 ( 
.A(n_522),
.B(n_290),
.C(n_289),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_509),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_568),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_509),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_543),
.B(n_525),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_572),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_572),
.B(n_477),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_537),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_572),
.B(n_478),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_543),
.B(n_418),
.Y(n_631)
);

INVx4_ASAP7_75t_SL g632 ( 
.A(n_514),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_512),
.A2(n_314),
.B1(n_316),
.B2(n_299),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_574),
.B(n_571),
.C(n_443),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_573),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_568),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_533),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_574),
.B(n_490),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_569),
.A2(n_229),
.B1(n_246),
.B2(n_237),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_537),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_509),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_525),
.B(n_418),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_533),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_570),
.A2(n_321),
.B1(n_323),
.B2(n_319),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_509),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_570),
.A2(n_329),
.B1(n_342),
.B2(n_328),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_511),
.Y(n_648)
);

OAI22xp33_ASAP7_75t_L g649 ( 
.A1(n_574),
.A2(n_467),
.B1(n_347),
.B2(n_350),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_570),
.A2(n_348),
.B1(n_355),
.B2(n_354),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_533),
.Y(n_651)
);

CKINVDCx11_ASAP7_75t_R g652 ( 
.A(n_529),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_574),
.B(n_491),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_L g654 ( 
.A(n_574),
.B(n_420),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_567),
.B(n_313),
.Y(n_655)
);

CKINVDCx16_ASAP7_75t_R g656 ( 
.A(n_522),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_507),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_574),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_574),
.B(n_417),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_574),
.B(n_494),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_577),
.B(n_335),
.C(n_333),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_577),
.B(n_335),
.C(n_333),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_522),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_515),
.A2(n_334),
.B1(n_255),
.B2(n_268),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_525),
.B(n_420),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_533),
.Y(n_666)
);

INVx6_ASAP7_75t_L g667 ( 
.A(n_514),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_541),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_L g669 ( 
.A(n_577),
.B(n_353),
.C(n_341),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_533),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_537),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_567),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_511),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_525),
.B(n_432),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_533),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_525),
.B(n_432),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_575),
.B(n_437),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_567),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_544),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_576),
.B(n_450),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_537),
.Y(n_681)
);

AND2x2_ASAP7_75t_SL g682 ( 
.A(n_577),
.B(n_290),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_576),
.B(n_436),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_544),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_511),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_525),
.B(n_437),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_528),
.B(n_440),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_544),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_511),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_544),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_528),
.B(n_440),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_544),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_515),
.A2(n_288),
.B1(n_229),
.B2(n_237),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_544),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_571),
.A2(n_363),
.B1(n_364),
.B2(n_360),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_537),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_507),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_576),
.B(n_451),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_513),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_513),
.Y(n_700)
);

AO21x1_ASAP7_75t_L g701 ( 
.A1(n_535),
.A2(n_353),
.B(n_341),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_513),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_513),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_528),
.B(n_451),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_548),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_548),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_517),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_548),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_535),
.A2(n_285),
.B1(n_246),
.B2(n_255),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_567),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_548),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_517),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_517),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_517),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_541),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_548),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_575),
.B(n_454),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_575),
.B(n_454),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_559),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_548),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_501),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_528),
.B(n_458),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_520),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_520),
.Y(n_724)
);

BUFx8_ASAP7_75t_SL g725 ( 
.A(n_541),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_567),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_501),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_577),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_575),
.B(n_406),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_507),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_577),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_520),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_698),
.B(n_462),
.C(n_458),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_583),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_583),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_589),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_631),
.B(n_579),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_626),
.B(n_528),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_613),
.B(n_528),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_589),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_590),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_683),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_588),
.B(n_618),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_597),
.B(n_579),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_616),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_701),
.A2(n_565),
.B1(n_558),
.B2(n_268),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_604),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_585),
.B(n_579),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_590),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_613),
.B(n_220),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_683),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_604),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_659),
.B(n_567),
.Y(n_753)
);

INVx4_ASAP7_75t_SL g754 ( 
.A(n_667),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_608),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_602),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_659),
.B(n_567),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_698),
.B(n_575),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_608),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_L g760 ( 
.A(n_634),
.B(n_462),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_SL g761 ( 
.A(n_595),
.B(n_514),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_586),
.B(n_551),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_597),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_680),
.B(n_480),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_627),
.B(n_551),
.Y(n_765)
);

BUFx5_ASAP7_75t_L g766 ( 
.A(n_731),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_581),
.B(n_576),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_602),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_L g769 ( 
.A(n_581),
.B(n_236),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_606),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_606),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_582),
.B(n_520),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_654),
.A2(n_424),
.B1(n_426),
.B2(n_410),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_680),
.B(n_480),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_582),
.B(n_547),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_623),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_657),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_682),
.B(n_547),
.Y(n_778)
);

AOI22x1_ASAP7_75t_L g779 ( 
.A1(n_612),
.A2(n_565),
.B1(n_558),
.B2(n_482),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_642),
.B(n_481),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_657),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_674),
.B(n_575),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_682),
.B(n_547),
.Y(n_783)
);

AND2x6_ASAP7_75t_SL g784 ( 
.A(n_620),
.B(n_285),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_706),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_599),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_584),
.B(n_482),
.C(n_481),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_682),
.B(n_547),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_665),
.B(n_484),
.Y(n_789)
);

INVx5_ASAP7_75t_L g790 ( 
.A(n_667),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_676),
.B(n_578),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_686),
.B(n_484),
.Y(n_792)
);

INVx8_ASAP7_75t_L g793 ( 
.A(n_710),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_687),
.B(n_492),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_L g795 ( 
.A(n_728),
.B(n_240),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_613),
.B(n_731),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_697),
.B(n_538),
.Y(n_797)
);

INVx8_ASAP7_75t_L g798 ( 
.A(n_655),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_697),
.B(n_368),
.Y(n_799)
);

OR2x2_ASAP7_75t_SL g800 ( 
.A(n_656),
.B(n_571),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_730),
.Y(n_801)
);

NOR2x1p5_ASAP7_75t_L g802 ( 
.A(n_663),
.B(n_492),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_730),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_656),
.B(n_496),
.C(n_538),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_SL g805 ( 
.A(n_611),
.B(n_578),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_623),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_SL g807 ( 
.A(n_595),
.B(n_514),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_691),
.B(n_510),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_704),
.B(n_510),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_625),
.Y(n_810)
);

NAND2x1_ASAP7_75t_L g811 ( 
.A(n_595),
.B(n_621),
.Y(n_811)
);

AOI22x1_ASAP7_75t_L g812 ( 
.A1(n_612),
.A2(n_558),
.B1(n_565),
.B2(n_496),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_580),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_715),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_722),
.B(n_510),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_706),
.B(n_510),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_706),
.B(n_708),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_715),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_598),
.B(n_578),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_622),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_708),
.B(n_510),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_708),
.Y(n_822)
);

NAND2xp33_ASAP7_75t_L g823 ( 
.A(n_728),
.B(n_249),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_625),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_633),
.B(n_609),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_580),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_633),
.B(n_242),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_716),
.B(n_220),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_592),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_592),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_716),
.B(n_510),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_609),
.B(n_308),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_716),
.B(n_521),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_645),
.B(n_322),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_663),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_645),
.B(n_538),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_593),
.B(n_521),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_593),
.B(n_521),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_628),
.B(n_578),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_601),
.B(n_523),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_655),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_630),
.A2(n_439),
.B1(n_446),
.B2(n_455),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_601),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_607),
.B(n_610),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_647),
.B(n_367),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_607),
.B(n_523),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_701),
.A2(n_286),
.B1(n_288),
.B2(n_291),
.Y(n_847)
);

O2A1O1Ixp5_ASAP7_75t_L g848 ( 
.A1(n_661),
.A2(n_542),
.B(n_526),
.C(n_534),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_610),
.B(n_523),
.Y(n_849)
);

NAND2x1_ASAP7_75t_L g850 ( 
.A(n_621),
.B(n_514),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_614),
.B(n_559),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_641),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_614),
.B(n_615),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_668),
.B(n_377),
.C(n_375),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_615),
.B(n_559),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_617),
.B(n_559),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_647),
.B(n_380),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_617),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_638),
.A2(n_460),
.B1(n_468),
.B2(n_324),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_619),
.B(n_559),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_653),
.B(n_578),
.Y(n_861)
);

AND2x2_ASAP7_75t_SL g862 ( 
.A(n_660),
.B(n_605),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_619),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_624),
.B(n_559),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_624),
.B(n_559),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_641),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_655),
.A2(n_383),
.B1(n_306),
.B2(n_318),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_672),
.B(n_220),
.Y(n_868)
);

NAND2x1_ASAP7_75t_L g869 ( 
.A(n_621),
.B(n_501),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_636),
.B(n_559),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_655),
.A2(n_369),
.B1(n_368),
.B2(n_373),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_SL g872 ( 
.A(n_729),
.B(n_578),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_636),
.B(n_559),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_637),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_658),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_672),
.B(n_220),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_596),
.B(n_382),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_658),
.B(n_373),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_637),
.B(n_562),
.Y(n_879)
);

NOR3xp33_ASAP7_75t_L g880 ( 
.A(n_668),
.B(n_390),
.C(n_388),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_655),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_650),
.B(n_391),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_661),
.A2(n_291),
.B1(n_286),
.B2(n_296),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_643),
.B(n_562),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_643),
.B(n_562),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_672),
.B(n_220),
.Y(n_886)
);

INVx8_ASAP7_75t_L g887 ( 
.A(n_725),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_651),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_651),
.B(n_562),
.Y(n_889)
);

INVx8_ASAP7_75t_L g890 ( 
.A(n_616),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_695),
.B(n_650),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_649),
.B(n_250),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_666),
.B(n_670),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_662),
.B(n_669),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_L g895 ( 
.A(n_695),
.B(n_393),
.C(n_392),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_666),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_670),
.B(n_562),
.Y(n_897)
);

O2A1O1Ixp5_ASAP7_75t_L g898 ( 
.A1(n_662),
.A2(n_542),
.B(n_526),
.C(n_534),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_675),
.B(n_394),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_675),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_672),
.B(n_678),
.Y(n_901)
);

NOR2xp67_ASAP7_75t_L g902 ( 
.A(n_669),
.B(n_556),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_679),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_L g904 ( 
.A(n_679),
.B(n_251),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_684),
.B(n_562),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_744),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_743),
.B(n_684),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_743),
.A2(n_717),
.B1(n_718),
.B2(n_677),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_811),
.A2(n_850),
.B(n_901),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_901),
.A2(n_591),
.B(n_587),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_L g911 ( 
.A(n_766),
.B(n_798),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_762),
.A2(n_667),
.B1(n_600),
.B2(n_639),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_737),
.B(n_688),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_L g914 ( 
.A(n_733),
.B(n_664),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_843),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_SL g916 ( 
.A(n_745),
.B(n_635),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_737),
.B(n_780),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_734),
.B(n_688),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_825),
.A2(n_827),
.B(n_832),
.C(n_834),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_843),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_780),
.B(n_690),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_789),
.B(n_690),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_789),
.B(n_692),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_734),
.B(n_692),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_825),
.A2(n_705),
.B(n_711),
.C(n_694),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_797),
.B(n_694),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_748),
.B(n_705),
.Y(n_927)
);

AOI33xp33_ASAP7_75t_L g928 ( 
.A1(n_891),
.A2(n_693),
.A3(n_709),
.B1(n_298),
.B2(n_300),
.B3(n_296),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_792),
.B(n_711),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_858),
.Y(n_930)
);

NOR2xp67_ASAP7_75t_SL g931 ( 
.A(n_819),
.B(n_841),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_792),
.B(n_720),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_827),
.A2(n_720),
.B(n_724),
.C(n_603),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_862),
.A2(n_667),
.B1(n_369),
.B2(n_386),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_794),
.B(n_594),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_858),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_766),
.B(n_678),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_794),
.B(n_594),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_863),
.B(n_594),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_778),
.A2(n_724),
.B(n_648),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_863),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_763),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_783),
.A2(n_648),
.B(n_646),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_874),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_788),
.A2(n_775),
.B(n_772),
.Y(n_945)
);

O2A1O1Ixp5_ASAP7_75t_L g946 ( 
.A1(n_738),
.A2(n_696),
.B(n_629),
.C(n_640),
.Y(n_946)
);

AOI21x1_ASAP7_75t_L g947 ( 
.A1(n_750),
.A2(n_673),
.B(n_646),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_765),
.A2(n_591),
.B(n_587),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_862),
.A2(n_386),
.B1(n_253),
.B2(n_727),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_742),
.B(n_629),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_738),
.A2(n_591),
.B(n_587),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_795),
.A2(n_591),
.B(n_587),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_823),
.A2(n_591),
.B(n_587),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_751),
.B(n_629),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_739),
.A2(n_681),
.B(n_644),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_764),
.B(n_652),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_748),
.B(n_640),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_890),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_739),
.A2(n_681),
.B(n_644),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_767),
.B(n_640),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_832),
.A2(n_671),
.B1(n_696),
.B2(n_726),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_750),
.A2(n_681),
.B(n_644),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_796),
.A2(n_681),
.B(n_644),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_813),
.B(n_671),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_888),
.Y(n_965)
);

OAI21xp33_ASAP7_75t_L g966 ( 
.A1(n_834),
.A2(n_349),
.B(n_346),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_796),
.A2(n_681),
.B(n_644),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_892),
.A2(n_732),
.B(n_673),
.C(n_723),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_764),
.B(n_671),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_826),
.B(n_696),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_836),
.A2(n_732),
.B(n_723),
.C(n_714),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_822),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_890),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_894),
.A2(n_719),
.B(n_689),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_868),
.A2(n_719),
.B(n_689),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_848),
.A2(n_699),
.B(n_685),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_829),
.B(n_685),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_SL g978 ( 
.A(n_890),
.B(n_453),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_830),
.Y(n_979)
);

NOR2x1p5_ASAP7_75t_L g980 ( 
.A(n_882),
.B(n_298),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_797),
.B(n_721),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_836),
.B(n_678),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_868),
.A2(n_719),
.B(n_700),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_753),
.B(n_699),
.Y(n_984)
);

AOI21xp33_ASAP7_75t_L g985 ( 
.A1(n_845),
.A2(n_258),
.B(n_252),
.Y(n_985)
);

AOI21x1_ASAP7_75t_L g986 ( 
.A1(n_817),
.A2(n_702),
.B(n_700),
.Y(n_986)
);

NOR3xp33_ASAP7_75t_L g987 ( 
.A(n_845),
.B(n_320),
.C(n_300),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_774),
.B(n_678),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_876),
.A2(n_719),
.B(n_703),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_774),
.B(n_702),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_766),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_896),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_876),
.A2(n_886),
.B(n_869),
.Y(n_993)
);

OAI21xp33_ASAP7_75t_L g994 ( 
.A1(n_857),
.A2(n_332),
.B(n_320),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_SL g995 ( 
.A(n_805),
.B(n_459),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_886),
.A2(n_719),
.B(n_707),
.Y(n_996)
);

OAI21xp33_ASAP7_75t_SL g997 ( 
.A1(n_817),
.A2(n_853),
.B(n_844),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_808),
.A2(n_707),
.B(n_703),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_898),
.A2(n_902),
.B(n_833),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_L g1000 ( 
.A(n_766),
.B(n_356),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_900),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_816),
.A2(n_713),
.B(n_712),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_753),
.B(n_712),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_857),
.A2(n_714),
.B(n_713),
.C(n_556),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_809),
.A2(n_727),
.B1(n_721),
.B2(n_278),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_815),
.A2(n_632),
.B(n_727),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_757),
.B(n_721),
.Y(n_1007)
);

AOI21x1_ASAP7_75t_L g1008 ( 
.A1(n_821),
.A2(n_503),
.B(n_500),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_903),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_831),
.A2(n_632),
.B(n_726),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_736),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_837),
.A2(n_556),
.B(n_561),
.C(n_560),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_752),
.B(n_556),
.Y(n_1013)
);

NOR2x1_ASAP7_75t_L g1014 ( 
.A(n_757),
.B(n_560),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_766),
.B(n_726),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_899),
.B(n_726),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_785),
.A2(n_632),
.B(n_561),
.Y(n_1017)
);

AOI21xp33_ASAP7_75t_L g1018 ( 
.A1(n_877),
.A2(n_262),
.B(n_261),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_899),
.B(n_838),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_740),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_741),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_893),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_840),
.B(n_560),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_847),
.A2(n_332),
.B(n_334),
.C(n_337),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_747),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_SL g1026 ( 
.A1(n_828),
.A2(n_879),
.B(n_885),
.C(n_884),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_846),
.A2(n_632),
.B(n_561),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_849),
.B(n_560),
.Y(n_1028)
);

NOR2x1p5_ASAP7_75t_SL g1029 ( 
.A(n_766),
.B(n_561),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_875),
.A2(n_534),
.B(n_526),
.Y(n_1030)
);

OAI321xp33_ASAP7_75t_L g1031 ( 
.A1(n_895),
.A2(n_847),
.A3(n_746),
.B1(n_814),
.B2(n_883),
.C(n_859),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_878),
.B(n_755),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_763),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_878),
.B(n_562),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_759),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_822),
.B(n_356),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_822),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_818),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_777),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_822),
.B(n_356),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_752),
.B(n_526),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_851),
.A2(n_856),
.B(n_855),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_875),
.A2(n_534),
.B(n_526),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_781),
.B(n_562),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_801),
.B(n_562),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_818),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_SL g1047 ( 
.A(n_872),
.B(n_459),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_860),
.A2(n_534),
.B(n_526),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_864),
.A2(n_542),
.B(n_534),
.Y(n_1049)
);

CKINVDCx10_ASAP7_75t_R g1050 ( 
.A(n_887),
.Y(n_1050)
);

AO21x1_ASAP7_75t_L g1051 ( 
.A1(n_782),
.A2(n_542),
.B(n_385),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_803),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_749),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_756),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_746),
.B(n_563),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_793),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_769),
.A2(n_542),
.B(n_563),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_786),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_865),
.A2(n_542),
.B(n_536),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_768),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_761),
.A2(n_564),
.B(n_563),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_760),
.B(n_563),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_835),
.Y(n_1063)
);

O2A1O1Ixp5_ASAP7_75t_L g1064 ( 
.A1(n_839),
.A2(n_505),
.B(n_503),
.C(n_504),
.Y(n_1064)
);

O2A1O1Ixp5_ASAP7_75t_L g1065 ( 
.A1(n_861),
.A2(n_505),
.B(n_503),
.C(n_504),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_770),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_758),
.A2(n_396),
.B(n_371),
.C(n_362),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_841),
.B(n_500),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_807),
.A2(n_564),
.B(n_563),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_842),
.B(n_337),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_752),
.B(n_563),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_771),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_787),
.B(n_351),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_752),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_883),
.A2(n_362),
.B1(n_371),
.B2(n_396),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_790),
.A2(n_564),
.B(n_563),
.Y(n_1076)
);

NOR2x2_ASAP7_75t_L g1077 ( 
.A(n_784),
.B(n_459),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_773),
.B(n_351),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_870),
.A2(n_524),
.B(n_500),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_800),
.B(n_264),
.Y(n_1080)
);

OR2x6_ASAP7_75t_L g1081 ( 
.A(n_798),
.B(n_356),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_793),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_735),
.B(n_563),
.Y(n_1083)
);

INVxp67_ASAP7_75t_SL g1084 ( 
.A(n_881),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_790),
.A2(n_873),
.B(n_889),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_735),
.A2(n_378),
.B1(n_266),
.B2(n_272),
.Y(n_1086)
);

BUFx12f_ASAP7_75t_L g1087 ( 
.A(n_820),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_779),
.B(n_563),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_776),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_881),
.B(n_504),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_L g1091 ( 
.A(n_804),
.B(n_358),
.C(n_357),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_897),
.A2(n_905),
.B(n_799),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_812),
.B(n_799),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_802),
.B(n_357),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_806),
.B(n_564),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_810),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_854),
.B(n_265),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_880),
.B(n_505),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_824),
.B(n_852),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_979),
.Y(n_1100)
);

AOI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_919),
.A2(n_385),
.B1(n_389),
.B2(n_358),
.C(n_379),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_917),
.A2(n_908),
.B(n_914),
.C(n_1031),
.Y(n_1102)
);

INVx4_ASAP7_75t_L g1103 ( 
.A(n_958),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_926),
.B(n_754),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1070),
.B(n_793),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1078),
.B(n_867),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_981),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1022),
.B(n_798),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_906),
.B(n_791),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_992),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_981),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1019),
.B(n_866),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_SL g1113 ( 
.A1(n_925),
.A2(n_871),
.B(n_379),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_982),
.A2(n_904),
.B1(n_273),
.B2(n_330),
.Y(n_1114)
);

BUFx12f_ASAP7_75t_L g1115 ( 
.A(n_1087),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_979),
.Y(n_1116)
);

BUFx12f_ASAP7_75t_L g1117 ( 
.A(n_1087),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_956),
.B(n_389),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_913),
.B(n_828),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_981),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_991),
.A2(n_790),
.B(n_754),
.Y(n_1121)
);

NAND2xp33_ASAP7_75t_L g1122 ( 
.A(n_982),
.B(n_790),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1013),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1050),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_913),
.B(n_754),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_927),
.B(n_990),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_927),
.B(n_506),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1073),
.B(n_887),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_990),
.B(n_506),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_991),
.A2(n_356),
.B(n_359),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1001),
.Y(n_1131)
);

BUFx12f_ASAP7_75t_L g1132 ( 
.A(n_1056),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1056),
.Y(n_1133)
);

OAI22x1_ASAP7_75t_L g1134 ( 
.A1(n_980),
.A2(n_887),
.B1(n_384),
.B2(n_374),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_988),
.B(n_506),
.Y(n_1135)
);

BUFx8_ASAP7_75t_L g1136 ( 
.A(n_958),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1038),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_985),
.A2(n_539),
.B(n_516),
.C(n_518),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_918),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_991),
.A2(n_387),
.B(n_359),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_907),
.B(n_516),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_920),
.B(n_274),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_942),
.B(n_292),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_957),
.B(n_516),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1000),
.A2(n_359),
.B(n_387),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1033),
.B(n_293),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1046),
.B(n_294),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_920),
.B(n_936),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1000),
.A2(n_359),
.B(n_387),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_957),
.B(n_969),
.Y(n_1150)
);

INVx4_ASAP7_75t_L g1151 ( 
.A(n_973),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1001),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_1084),
.A2(n_303),
.B1(n_295),
.B2(n_325),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_987),
.A2(n_540),
.B(n_518),
.C(n_519),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_969),
.B(n_518),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_945),
.A2(n_524),
.B(n_519),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_973),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_SL g1158 ( 
.A1(n_931),
.A2(n_524),
.B(n_519),
.C(n_527),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1058),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1009),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1016),
.A2(n_359),
.B(n_387),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1009),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_937),
.A2(n_387),
.B(n_564),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1063),
.B(n_326),
.Y(n_1164)
);

CKINVDCx16_ASAP7_75t_R g1165 ( 
.A(n_916),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_944),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_936),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1094),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_965),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_997),
.A2(n_336),
.B(n_338),
.C(n_343),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1068),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_1097),
.B(n_345),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1068),
.B(n_527),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_SL g1174 ( 
.A1(n_995),
.A2(n_352),
.B1(n_365),
.B2(n_370),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1090),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1090),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_915),
.B(n_372),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1075),
.A2(n_545),
.B1(n_527),
.B2(n_532),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_930),
.B(n_7),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_1082),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_L g1181 ( 
.A1(n_1093),
.A2(n_546),
.B(n_536),
.C(n_539),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_941),
.B(n_564),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_926),
.B(n_564),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_926),
.B(n_564),
.Y(n_1184)
);

NAND2x2_ASAP7_75t_L g1185 ( 
.A(n_1077),
.B(n_8),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1011),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_918),
.Y(n_1187)
);

OAI21xp33_ASAP7_75t_SL g1188 ( 
.A1(n_999),
.A2(n_546),
.B(n_532),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_937),
.A2(n_564),
.B(n_554),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_1098),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_921),
.A2(n_923),
.B1(n_929),
.B2(n_922),
.Y(n_1191)
);

AOI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_1018),
.A2(n_9),
.B(n_10),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_SL g1193 ( 
.A(n_978),
.B(n_532),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_932),
.B(n_536),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1011),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1020),
.Y(n_1196)
);

BUFx4f_ASAP7_75t_SL g1197 ( 
.A(n_1098),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1025),
.B(n_10),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1035),
.B(n_11),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_994),
.A2(n_546),
.B(n_539),
.C(n_552),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_933),
.A2(n_549),
.B(n_540),
.C(n_552),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1039),
.B(n_540),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1052),
.B(n_545),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_918),
.B(n_78),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_SL g1205 ( 
.A(n_1047),
.B(n_545),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1032),
.B(n_966),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1021),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_R g1208 ( 
.A(n_911),
.B(n_193),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_924),
.B(n_552),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1015),
.A2(n_554),
.B(n_553),
.Y(n_1210)
);

NAND2x2_ASAP7_75t_L g1211 ( 
.A(n_1077),
.B(n_12),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_928),
.B(n_549),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1021),
.Y(n_1213)
);

NAND2x1p5_ASAP7_75t_L g1214 ( 
.A(n_972),
.B(n_501),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_928),
.B(n_549),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1097),
.B(n_16),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_924),
.B(n_1080),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1080),
.B(n_17),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_949),
.A2(n_553),
.B(n_550),
.C(n_554),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_924),
.B(n_19),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1007),
.B(n_554),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1013),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_935),
.A2(n_553),
.B1(n_550),
.B2(n_501),
.Y(n_1223)
);

BUFx12f_ASAP7_75t_L g1224 ( 
.A(n_1081),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1054),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1013),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_984),
.B(n_1003),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1015),
.A2(n_553),
.B(n_550),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_974),
.A2(n_550),
.B(n_501),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1074),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1054),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1091),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1075),
.B(n_24),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1086),
.B(n_80),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_938),
.B(n_27),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_950),
.B(n_27),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_972),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1055),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_954),
.B(n_36),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_909),
.A2(n_89),
.B(n_187),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1060),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_911),
.A2(n_84),
.B(n_178),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1053),
.B(n_36),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_972),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1024),
.A2(n_37),
.B(n_40),
.C(n_42),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1023),
.B(n_44),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1037),
.B(n_97),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1060),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_952),
.A2(n_93),
.B(n_169),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1089),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1066),
.B(n_45),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_953),
.A2(n_91),
.B(n_159),
.Y(n_1252)
);

AOI21xp33_ASAP7_75t_L g1253 ( 
.A1(n_912),
.A2(n_45),
.B(n_46),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1028),
.B(n_49),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1072),
.B(n_49),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1089),
.B(n_52),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_960),
.B(n_53),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1096),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_948),
.A2(n_108),
.B(n_152),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_L g1260 ( 
.A(n_1024),
.B(n_55),
.C(n_60),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1067),
.B(n_1037),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1096),
.B(n_61),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1042),
.B(n_61),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1189),
.A2(n_1092),
.B(n_947),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1190),
.B(n_1168),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1126),
.B(n_1014),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1102),
.A2(n_998),
.B(n_1004),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1171),
.B(n_977),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1122),
.A2(n_1010),
.B(n_1026),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1150),
.A2(n_971),
.B(n_946),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1216),
.A2(n_934),
.B1(n_1051),
.B2(n_1081),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_1137),
.Y(n_1272)
);

OAI22x1_ASAP7_75t_L g1273 ( 
.A1(n_1216),
.A2(n_1190),
.B1(n_1218),
.B2(n_1106),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1227),
.A2(n_1026),
.B(n_993),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1191),
.A2(n_1059),
.B(n_940),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1192),
.A2(n_1064),
.B(n_1065),
.C(n_1040),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1263),
.A2(n_1005),
.B(n_1043),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1206),
.A2(n_1197),
.B1(n_1220),
.B2(n_1217),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1188),
.A2(n_1170),
.B(n_1181),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1105),
.B(n_1037),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1110),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1135),
.A2(n_1006),
.B(n_955),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1112),
.A2(n_959),
.B(n_951),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1165),
.B(n_1099),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1119),
.A2(n_1057),
.B(n_910),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1221),
.A2(n_1049),
.B(n_1048),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1161),
.A2(n_1088),
.A3(n_1062),
.B(n_962),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1206),
.A2(n_1081),
.B1(n_1034),
.B2(n_939),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1175),
.B(n_964),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1155),
.A2(n_1125),
.B(n_1144),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1129),
.A2(n_1083),
.B(n_1085),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1127),
.A2(n_1081),
.B(n_976),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_SL g1293 ( 
.A1(n_1234),
.A2(n_1040),
.B(n_1036),
.C(n_970),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1137),
.B(n_1041),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1166),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1253),
.A2(n_1029),
.B(n_1012),
.C(n_1092),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1201),
.A2(n_1061),
.A3(n_1069),
.B(n_963),
.Y(n_1297)
);

NOR2xp67_ASAP7_75t_L g1298 ( 
.A(n_1108),
.B(n_1071),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1172),
.A2(n_961),
.B(n_968),
.C(n_1030),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1176),
.B(n_943),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1167),
.B(n_1041),
.Y(n_1301)
);

AOI211x1_ASAP7_75t_L g1302 ( 
.A1(n_1233),
.A2(n_1036),
.B(n_1008),
.C(n_1079),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1210),
.A2(n_986),
.B(n_1228),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1139),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1167),
.B(n_1002),
.Y(n_1305)
);

INVx5_ASAP7_75t_L g1306 ( 
.A(n_1139),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1235),
.A2(n_1044),
.B(n_1045),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1159),
.B(n_967),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1160),
.Y(n_1309)
);

OAI22x1_ASAP7_75t_L g1310 ( 
.A1(n_1109),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_1310)
);

INVxp67_ASAP7_75t_SL g1311 ( 
.A(n_1187),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1163),
.A2(n_1027),
.A3(n_975),
.B(n_996),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1257),
.A2(n_989),
.B(n_983),
.Y(n_1313)
);

NOR2xp67_ASAP7_75t_L g1314 ( 
.A(n_1123),
.B(n_1017),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1187),
.B(n_1095),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1159),
.B(n_1076),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1246),
.A2(n_1254),
.B(n_1261),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1236),
.A2(n_1239),
.B(n_1101),
.C(n_1232),
.Y(n_1318)
);

AO21x2_ASAP7_75t_L g1319 ( 
.A1(n_1158),
.A2(n_112),
.B(n_139),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1141),
.A2(n_110),
.B(n_137),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1194),
.A2(n_107),
.B(n_126),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1118),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1169),
.B(n_67),
.Y(n_1323)
);

CKINVDCx16_ASAP7_75t_R g1324 ( 
.A(n_1132),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1229),
.A2(n_115),
.B(n_119),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1222),
.B(n_69),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1107),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1156),
.A2(n_101),
.B(n_118),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_SL g1329 ( 
.A1(n_1158),
.A2(n_117),
.B(n_189),
.C(n_75),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1147),
.B(n_1146),
.Y(n_1330)
);

O2A1O1Ixp5_ASAP7_75t_L g1331 ( 
.A1(n_1236),
.A2(n_69),
.B(n_74),
.C(n_76),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1222),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_SL g1333 ( 
.A(n_1205),
.B(n_1193),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1128),
.B(n_1164),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1104),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1197),
.B(n_1107),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_R g1337 ( 
.A(n_1180),
.B(n_1124),
.Y(n_1337)
);

AND2x6_ASAP7_75t_L g1338 ( 
.A(n_1204),
.B(n_1104),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1226),
.B(n_1239),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1130),
.A2(n_1140),
.A3(n_1223),
.B(n_1256),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1143),
.B(n_1220),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1181),
.A2(n_1121),
.B(n_1259),
.Y(n_1342)
);

OAI22x1_ASAP7_75t_L g1343 ( 
.A1(n_1198),
.A2(n_1199),
.B1(n_1179),
.B2(n_1260),
.Y(n_1343)
);

NAND4xp25_ASAP7_75t_SL g1344 ( 
.A(n_1238),
.B(n_1245),
.C(n_1174),
.D(n_1242),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1136),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1198),
.A2(n_1199),
.B1(n_1238),
.B2(n_1179),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1107),
.B(n_1111),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1100),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1116),
.Y(n_1349)
);

NAND2xp33_ASAP7_75t_SL g1350 ( 
.A(n_1208),
.B(n_1103),
.Y(n_1350)
);

AOI221x1_ASAP7_75t_L g1351 ( 
.A1(n_1113),
.A2(n_1153),
.B1(n_1149),
.B2(n_1145),
.C(n_1252),
.Y(n_1351)
);

INVx3_ASAP7_75t_SL g1352 ( 
.A(n_1133),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1139),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1131),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1143),
.B(n_1107),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1356)
);

AOI221xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1212),
.A2(n_1215),
.B1(n_1256),
.B2(n_1262),
.C(n_1173),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1138),
.A2(n_1219),
.B(n_1240),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1136),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1262),
.A2(n_1249),
.A3(n_1251),
.B(n_1162),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1182),
.A2(n_1214),
.B(n_1148),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1183),
.A2(n_1184),
.B(n_1142),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1202),
.A2(n_1203),
.B(n_1207),
.Y(n_1363)
);

INVx6_ASAP7_75t_L g1364 ( 
.A(n_1115),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1251),
.A2(n_1114),
.B(n_1204),
.C(n_1152),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1226),
.A2(n_1139),
.B1(n_1123),
.B2(n_1230),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1186),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1177),
.A2(n_1209),
.B(n_1247),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1111),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1120),
.A2(n_1174),
.B1(n_1250),
.B2(n_1241),
.Y(n_1371)
);

AO221x1_ASAP7_75t_L g1372 ( 
.A1(n_1134),
.A2(n_1244),
.B1(n_1237),
.B2(n_1258),
.C(n_1196),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1120),
.B(n_1213),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1225),
.B(n_1248),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1243),
.A2(n_1255),
.B1(n_1224),
.B2(n_1195),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1154),
.A2(n_1200),
.B(n_1231),
.C(n_1247),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1103),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1185),
.A2(n_1211),
.B1(n_1178),
.B2(n_1157),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1214),
.A2(n_1178),
.B(n_1151),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1208),
.A2(n_1151),
.A3(n_1157),
.B(n_1237),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1237),
.A2(n_1244),
.B(n_1185),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1237),
.A2(n_1244),
.B(n_1211),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1244),
.Y(n_1383)
);

CKINVDCx9p33_ASAP7_75t_R g1384 ( 
.A(n_1117),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1126),
.A2(n_917),
.B1(n_919),
.B2(n_908),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1136),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1165),
.B(n_919),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1166),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1126),
.B(n_917),
.Y(n_1389)
);

CKINVDCx6p67_ASAP7_75t_R g1390 ( 
.A(n_1115),
.Y(n_1390)
);

OR2x2_ASAP7_75t_SL g1391 ( 
.A(n_1165),
.B(n_656),
.Y(n_1391)
);

INVx4_ASAP7_75t_L g1392 ( 
.A(n_1103),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1190),
.B(n_919),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1126),
.A2(n_917),
.B1(n_919),
.B2(n_908),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1102),
.A2(n_1170),
.A3(n_1191),
.B(n_1051),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1102),
.A2(n_919),
.B(n_917),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1104),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1189),
.A2(n_1092),
.B(n_947),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1122),
.A2(n_991),
.B(n_811),
.Y(n_1399)
);

OAI22x1_ASAP7_75t_L g1400 ( 
.A1(n_1216),
.A2(n_825),
.B1(n_908),
.B2(n_1190),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1216),
.A2(n_825),
.B1(n_611),
.B2(n_832),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1133),
.Y(n_1402)
);

AO31x2_ASAP7_75t_L g1403 ( 
.A1(n_1102),
.A2(n_1170),
.A3(n_1191),
.B(n_1051),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1126),
.B(n_917),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1110),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1126),
.B(n_917),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1126),
.B(n_917),
.Y(n_1407)
);

CKINVDCx11_ASAP7_75t_R g1408 ( 
.A(n_1115),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1122),
.A2(n_991),
.B(n_811),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1122),
.A2(n_991),
.B(n_811),
.Y(n_1410)
);

BUFx12f_ASAP7_75t_L g1411 ( 
.A(n_1115),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1102),
.A2(n_919),
.B(n_1150),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1216),
.A2(n_919),
.B(n_917),
.C(n_825),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1105),
.B(n_1106),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1122),
.A2(n_991),
.B(n_811),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1104),
.B(n_1120),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1102),
.A2(n_919),
.B(n_1150),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1126),
.B(n_917),
.Y(n_1418)
);

AO31x2_ASAP7_75t_L g1419 ( 
.A1(n_1102),
.A2(n_1170),
.A3(n_1191),
.B(n_1051),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1104),
.B(n_1120),
.Y(n_1420)
);

OR2x6_ASAP7_75t_L g1421 ( 
.A(n_1132),
.B(n_798),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1190),
.B(n_919),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1122),
.A2(n_991),
.B(n_811),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1166),
.Y(n_1424)
);

AO31x2_ASAP7_75t_L g1425 ( 
.A1(n_1102),
.A2(n_1170),
.A3(n_1191),
.B(n_1051),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1126),
.B(n_917),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1126),
.A2(n_917),
.B1(n_919),
.B2(n_908),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1190),
.B(n_919),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1110),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1126),
.B(n_917),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1122),
.A2(n_991),
.B(n_811),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1126),
.B(n_917),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1136),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1352),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1388),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1401),
.A2(n_1346),
.B1(n_1343),
.B2(n_1396),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1346),
.A2(n_1394),
.B1(n_1385),
.B2(n_1427),
.Y(n_1437)
);

BUFx8_ASAP7_75t_SL g1438 ( 
.A(n_1411),
.Y(n_1438)
);

INVx6_ASAP7_75t_L g1439 ( 
.A(n_1304),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1344),
.A2(n_1387),
.B1(n_1400),
.B2(n_1428),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1408),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1424),
.Y(n_1442)
);

BUFx8_ASAP7_75t_L g1443 ( 
.A(n_1334),
.Y(n_1443)
);

BUFx12f_ASAP7_75t_L g1444 ( 
.A(n_1364),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1281),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1412),
.A2(n_1417),
.B1(n_1393),
.B2(n_1422),
.Y(n_1446)
);

INVx6_ASAP7_75t_L g1447 ( 
.A(n_1304),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1412),
.A2(n_1417),
.B1(n_1310),
.B2(n_1341),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1390),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1348),
.Y(n_1450)
);

BUFx8_ASAP7_75t_L g1451 ( 
.A(n_1345),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1402),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1327),
.Y(n_1453)
);

BUFx12f_ASAP7_75t_L g1454 ( 
.A(n_1364),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1349),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1389),
.B(n_1404),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1354),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1333),
.A2(n_1414),
.B1(n_1275),
.B2(n_1407),
.Y(n_1458)
);

INVx6_ASAP7_75t_L g1459 ( 
.A(n_1306),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1273),
.A2(n_1333),
.B1(n_1372),
.B2(n_1278),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1367),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1278),
.A2(n_1284),
.B1(n_1330),
.B2(n_1406),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1418),
.A2(n_1426),
.B1(n_1430),
.B2(n_1432),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1413),
.A2(n_1318),
.B1(n_1375),
.B2(n_1365),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1309),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1322),
.B(n_1339),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1371),
.A2(n_1355),
.B1(n_1338),
.B2(n_1328),
.Y(n_1467)
);

INVx5_ASAP7_75t_SL g1468 ( 
.A(n_1384),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1265),
.A2(n_1375),
.B1(n_1368),
.B2(n_1338),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1338),
.A2(n_1271),
.B1(n_1326),
.B2(n_1317),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1405),
.Y(n_1471)
);

CKINVDCx11_ASAP7_75t_R g1472 ( 
.A(n_1324),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1429),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1337),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1359),
.Y(n_1475)
);

AOI21xp33_ASAP7_75t_L g1476 ( 
.A1(n_1357),
.A2(n_1277),
.B(n_1271),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1338),
.A2(n_1323),
.B1(n_1279),
.B2(n_1379),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1378),
.A2(n_1336),
.B1(n_1280),
.B2(n_1350),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1374),
.Y(n_1479)
);

BUFx12f_ASAP7_75t_L g1480 ( 
.A(n_1391),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1373),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1386),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1266),
.A2(n_1268),
.B1(n_1358),
.B2(n_1279),
.Y(n_1483)
);

BUFx12f_ASAP7_75t_L g1484 ( 
.A(n_1421),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1332),
.B(n_1272),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1358),
.A2(n_1267),
.B1(n_1286),
.B2(n_1289),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1316),
.A2(n_1308),
.B1(n_1378),
.B2(n_1362),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1294),
.B(n_1311),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1433),
.A2(n_1421),
.B1(n_1377),
.B2(n_1392),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1369),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1267),
.A2(n_1292),
.B1(n_1300),
.B2(n_1290),
.Y(n_1491)
);

NAND2x1p5_ASAP7_75t_L g1492 ( 
.A(n_1306),
.B(n_1377),
.Y(n_1492)
);

BUFx8_ASAP7_75t_L g1493 ( 
.A(n_1416),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1370),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1298),
.A2(n_1357),
.B1(n_1366),
.B2(n_1420),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1320),
.A2(n_1321),
.B(n_1288),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1363),
.Y(n_1497)
);

INVx6_ASAP7_75t_L g1498 ( 
.A(n_1392),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1416),
.B(n_1420),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1315),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1301),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1298),
.A2(n_1314),
.B1(n_1288),
.B2(n_1356),
.Y(n_1502)
);

BUFx10_ASAP7_75t_L g1503 ( 
.A(n_1421),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1305),
.A2(n_1376),
.B1(n_1397),
.B2(n_1335),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1335),
.B(n_1397),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1383),
.Y(n_1506)
);

INVx6_ASAP7_75t_L g1507 ( 
.A(n_1356),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1382),
.A2(n_1302),
.B1(n_1353),
.B2(n_1347),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1381),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1270),
.A2(n_1351),
.B1(n_1331),
.B2(n_1274),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1360),
.B(n_1380),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1380),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1380),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1361),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1360),
.Y(n_1515)
);

CKINVDCx11_ASAP7_75t_R g1516 ( 
.A(n_1329),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1313),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1283),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1319),
.A2(n_1285),
.B1(n_1325),
.B2(n_1291),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1319),
.A2(n_1282),
.B1(n_1269),
.B2(n_1303),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1342),
.A2(n_1264),
.B1(n_1398),
.B2(n_1431),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1293),
.A2(n_1299),
.B1(n_1296),
.B2(n_1415),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1399),
.A2(n_1423),
.B1(n_1410),
.B2(n_1409),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1307),
.B(n_1425),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1395),
.Y(n_1525)
);

CKINVDCx6p67_ASAP7_75t_R g1526 ( 
.A(n_1276),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1395),
.A2(n_1403),
.B1(n_1419),
.B2(n_1425),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1395),
.Y(n_1528)
);

INVx8_ASAP7_75t_L g1529 ( 
.A(n_1403),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1403),
.Y(n_1530)
);

BUFx4f_ASAP7_75t_SL g1531 ( 
.A(n_1419),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1419),
.Y(n_1532)
);

CKINVDCx8_ASAP7_75t_R g1533 ( 
.A(n_1425),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1297),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1340),
.A2(n_1297),
.B1(n_1287),
.B2(n_1312),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1312),
.Y(n_1536)
);

BUFx8_ASAP7_75t_L g1537 ( 
.A(n_1340),
.Y(n_1537)
);

INVx6_ASAP7_75t_L g1538 ( 
.A(n_1287),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1295),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1333),
.A2(n_825),
.B1(n_1216),
.B2(n_832),
.Y(n_1540)
);

INVx6_ASAP7_75t_L g1541 ( 
.A(n_1304),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_1337),
.Y(n_1542)
);

BUFx4f_ASAP7_75t_SL g1543 ( 
.A(n_1411),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1401),
.A2(n_919),
.B1(n_917),
.B2(n_1346),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1281),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1337),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1337),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1389),
.B(n_1404),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1332),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1332),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_1337),
.Y(n_1551)
);

BUFx12f_ASAP7_75t_L g1552 ( 
.A(n_1408),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1304),
.B(n_1306),
.Y(n_1553)
);

BUFx8_ASAP7_75t_L g1554 ( 
.A(n_1411),
.Y(n_1554)
);

INVx6_ASAP7_75t_L g1555 ( 
.A(n_1304),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1401),
.A2(n_1216),
.B1(n_1346),
.B2(n_825),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1333),
.A2(n_825),
.B1(n_1216),
.B2(n_832),
.Y(n_1557)
);

BUFx12f_ASAP7_75t_L g1558 ( 
.A(n_1408),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1281),
.Y(n_1559)
);

INVx6_ASAP7_75t_L g1560 ( 
.A(n_1304),
.Y(n_1560)
);

OAI22xp33_ASAP7_75t_R g1561 ( 
.A1(n_1265),
.A2(n_825),
.B1(n_857),
.B2(n_845),
.Y(n_1561)
);

CKINVDCx11_ASAP7_75t_R g1562 ( 
.A(n_1408),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1401),
.A2(n_1216),
.B1(n_825),
.B2(n_1346),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1414),
.B(n_1341),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1304),
.B(n_1306),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1281),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1281),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_SL g1568 ( 
.A1(n_1310),
.A2(n_1216),
.B1(n_825),
.B2(n_832),
.Y(n_1568)
);

CKINVDCx11_ASAP7_75t_R g1569 ( 
.A(n_1408),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1352),
.Y(n_1570)
);

INVx8_ASAP7_75t_L g1571 ( 
.A(n_1304),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1332),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1401),
.A2(n_1216),
.B1(n_825),
.B2(n_1346),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1333),
.A2(n_825),
.B1(n_1216),
.B2(n_832),
.Y(n_1574)
);

BUFx2_ASAP7_75t_SL g1575 ( 
.A(n_1402),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1295),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1333),
.A2(n_825),
.B1(n_1216),
.B2(n_832),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1401),
.A2(n_1216),
.B1(n_1346),
.B2(n_825),
.Y(n_1578)
);

INVx4_ASAP7_75t_L g1579 ( 
.A(n_1304),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1401),
.A2(n_919),
.B(n_584),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1401),
.A2(n_1216),
.B1(n_1346),
.B2(n_825),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1295),
.Y(n_1582)
);

CKINVDCx11_ASAP7_75t_R g1583 ( 
.A(n_1408),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1401),
.A2(n_1216),
.B1(n_1346),
.B2(n_825),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1401),
.A2(n_1216),
.B1(n_825),
.B2(n_1346),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1295),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1521),
.A2(n_1523),
.B(n_1520),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1511),
.B(n_1532),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1520),
.A2(n_1524),
.B(n_1519),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1522),
.A2(n_1534),
.B(n_1491),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1497),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1549),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1450),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1455),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1564),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1497),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1457),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1528),
.Y(n_1598)
);

OAI211xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1540),
.A2(n_1574),
.B(n_1577),
.C(n_1557),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1515),
.A2(n_1509),
.B(n_1530),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1561),
.A2(n_1540),
.B1(n_1577),
.B2(n_1574),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1568),
.A2(n_1544),
.B1(n_1464),
.B2(n_1517),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1549),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1435),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1442),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1512),
.Y(n_1606)
);

AO21x2_ASAP7_75t_L g1607 ( 
.A1(n_1510),
.A2(n_1476),
.B(n_1527),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1550),
.Y(n_1608)
);

INVx8_ASAP7_75t_L g1609 ( 
.A(n_1571),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1525),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1456),
.B(n_1548),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1441),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1550),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1533),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1536),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1446),
.B(n_1437),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1538),
.Y(n_1617)
);

AO21x2_ASAP7_75t_L g1618 ( 
.A1(n_1510),
.A2(n_1496),
.B(n_1495),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1461),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1538),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1487),
.A2(n_1508),
.B(n_1486),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1538),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1514),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1539),
.Y(n_1624)
);

OAI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1580),
.A2(n_1526),
.B1(n_1478),
.B2(n_1557),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1513),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1437),
.A2(n_1563),
.B(n_1585),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1446),
.B(n_1436),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1529),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1531),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1531),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1572),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1535),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1537),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1537),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1571),
.B(n_1504),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1452),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1485),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1573),
.A2(n_1584),
.B1(n_1581),
.B2(n_1556),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1576),
.Y(n_1640)
);

OR2x6_ASAP7_75t_L g1641 ( 
.A(n_1571),
.B(n_1484),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1582),
.B(n_1586),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1501),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1463),
.B(n_1500),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1436),
.B(n_1440),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1570),
.Y(n_1646)
);

NAND4xp25_ASAP7_75t_SL g1647 ( 
.A(n_1556),
.B(n_1584),
.C(n_1578),
.D(n_1581),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1466),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1448),
.B(n_1483),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1465),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1448),
.B(n_1483),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1471),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1486),
.A2(n_1518),
.B(n_1460),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1479),
.Y(n_1654)
);

BUFx2_ASAP7_75t_SL g1655 ( 
.A(n_1503),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1481),
.B(n_1490),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1445),
.Y(n_1657)
);

INVx5_ASAP7_75t_L g1658 ( 
.A(n_1439),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1503),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1439),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1578),
.A2(n_1458),
.B1(n_1477),
.B2(n_1470),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1488),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1473),
.Y(n_1663)
);

AOI21xp33_ASAP7_75t_L g1664 ( 
.A1(n_1458),
.A2(n_1477),
.B(n_1462),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1494),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1506),
.Y(n_1666)
);

OA21x2_ASAP7_75t_L g1667 ( 
.A1(n_1502),
.A2(n_1469),
.B(n_1567),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1545),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1575),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1443),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1559),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1566),
.Y(n_1672)
);

AOI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1505),
.A2(n_1499),
.B(n_1516),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1467),
.B(n_1507),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1467),
.B(n_1507),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1453),
.Y(n_1676)
);

OAI21x1_ASAP7_75t_SL g1677 ( 
.A1(n_1579),
.A2(n_1434),
.B(n_1480),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1493),
.Y(n_1678)
);

INVx8_ASAP7_75t_L g1679 ( 
.A(n_1444),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1507),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1553),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1565),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1542),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1551),
.A2(n_1489),
.B1(n_1443),
.B2(n_1482),
.Y(n_1684)
);

AO31x2_ASAP7_75t_L g1685 ( 
.A1(n_1565),
.A2(n_1541),
.A3(n_1447),
.B(n_1555),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1447),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1493),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1447),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1459),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1541),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1541),
.Y(n_1691)
);

AO21x1_ASAP7_75t_L g1692 ( 
.A1(n_1492),
.A2(n_1560),
.B(n_1555),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1560),
.Y(n_1693)
);

OA21x2_ASAP7_75t_L g1694 ( 
.A1(n_1492),
.A2(n_1474),
.B(n_1546),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1468),
.B(n_1498),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1468),
.B(n_1498),
.Y(n_1696)
);

BUFx2_ASAP7_75t_SL g1697 ( 
.A(n_1475),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1498),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1454),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1472),
.B(n_1547),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1451),
.A2(n_1543),
.B1(n_1554),
.B2(n_1449),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1662),
.B(n_1583),
.Y(n_1702)
);

NAND4xp25_ASAP7_75t_L g1703 ( 
.A(n_1601),
.B(n_1543),
.C(n_1554),
.D(n_1569),
.Y(n_1703)
);

OR2x6_ASAP7_75t_L g1704 ( 
.A(n_1636),
.B(n_1552),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1595),
.B(n_1562),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1602),
.A2(n_1451),
.B(n_1438),
.C(n_1558),
.Y(n_1706)
);

INVx2_ASAP7_75t_SL g1707 ( 
.A(n_1637),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1675),
.B(n_1656),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1675),
.B(n_1656),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1627),
.A2(n_1599),
.B(n_1664),
.C(n_1661),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1630),
.B(n_1631),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1625),
.A2(n_1647),
.B(n_1639),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1637),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1656),
.B(n_1603),
.Y(n_1714)
);

INVx4_ASAP7_75t_L g1715 ( 
.A(n_1658),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1603),
.B(n_1642),
.Y(n_1716)
);

AO32x2_ASAP7_75t_L g1717 ( 
.A1(n_1588),
.A2(n_1607),
.A3(n_1592),
.B1(n_1613),
.B2(n_1632),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1611),
.B(n_1683),
.Y(n_1718)
);

AO32x2_ASAP7_75t_L g1719 ( 
.A1(n_1588),
.A2(n_1607),
.A3(n_1608),
.B1(n_1633),
.B2(n_1626),
.Y(n_1719)
);

AO21x1_ASAP7_75t_L g1720 ( 
.A1(n_1645),
.A2(n_1644),
.B(n_1628),
.Y(n_1720)
);

A2O1A1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1628),
.A2(n_1645),
.B(n_1616),
.C(n_1649),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1616),
.A2(n_1648),
.B1(n_1649),
.B2(n_1651),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1654),
.B(n_1651),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1634),
.B(n_1635),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1634),
.B(n_1635),
.Y(n_1725)
);

BUFx4f_ASAP7_75t_SL g1726 ( 
.A(n_1646),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1654),
.B(n_1593),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_1612),
.Y(n_1728)
);

A2O1A1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1621),
.A2(n_1669),
.B(n_1674),
.C(n_1590),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1653),
.A2(n_1638),
.B1(n_1666),
.B2(n_1643),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1618),
.A2(n_1607),
.B1(n_1665),
.B2(n_1633),
.C(n_1604),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1614),
.B(n_1593),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1594),
.B(n_1597),
.Y(n_1733)
);

NAND3xp33_ASAP7_75t_L g1734 ( 
.A(n_1653),
.B(n_1667),
.C(n_1668),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1646),
.B(n_1700),
.Y(n_1735)
);

O2A1O1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1618),
.A2(n_1653),
.B(n_1677),
.C(n_1636),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1619),
.B(n_1624),
.Y(n_1737)
);

OAI211xp5_ASAP7_75t_SL g1738 ( 
.A1(n_1684),
.A2(n_1701),
.B(n_1670),
.C(n_1605),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1618),
.A2(n_1587),
.B(n_1589),
.Y(n_1739)
);

AOI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1653),
.A2(n_1636),
.B1(n_1667),
.B2(n_1695),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1667),
.A2(n_1636),
.B1(n_1680),
.B2(n_1687),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1697),
.A2(n_1678),
.B1(n_1687),
.B2(n_1658),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1640),
.A2(n_1650),
.B1(n_1652),
.B2(n_1672),
.C(n_1671),
.Y(n_1743)
);

INVx4_ASAP7_75t_L g1744 ( 
.A(n_1658),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1697),
.A2(n_1678),
.B1(n_1658),
.B2(n_1641),
.Y(n_1745)
);

A2O1A1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1659),
.A2(n_1695),
.B(n_1696),
.C(n_1658),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1700),
.B(n_1673),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1667),
.A2(n_1659),
.B1(n_1655),
.B2(n_1694),
.Y(n_1748)
);

BUFx4f_ASAP7_75t_SL g1749 ( 
.A(n_1699),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1598),
.Y(n_1750)
);

NOR2x1_ASAP7_75t_SL g1751 ( 
.A(n_1673),
.B(n_1626),
.Y(n_1751)
);

NOR2x1_ASAP7_75t_SL g1752 ( 
.A(n_1610),
.B(n_1591),
.Y(n_1752)
);

A2O1A1Ixp33_ASAP7_75t_L g1753 ( 
.A1(n_1659),
.A2(n_1696),
.B(n_1681),
.C(n_1682),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1596),
.B(n_1615),
.Y(n_1754)
);

OR2x6_ASAP7_75t_L g1755 ( 
.A(n_1692),
.B(n_1694),
.Y(n_1755)
);

AOI211xp5_ASAP7_75t_L g1756 ( 
.A1(n_1692),
.A2(n_1691),
.B(n_1686),
.C(n_1688),
.Y(n_1756)
);

OR2x6_ASAP7_75t_L g1757 ( 
.A(n_1694),
.B(n_1629),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1612),
.B(n_1699),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1663),
.B(n_1606),
.Y(n_1759)
);

AO21x2_ASAP7_75t_L g1760 ( 
.A1(n_1600),
.A2(n_1617),
.B(n_1622),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1657),
.Y(n_1761)
);

OA21x2_ASAP7_75t_L g1762 ( 
.A1(n_1617),
.A2(n_1620),
.B(n_1622),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_1757),
.Y(n_1763)
);

INVx4_ASAP7_75t_L g1764 ( 
.A(n_1704),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1750),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1762),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1723),
.B(n_1623),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1760),
.Y(n_1768)
);

INVxp67_ASAP7_75t_SL g1769 ( 
.A(n_1734),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1755),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1754),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1723),
.B(n_1623),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1717),
.B(n_1620),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1717),
.B(n_1676),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1717),
.B(n_1719),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1719),
.B(n_1739),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1719),
.B(n_1676),
.Y(n_1777)
);

INVxp67_ASAP7_75t_SL g1778 ( 
.A(n_1752),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1755),
.B(n_1685),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1755),
.B(n_1685),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1712),
.B(n_1698),
.C(n_1686),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1761),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1757),
.B(n_1693),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1712),
.A2(n_1679),
.B1(n_1641),
.B2(n_1693),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1727),
.B(n_1690),
.Y(n_1785)
);

AND2x4_ASAP7_75t_SL g1786 ( 
.A(n_1704),
.B(n_1641),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1759),
.Y(n_1787)
);

INVx8_ASAP7_75t_L g1788 ( 
.A(n_1704),
.Y(n_1788)
);

NOR2xp67_ASAP7_75t_L g1789 ( 
.A(n_1730),
.B(n_1688),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1737),
.B(n_1689),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1757),
.B(n_1685),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1733),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1767),
.B(n_1716),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1765),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1767),
.B(n_1772),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1781),
.A2(n_1710),
.B(n_1731),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1763),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1783),
.B(n_1791),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1784),
.A2(n_1721),
.B1(n_1706),
.B2(n_1747),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1788),
.Y(n_1800)
);

AOI33xp33_ASAP7_75t_L g1801 ( 
.A1(n_1776),
.A2(n_1732),
.A3(n_1748),
.B1(n_1708),
.B2(n_1709),
.B3(n_1756),
.Y(n_1801)
);

AND2x4_ASAP7_75t_SL g1802 ( 
.A(n_1764),
.B(n_1715),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1783),
.B(n_1740),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1772),
.B(n_1714),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1791),
.B(n_1711),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1783),
.B(n_1791),
.Y(n_1806)
);

BUFx3_ASAP7_75t_L g1807 ( 
.A(n_1788),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1765),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1790),
.B(n_1720),
.Y(n_1809)
);

INVx5_ASAP7_75t_L g1810 ( 
.A(n_1768),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1765),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1765),
.Y(n_1812)
);

NAND2x1_ASAP7_75t_L g1813 ( 
.A(n_1791),
.B(n_1744),
.Y(n_1813)
);

NOR3xp33_ASAP7_75t_L g1814 ( 
.A(n_1781),
.B(n_1738),
.C(n_1703),
.Y(n_1814)
);

AO21x2_ASAP7_75t_L g1815 ( 
.A1(n_1769),
.A2(n_1751),
.B(n_1729),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1788),
.A2(n_1703),
.B1(n_1722),
.B2(n_1711),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1791),
.B(n_1724),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1770),
.B(n_1792),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1770),
.B(n_1725),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1785),
.B(n_1722),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1777),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1771),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1788),
.A2(n_1764),
.B1(n_1784),
.B2(n_1786),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1789),
.A2(n_1741),
.B1(n_1726),
.B2(n_1736),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1764),
.B(n_1735),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1770),
.B(n_1725),
.Y(n_1826)
);

OAI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1769),
.A2(n_1746),
.B1(n_1736),
.B2(n_1753),
.C(n_1718),
.Y(n_1827)
);

AOI33xp33_ASAP7_75t_L g1828 ( 
.A1(n_1776),
.A2(n_1724),
.A3(n_1743),
.B1(n_1702),
.B2(n_1707),
.B3(n_1713),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1782),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1794),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1821),
.B(n_1776),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1794),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1811),
.Y(n_1833)
);

NOR2x1_ASAP7_75t_L g1834 ( 
.A(n_1796),
.B(n_1815),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1809),
.B(n_1787),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1802),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1811),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1821),
.B(n_1775),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1808),
.Y(n_1839)
);

NAND2x1_ASAP7_75t_L g1840 ( 
.A(n_1797),
.B(n_1775),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1812),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1812),
.Y(n_1842)
);

BUFx2_ASAP7_75t_L g1843 ( 
.A(n_1815),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1821),
.B(n_1798),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1808),
.B(n_1766),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1798),
.B(n_1806),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1810),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1806),
.B(n_1775),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1818),
.B(n_1763),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1818),
.B(n_1763),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1802),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1803),
.B(n_1763),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1803),
.B(n_1773),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1822),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1797),
.B(n_1773),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1829),
.B(n_1766),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1805),
.B(n_1773),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1805),
.B(n_1774),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1805),
.B(n_1774),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1813),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1815),
.B(n_1777),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1817),
.B(n_1777),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1810),
.B(n_1779),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1854),
.Y(n_1864)
);

INVxp67_ASAP7_75t_SL g1865 ( 
.A(n_1834),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1835),
.B(n_1820),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1854),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1830),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1830),
.Y(n_1869)
);

NAND2x1p5_ASAP7_75t_L g1870 ( 
.A(n_1834),
.B(n_1764),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1830),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1835),
.B(n_1793),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1834),
.B(n_1828),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1832),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1832),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1853),
.B(n_1793),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1832),
.Y(n_1877)
);

AND2x4_ASAP7_75t_SL g1878 ( 
.A(n_1860),
.B(n_1764),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1833),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1852),
.B(n_1817),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1845),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1833),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1833),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1837),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1837),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1852),
.B(n_1796),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1837),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1853),
.B(n_1804),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1841),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1841),
.Y(n_1890)
);

INVxp33_ASAP7_75t_L g1891 ( 
.A(n_1852),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1843),
.A2(n_1814),
.B1(n_1799),
.B2(n_1827),
.Y(n_1892)
);

AOI32xp33_ASAP7_75t_L g1893 ( 
.A1(n_1861),
.A2(n_1824),
.A3(n_1816),
.B1(n_1819),
.B2(n_1826),
.Y(n_1893)
);

AND2x4_ASAP7_75t_SL g1894 ( 
.A(n_1860),
.B(n_1819),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1841),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1846),
.B(n_1826),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1861),
.B(n_1801),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1836),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1853),
.B(n_1804),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1845),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1836),
.B(n_1851),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1848),
.B(n_1795),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1845),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1842),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1842),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1843),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1836),
.B(n_1807),
.Y(n_1907)
);

INVx2_ASAP7_75t_SL g1908 ( 
.A(n_1836),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1851),
.Y(n_1909)
);

NAND3xp33_ASAP7_75t_L g1910 ( 
.A(n_1892),
.B(n_1843),
.C(n_1861),
.Y(n_1910)
);

INVx1_ASAP7_75t_SL g1911 ( 
.A(n_1901),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1894),
.B(n_1846),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1894),
.B(n_1901),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1901),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1892),
.B(n_1897),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1881),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1880),
.B(n_1846),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1864),
.B(n_1840),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1907),
.B(n_1846),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1907),
.B(n_1857),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1867),
.B(n_1840),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1865),
.B(n_1847),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1907),
.B(n_1857),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1896),
.B(n_1857),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1872),
.B(n_1840),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1886),
.B(n_1855),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1868),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1881),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1876),
.B(n_1848),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1866),
.B(n_1873),
.Y(n_1930)
);

NOR2x1p5_ASAP7_75t_L g1931 ( 
.A(n_1865),
.B(n_1851),
.Y(n_1931)
);

AOI211xp5_ASAP7_75t_L g1932 ( 
.A1(n_1891),
.A2(n_1824),
.B(n_1789),
.C(n_1742),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1870),
.B(n_1858),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1869),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1888),
.B(n_1848),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1900),
.B(n_1855),
.Y(n_1936)
);

NAND2x1p5_ASAP7_75t_L g1937 ( 
.A(n_1909),
.B(n_1851),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1900),
.B(n_1855),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1870),
.A2(n_1891),
.B(n_1906),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1898),
.B(n_1858),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1898),
.B(n_1858),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1908),
.B(n_1859),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1871),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1906),
.Y(n_1944)
);

NAND2xp33_ASAP7_75t_SL g1945 ( 
.A(n_1908),
.B(n_1728),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1874),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1875),
.Y(n_1947)
);

OAI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1910),
.A2(n_1915),
.B1(n_1930),
.B2(n_1911),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1922),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1913),
.B(n_1909),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1922),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1937),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1915),
.B(n_1893),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1922),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1910),
.A2(n_1932),
.B1(n_1914),
.B2(n_1911),
.Y(n_1955)
);

INVxp67_ASAP7_75t_L g1956 ( 
.A(n_1914),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1930),
.B(n_1899),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1946),
.Y(n_1958)
);

AOI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1932),
.A2(n_1903),
.B1(n_1904),
.B2(n_1905),
.C(n_1877),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1922),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1946),
.Y(n_1961)
);

AOI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1945),
.A2(n_1878),
.B1(n_1825),
.B2(n_1823),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1926),
.B(n_1902),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1939),
.A2(n_1926),
.B(n_1944),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1944),
.Y(n_1965)
);

OAI32xp33_ASAP7_75t_L g1966 ( 
.A1(n_1939),
.A2(n_1847),
.A3(n_1863),
.B1(n_1780),
.B2(n_1779),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1927),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1929),
.B(n_1903),
.Y(n_1968)
);

AND2x2_ASAP7_75t_SL g1969 ( 
.A(n_1913),
.B(n_1786),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1931),
.A2(n_1878),
.B1(n_1779),
.B2(n_1780),
.Y(n_1970)
);

AOI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1936),
.A2(n_1895),
.B1(n_1890),
.B2(n_1889),
.C(n_1887),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1919),
.B(n_1920),
.Y(n_1972)
);

AOI322xp5_ASAP7_75t_L g1973 ( 
.A1(n_1919),
.A2(n_1838),
.A3(n_1831),
.B1(n_1844),
.B2(n_1862),
.C1(n_1863),
.C2(n_1859),
.Y(n_1973)
);

INVxp67_ASAP7_75t_SL g1974 ( 
.A(n_1931),
.Y(n_1974)
);

OAI221xp5_ASAP7_75t_L g1975 ( 
.A1(n_1953),
.A2(n_1937),
.B1(n_1936),
.B2(n_1938),
.C(n_1925),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1974),
.B(n_1758),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1965),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1958),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1956),
.B(n_1917),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1969),
.B(n_1937),
.Y(n_1980)
);

OAI21xp33_ASAP7_75t_L g1981 ( 
.A1(n_1955),
.A2(n_1941),
.B(n_1940),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1972),
.B(n_1920),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1952),
.Y(n_1983)
);

OAI21xp33_ASAP7_75t_L g1984 ( 
.A1(n_1959),
.A2(n_1941),
.B(n_1940),
.Y(n_1984)
);

OAI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1948),
.A2(n_1937),
.B1(n_1929),
.B2(n_1935),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1961),
.Y(n_1986)
);

INVx1_ASAP7_75t_SL g1987 ( 
.A(n_1950),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1964),
.B(n_1950),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1952),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1972),
.B(n_1923),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1967),
.Y(n_1991)
);

OAI32xp33_ASAP7_75t_L g1992 ( 
.A1(n_1949),
.A2(n_1918),
.A3(n_1921),
.B1(n_1925),
.B2(n_1938),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1969),
.B(n_1923),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1949),
.B(n_1917),
.Y(n_1994)
);

O2A1O1Ixp5_ASAP7_75t_L g1995 ( 
.A1(n_1966),
.A2(n_1916),
.B(n_1928),
.C(n_1933),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1982),
.B(n_1962),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1987),
.B(n_1951),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1982),
.B(n_1951),
.Y(n_1998)
);

NAND3xp33_ASAP7_75t_L g1999 ( 
.A(n_1985),
.B(n_1971),
.C(n_1960),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1983),
.Y(n_2000)
);

OAI32xp33_ASAP7_75t_L g2001 ( 
.A1(n_1988),
.A2(n_1960),
.A3(n_1954),
.B1(n_1921),
.B2(n_1918),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1983),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1979),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1976),
.B(n_1954),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1977),
.Y(n_2005)
);

AOI221xp5_ASAP7_75t_L g2006 ( 
.A1(n_1992),
.A2(n_1966),
.B1(n_1970),
.B2(n_1957),
.C(n_1968),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1977),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1978),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_2000),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1998),
.B(n_1990),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_2000),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_2004),
.B(n_1993),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_2003),
.B(n_1993),
.Y(n_2013)
);

OAI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1999),
.A2(n_1995),
.B(n_1980),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_2006),
.B(n_1981),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1998),
.B(n_1990),
.Y(n_2016)
);

AOI221xp5_ASAP7_75t_L g2017 ( 
.A1(n_2001),
.A2(n_1992),
.B1(n_1975),
.B2(n_1984),
.C(n_1986),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_2002),
.Y(n_2018)
);

NAND3xp33_ASAP7_75t_L g2019 ( 
.A(n_1997),
.B(n_1986),
.C(n_1978),
.Y(n_2019)
);

OAI211xp5_ASAP7_75t_L g2020 ( 
.A1(n_2014),
.A2(n_2002),
.B(n_2007),
.C(n_2005),
.Y(n_2020)
);

AOI221xp5_ASAP7_75t_L g2021 ( 
.A1(n_2015),
.A2(n_1996),
.B1(n_2008),
.B2(n_1991),
.C(n_1994),
.Y(n_2021)
);

AOI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_2017),
.A2(n_1989),
.B1(n_1916),
.B2(n_1928),
.C(n_1968),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_2012),
.B(n_2010),
.Y(n_2023)
);

AOI321xp33_ASAP7_75t_L g2024 ( 
.A1(n_2013),
.A2(n_1989),
.A3(n_1928),
.B1(n_1916),
.B2(n_1963),
.C(n_1933),
.Y(n_2024)
);

AOI221xp5_ASAP7_75t_SL g2025 ( 
.A1(n_2016),
.A2(n_1933),
.B1(n_1934),
.B2(n_1927),
.C(n_1947),
.Y(n_2025)
);

AOI222xp33_ASAP7_75t_L g2026 ( 
.A1(n_2020),
.A2(n_2019),
.B1(n_2011),
.B2(n_2009),
.C1(n_2018),
.C2(n_1943),
.Y(n_2026)
);

INVxp67_ASAP7_75t_SL g2027 ( 
.A(n_2023),
.Y(n_2027)
);

AOI211xp5_ASAP7_75t_L g2028 ( 
.A1(n_2022),
.A2(n_1963),
.B(n_1934),
.C(n_1943),
.Y(n_2028)
);

AOI321xp33_ASAP7_75t_L g2029 ( 
.A1(n_2021),
.A2(n_1942),
.A3(n_1912),
.B1(n_1947),
.B2(n_1705),
.C(n_1924),
.Y(n_2029)
);

AOI221xp5_ASAP7_75t_L g2030 ( 
.A1(n_2025),
.A2(n_1942),
.B1(n_1912),
.B2(n_1847),
.C(n_1924),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_2024),
.Y(n_2031)
);

OAI211xp5_ASAP7_75t_L g2032 ( 
.A1(n_2020),
.A2(n_1973),
.B(n_1679),
.C(n_1847),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2027),
.Y(n_2033)
);

NOR2x1_ASAP7_75t_L g2034 ( 
.A(n_2032),
.B(n_1860),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_2031),
.Y(n_2035)
);

XOR2xp5_ASAP7_75t_L g2036 ( 
.A(n_2029),
.B(n_2026),
.Y(n_2036)
);

XNOR2x1_ASAP7_75t_L g2037 ( 
.A(n_2028),
.B(n_1641),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2030),
.Y(n_2038)
);

AOI21xp33_ASAP7_75t_SL g2039 ( 
.A1(n_2035),
.A2(n_1679),
.B(n_1935),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_2033),
.B(n_1860),
.Y(n_2040)
);

AOI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_2036),
.A2(n_1885),
.B1(n_1884),
.B2(n_1883),
.C(n_1882),
.Y(n_2041)
);

OAI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_2037),
.A2(n_1860),
.B(n_1879),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2040),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_2043),
.A2(n_2038),
.B1(n_2034),
.B2(n_2041),
.Y(n_2044)
);

OA21x2_ASAP7_75t_L g2045 ( 
.A1(n_2044),
.A2(n_2042),
.B(n_2039),
.Y(n_2045)
);

NOR2x1p5_ASAP7_75t_L g2046 ( 
.A(n_2044),
.B(n_1749),
.Y(n_2046)
);

XOR2xp5_ASAP7_75t_L g2047 ( 
.A(n_2045),
.B(n_1800),
.Y(n_2047)
);

OAI22x1_ASAP7_75t_L g2048 ( 
.A1(n_2046),
.A2(n_1860),
.B1(n_1863),
.B2(n_1778),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_2048),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_2047),
.A2(n_1863),
.B1(n_1849),
.B2(n_1850),
.Y(n_2050)
);

OAI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_2049),
.A2(n_1856),
.B1(n_1839),
.B2(n_1810),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_2051),
.A2(n_2050),
.B(n_1839),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_2052),
.Y(n_2053)
);

OAI221xp5_ASAP7_75t_R g2054 ( 
.A1(n_2053),
.A2(n_1788),
.B1(n_1609),
.B2(n_1856),
.C(n_1810),
.Y(n_2054)
);

AOI211xp5_ASAP7_75t_L g2055 ( 
.A1(n_2054),
.A2(n_1742),
.B(n_1745),
.C(n_1660),
.Y(n_2055)
);


endmodule