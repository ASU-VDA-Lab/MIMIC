module fake_jpeg_8932_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_2),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_0),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_1),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

OR2x2_ASAP7_75t_SL g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

OA22x2_ASAP7_75t_SL g27 ( 
.A1(n_17),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_26),
.B(n_24),
.C(n_15),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_13),
.B1(n_14),
.B2(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_5),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_32),
.B1(n_23),
.B2(n_11),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_11),
.C(n_16),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_39),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_6),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_32),
.B(n_11),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_36),
.B(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_44),
.B(n_41),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_43),
.C(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_46),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.C(n_16),
.Y(n_53)
);

OAI21x1_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_7),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_7),
.Y(n_55)
);


endmodule