module fake_jpeg_27556_n_118 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_118);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_17),
.Y(n_52)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_12),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_26),
.B(n_13),
.Y(n_50)
);

AND2x6_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_51),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_30),
.B1(n_20),
.B2(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_18),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_14),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_27),
.B1(n_29),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_20),
.B1(n_25),
.B2(n_29),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_36),
.B1(n_39),
.B2(n_14),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_35),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_50),
.C(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_55),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_11),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_15),
.Y(n_84)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_34),
.B1(n_32),
.B2(n_11),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_63),
.B1(n_51),
.B2(n_42),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_17),
.B1(n_22),
.B2(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_67),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_15),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_31),
.C(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_38),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_63),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_31),
.B(n_19),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_64),
.B(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_12),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_72),
.B(n_59),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_92),
.B(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_56),
.B(n_2),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_56),
.B1(n_77),
.B2(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_100),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_94),
.B1(n_85),
.B2(n_90),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_76),
.B1(n_84),
.B2(n_15),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_104),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_100),
.B(n_102),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_99),
.B(n_3),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_99),
.B(n_2),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_4),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_1),
.B(n_3),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_110),
.B(n_9),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_3),
.B1(n_4),
.B2(n_9),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_114),
.B(n_10),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_116),
.B(n_10),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_10),
.Y(n_118)
);


endmodule