module fake_jpeg_6155_n_291 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_291);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_30),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_18),
.B1(n_15),
.B2(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_20),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_36),
.Y(n_43)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_18),
.B1(n_16),
.B2(n_26),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_16),
.B1(n_26),
.B2(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_20),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_54),
.Y(n_63)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_60),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_17),
.B1(n_43),
.B2(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

XOR2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_19),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_28),
.A3(n_17),
.B1(n_20),
.B2(n_15),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_37),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_24),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_73),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_29),
.B(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_35),
.B1(n_28),
.B2(n_18),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_51),
.B1(n_17),
.B2(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_50),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_75),
.A2(n_38),
.B1(n_40),
.B2(n_50),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_56),
.B1(n_76),
.B2(n_64),
.Y(n_103)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_83),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_40),
.B1(n_50),
.B2(n_35),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_82),
.A2(n_45),
.B1(n_54),
.B2(n_60),
.Y(n_120)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_14),
.Y(n_114)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_88),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_67),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_93),
.B1(n_96),
.B2(n_56),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_94),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_63),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_35),
.B1(n_43),
.B2(n_31),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_95),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_37),
.B(n_51),
.C(n_19),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_31),
.B1(n_45),
.B2(n_49),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_98),
.B1(n_56),
.B2(n_57),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_72),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_81),
.C(n_85),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_110),
.B1(n_112),
.B2(n_119),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_R g106 ( 
.A(n_92),
.B(n_72),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_86),
.B1(n_89),
.B2(n_96),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_59),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_70),
.B1(n_55),
.B2(n_45),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_88),
.B1(n_84),
.B2(n_77),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_51),
.B1(n_31),
.B2(n_52),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_96),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_29),
.A3(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_116),
.B(n_117),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_63),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_64),
.B1(n_57),
.B2(n_58),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_97),
.B1(n_84),
.B2(n_77),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_29),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_131),
.C(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_138),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_145),
.B(n_132),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_86),
.C(n_91),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_104),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_139),
.B1(n_99),
.B2(n_79),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_114),
.B(n_117),
.C(n_115),
.D(n_110),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_88),
.B1(n_79),
.B2(n_14),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_78),
.B1(n_54),
.B2(n_66),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_143),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_141),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_14),
.A3(n_21),
.B1(n_23),
.B2(n_13),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_29),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_32),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_138),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_144),
.A2(n_116),
.B(n_117),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_152),
.B(n_157),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_153),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_158),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_134),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_155),
.Y(n_185)
);

XOR2x2_ASAP7_75t_SL g183 ( 
.A(n_156),
.B(n_34),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_113),
.B(n_105),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_164),
.B1(n_139),
.B2(n_129),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_160),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_88),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_169),
.B1(n_128),
.B2(n_14),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_127),
.B1(n_141),
.B2(n_126),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_131),
.C(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_170),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_151),
.A2(n_130),
.B1(n_124),
.B2(n_123),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_188),
.C(n_163),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_135),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_180),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_140),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_189),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_158),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_157),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_186),
.Y(n_213)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_32),
.C(n_33),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_33),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_95),
.B1(n_69),
.B2(n_21),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_171),
.A2(n_168),
.B(n_147),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_203),
.B1(n_191),
.B2(n_186),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_201),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_189),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_146),
.B(n_155),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_207),
.C(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_162),
.C(n_160),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_161),
.B(n_156),
.C(n_146),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_209),
.A2(n_178),
.B1(n_185),
.B2(n_190),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_193),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_210),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_164),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_180),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_224),
.C(n_225),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_222),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_225),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_223),
.C(n_200),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_188),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_181),
.C(n_173),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_175),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_174),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_196),
.B1(n_199),
.B2(n_198),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_195),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_227),
.B(n_230),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_172),
.B1(n_184),
.B2(n_157),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_203),
.B1(n_212),
.B2(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_159),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_231),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_23),
.C(n_13),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_221),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_202),
.B1(n_95),
.B2(n_21),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_1),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_12),
.B(n_2),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_243),
.A2(n_12),
.B(n_229),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_13),
.C(n_23),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_245),
.C(n_228),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_13),
.C(n_23),
.Y(n_245)
);

FAx1_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_1),
.CI(n_2),
.CON(n_246),
.SN(n_246)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_27),
.B(n_12),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_250),
.B(n_251),
.Y(n_262)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_247),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_259),
.C(n_4),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_235),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_257),
.Y(n_270)
);

AOI21x1_ASAP7_75t_SL g265 ( 
.A1(n_254),
.A2(n_255),
.B(n_1),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_23),
.C(n_3),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_13),
.C(n_3),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_5),
.C(n_6),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_23),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_246),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_1),
.C(n_3),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_238),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_265),
.B(n_267),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_245),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_SL g274 ( 
.A(n_263),
.B(n_260),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_268),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_271),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_13),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_4),
.Y(n_268)
);

AOI321xp33_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_265),
.A3(n_271),
.B1(n_9),
.B2(n_10),
.C(n_7),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_5),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_275),
.B(n_278),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_279),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_6),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_7),
.Y(n_279)
);

A2O1A1O1Ixp25_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_273),
.B(n_280),
.C(n_10),
.D(n_8),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g283 ( 
.A(n_276),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_284),
.C(n_272),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_7),
.B(n_8),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_282),
.B(n_286),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_8),
.B(n_9),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_9),
.C(n_10),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_290),
.A2(n_9),
.B(n_10),
.Y(n_291)
);


endmodule