module real_jpeg_7191_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_1),
.A2(n_24),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_44),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_2),
.A2(n_44),
.B1(n_82),
.B2(n_86),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_2),
.A2(n_44),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_2),
.A2(n_199),
.B(n_202),
.C(n_205),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_22),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_2),
.B(n_67),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_2),
.B(n_242),
.C(n_245),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_2),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_2),
.B(n_239),
.C(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_2),
.B(n_121),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_3),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_3),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_77),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_3),
.A2(n_77),
.B1(n_125),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_3),
.A2(n_77),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_4),
.Y(n_158)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_6),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_6),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_7),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_7),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_8),
.Y(n_128)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_8),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_8),
.Y(n_201)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_10),
.Y(n_141)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_215),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_213),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_187),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_15),
.B(n_187),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_143),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_79),
.C(n_115),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_18),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_49),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_19),
.A2(n_49),
.B1(n_237),
.B2(n_314),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_19),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_23),
.B(n_32),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_20),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_23),
.Y(n_153)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_27),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_28),
.Y(n_161)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_42),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_33),
.A2(n_153),
.B1(n_154),
.B2(n_162),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_33),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_34),
.A2(n_43),
.B1(n_208),
.B2(n_211),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_34),
.A2(n_43),
.B1(n_208),
.B2(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_36),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_41),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_43),
.B(n_183),
.Y(n_272)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_44),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_49),
.A2(n_237),
.B1(n_238),
.B2(n_247),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_49),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_49),
.A2(n_165),
.B1(n_166),
.B2(n_237),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_72),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_50),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_51),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_51),
.B(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_53),
.Y(n_240)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_56),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_67),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_61),
.Y(n_244)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_64),
.Y(n_177)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_66),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_67),
.A2(n_175),
.B(n_181),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_79),
.A2(n_115),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_79),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_89),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_81),
.A2(n_90),
.B1(n_106),
.B2(n_167),
.Y(n_166)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_81),
.A2(n_90),
.B1(n_106),
.B2(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_85),
.Y(n_170)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_106),
.Y(n_89)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_106),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_96),
.B1(n_101),
.B2(n_103),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_99),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_100),
.Y(n_266)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_102),
.Y(n_271)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_106),
.Y(n_254)
);

AOI22x1_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_115),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_115),
.A2(n_191),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_115),
.B(n_166),
.C(n_297),
.Y(n_315)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_120),
.B1(n_137),
.B2(n_142),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_120),
.B1(n_137),
.B2(n_142),
.Y(n_164)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_129),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_127),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_130),
.B1(n_132),
.B2(n_134),
.Y(n_129)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g203 ( 
.A(n_124),
.Y(n_203)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_172),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_163),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_152),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_147),
.B1(n_152),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_146),
.A2(n_147),
.B1(n_253),
.B2(n_255),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_146),
.A2(n_147),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_147),
.B(n_207),
.C(n_253),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_147),
.B(n_279),
.C(n_281),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_149),
.B(n_150),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_171),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_164),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_196),
.C(n_197),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_164),
.A2(n_171),
.B1(n_196),
.B2(n_287),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_165),
.B(n_237),
.C(n_261),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_165),
.A2(n_166),
.B1(n_297),
.B2(n_299),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_182),
.B2(n_186),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.C(n_195),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_188),
.A2(n_189),
.B1(n_193),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_193),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_195),
.B(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_196),
.A2(n_283),
.B1(n_284),
.B2(n_287),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_196),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_197),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_206),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_198),
.A2(n_206),
.B1(n_207),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_198),
.Y(n_305)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_207),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_232),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_210),
.Y(n_225)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_307),
.B(n_323),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_291),
.B(n_306),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_276),
.B(n_290),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_258),
.B(n_275),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_249),
.B(n_257),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_234),
.B(n_248),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_231),
.B(n_233),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_227),
.A2(n_235),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_236),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_235),
.B(n_285),
.C(n_287),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_247),
.Y(n_256)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_256),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_256),
.Y(n_257)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_253),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_260),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_274),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_272),
.B2(n_273),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_273),
.Y(n_279)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_289),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_289),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_281),
.B1(n_282),
.B2(n_288),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_279),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_293),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_300),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_302),
.C(n_303),
.Y(n_316)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_316),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_315),
.C(n_319),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_324),
.B(n_325),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_320),
.Y(n_325)
);


endmodule