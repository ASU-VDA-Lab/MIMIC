module real_jpeg_7512_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_286;
wire n_166;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_534;
wire n_181;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_0),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_0),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_0),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_0),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_0),
.B(n_164),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_0),
.B(n_346),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_0),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_0),
.B(n_442),
.Y(n_441)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_1),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_1),
.Y(n_176)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_1),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_1),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_1),
.Y(n_305)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_2),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_2),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_2),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_4),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_4),
.B(n_40),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_4),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_4),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_4),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_4),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_5),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_5),
.B(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_5),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_5),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_5),
.B(n_360),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_5),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_6),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_6),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_6),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_6),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_6),
.B(n_204),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_6),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_6),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_7),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_7),
.B(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_7),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_7),
.B(n_231),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_7),
.B(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_7),
.B(n_458),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_7),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_7),
.B(n_58),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_8),
.Y(n_116)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_8),
.Y(n_493)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g304 ( 
.A(n_10),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_10),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_10),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_10),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_10),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_10),
.B(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_11),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_11),
.Y(n_452)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_13),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_13),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_14),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_14),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g370 ( 
.A(n_14),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_14),
.B(n_451),
.Y(n_450)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_16),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_16),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_16),
.B(n_231),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_16),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_16),
.B(n_401),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_16),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_16),
.B(n_492),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_17),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_17),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_17),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_17),
.B(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_17),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_17),
.B(n_154),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_17),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_17),
.B(n_418),
.Y(n_417)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_19),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_19),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_19),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_19),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_19),
.B(n_231),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_19),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_19),
.B(n_42),
.Y(n_301)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_36),
.B(n_85),
.C(n_548),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_51),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_29),
.B(n_51),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_44),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_31),
.A2(n_32),
.B1(n_45),
.B2(n_66),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_45),
.C(n_49),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_33),
.B(n_394),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_34),
.B(n_169),
.Y(n_455)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_35),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_55),
.C(n_62),
.Y(n_82)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_47),
.Y(n_484)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_47),
.Y(n_509)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_48),
.Y(n_156)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_48),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_50),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_81),
.C(n_83),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_52),
.B(n_538),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_67),
.C(n_71),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_53),
.A2(n_54),
.B1(n_534),
.B2(n_535),
.Y(n_533)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_59),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_72),
.C(n_76),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_61),
.A2(n_62),
.B1(n_76),
.B2(n_494),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_65),
.Y(n_267)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_65),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_67),
.B(n_71),
.Y(n_535)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_72),
.A2(n_73),
.B1(n_496),
.B2(n_497),
.Y(n_495)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_76),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_76),
.A2(n_449),
.B1(n_450),
.B2(n_494),
.Y(n_513)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_78),
.Y(n_235)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_79),
.Y(n_264)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_79),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_79),
.Y(n_405)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_79),
.Y(n_463)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_539),
.Y(n_538)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_83),
.Y(n_539)
);

AO21x1_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_467),
.B(n_541),
.Y(n_85)
);

OAI21x1_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_428),
.B(n_466),
.Y(n_86)
);

AOI21x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_381),
.B(n_427),
.Y(n_87)
);

OAI21x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_332),
.B(n_380),
.Y(n_88)
);

AOI21x1_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_294),
.B(n_331),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_215),
.B(n_293),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_195),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_92),
.B(n_195),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_137),
.B2(n_194),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_93),
.B(n_138),
.C(n_177),
.Y(n_330)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_117),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_95),
.B(n_118),
.C(n_136),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_109),
.C(n_113),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_96),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_97),
.A2(n_98),
.B1(n_103),
.B2(n_104),
.Y(n_200)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_102),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_102),
.Y(n_396)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_108),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_109),
.B(n_113),
.Y(n_214)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_111),
.Y(n_447)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_116),
.Y(n_324)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_116),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_125),
.B1(n_135),
.B2(n_136),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B(n_124),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_120),
.Y(n_124)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_124),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_124),
.B(n_299),
.C(n_310),
.Y(n_339)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_126),
.B(n_128),
.C(n_131),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_137),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_177),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_150),
.C(n_167),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_139),
.B(n_197),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g551 ( 
.A(n_139),
.Y(n_551)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_143),
.CI(n_147),
.CON(n_139),
.SN(n_139)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_143),
.C(n_147),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_146),
.Y(n_205)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_146),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_149),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_150),
.A2(n_151),
.B1(n_167),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.C(n_162),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_152),
.A2(n_153),
.B1(n_162),
.B2(n_163),
.Y(n_286)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_156),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_157),
.B(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_165),
.Y(n_458)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_173),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_169),
.B(n_476),
.Y(n_475)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_172),
.Y(n_308)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_176),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_191),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_178),
.B(n_192),
.C(n_193),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g310 ( 
.A(n_179),
.B(n_186),
.C(n_189),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.C(n_213),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_196),
.B(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_199),
.B(n_213),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.C(n_206),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_200),
.B(n_201),
.Y(n_279)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_206),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_211),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_207),
.B(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_288),
.B(n_292),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_273),
.B(n_287),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_255),
.B(n_272),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_244),
.B(n_254),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_227),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_227),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_224),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_223),
.Y(n_369)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_236),
.B2(n_237),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_232),
.C(n_236),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_242),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_249),
.B(n_253),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_247),
.Y(n_253)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_248),
.Y(n_408)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_271),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_271),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_259),
.C(n_275),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_268),
.C(n_270),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_267),
.Y(n_402)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_276),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_283),
.C(n_284),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_290),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_330),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_330),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_312),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_298),
.C(n_312),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_309),
.B2(n_311),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_304),
.C(n_306),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_315),
.C(n_325),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_325),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_321),
.C(n_322),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_328),
.C(n_329),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_334),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_335),
.B(n_352),
.C(n_378),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_352),
.B1(n_378),
.B2(n_379),
.Y(n_336)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_340),
.B2(n_351),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_341),
.C(n_342),
.Y(n_383)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_340),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_350),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_344),
.B(n_345),
.C(n_350),
.Y(n_414)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_352),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_363),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_364),
.C(n_365),
.Y(n_412)
);

BUFx24_ASAP7_75t_SL g553 ( 
.A(n_353),
.Y(n_553)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_357),
.CI(n_359),
.CON(n_353),
.SN(n_353)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_354),
.B(n_357),
.C(n_359),
.Y(n_424)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_374),
.B2(n_375),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_370),
.B1(n_372),
.B2(n_373),
.Y(n_367)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_368),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_373),
.C(n_374),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_370),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_370),
.A2(n_373),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_373),
.B(n_388),
.C(n_393),
.Y(n_439)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_426),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_426),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_383),
.B(n_385),
.C(n_410),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_410),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_397),
.B2(n_409),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_398),
.C(n_399),
.Y(n_433)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_392),
.A2(n_393),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_392),
.B(n_446),
.C(n_449),
.Y(n_514)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_397),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_399),
.B(n_454),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_399),
.B(n_445),
.C(n_454),
.Y(n_473)
);

FAx1_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_403),
.CI(n_406),
.CON(n_399),
.SN(n_399)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_412),
.B1(n_413),
.B2(n_425),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_414),
.C(n_415),
.Y(n_430)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_424),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_419),
.B1(n_422),
.B2(n_423),
.Y(n_416)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_417),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_419),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_422),
.C(n_437),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_419),
.A2(n_423),
.B1(n_441),
.B2(n_443),
.Y(n_440)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_439),
.C(n_443),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_424),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_465),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_465),
.Y(n_466)
);

BUFx24_ASAP7_75t_SL g552 ( 
.A(n_429),
.Y(n_552)
);

FAx1_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.CI(n_444),
.CON(n_429),
.SN(n_429)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_430),
.B(n_431),
.C(n_444),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_434),
.B2(n_435),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_432),
.B(n_436),
.C(n_438),
.Y(n_522)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_438),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_441),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_453),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_449),
.B(n_491),
.C(n_494),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_455),
.B(n_459),
.C(n_464),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_459),
.B1(n_460),
.B2(n_464),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_457),
.Y(n_464)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

NOR3xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_526),
.C(n_536),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_523),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_470),
.A2(n_545),
.B(n_546),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_516),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_471),
.B(n_516),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_487),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_472),
.B(n_488),
.C(n_511),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.C(n_485),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_473),
.B(n_518),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_474),
.A2(n_485),
.B1(n_486),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_474),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_477),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_478),
.C(n_481),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_481),
.Y(n_477)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_511),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_500),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_495),
.B1(n_498),
.B2(n_499),
.Y(n_489)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_490),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_490),
.B(n_499),
.C(n_500),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_513),
.Y(n_512)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_495),
.Y(n_499)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_501),
.B(n_504),
.C(n_510),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_505),
.B2(n_510),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_503),
.Y(n_510)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_514),
.C(n_515),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_521),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_515),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.C(n_522),
.Y(n_516)
);

FAx1_ASAP7_75t_SL g524 ( 
.A(n_517),
.B(n_520),
.CI(n_522),
.CON(n_524),
.SN(n_524)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_525),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_524),
.B(n_525),
.Y(n_545)
);

BUFx24_ASAP7_75t_SL g550 ( 
.A(n_524),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_544),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_529),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_531),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_532),
.C(n_533),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_533),
.Y(n_531)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

A2O1A1Ixp33_ASAP7_75t_L g541 ( 
.A1(n_536),
.A2(n_542),
.B(n_543),
.C(n_547),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_540),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_537),
.B(n_540),
.Y(n_547)
);


endmodule