module real_aes_15604_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1694;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_1712;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1699;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1280;
wire n_729;
wire n_394;
wire n_1323;
wire n_1352;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_1705;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1344 ( .A(n_0), .Y(n_1344) );
OAI211xp5_ASAP7_75t_L g452 ( .A1(n_1), .A2(n_443), .B(n_453), .C(n_457), .Y(n_452) );
INVx1_ASAP7_75t_L g503 ( .A(n_1), .Y(n_503) );
INVx1_ASAP7_75t_L g652 ( .A(n_2), .Y(n_652) );
OAI211xp5_ASAP7_75t_L g698 ( .A1(n_2), .A2(n_699), .B(n_701), .C(n_710), .Y(n_698) );
INVx1_ASAP7_75t_L g326 ( .A(n_3), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_3), .B(n_336), .Y(n_351) );
AND2x2_ASAP7_75t_L g535 ( .A(n_3), .B(n_482), .Y(n_535) );
AND2x2_ASAP7_75t_L g602 ( .A(n_3), .B(n_225), .Y(n_602) );
OAI211xp5_ASAP7_75t_SL g1363 ( .A1(n_4), .A2(n_1196), .B(n_1274), .C(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1375 ( .A(n_4), .Y(n_1375) );
INVx1_ASAP7_75t_L g782 ( .A(n_5), .Y(n_782) );
INVx1_ASAP7_75t_L g1384 ( .A(n_6), .Y(n_1384) );
OAI22xp5_ASAP7_75t_L g1185 ( .A1(n_7), .A2(n_135), .B1(n_1060), .B2(n_1186), .Y(n_1185) );
OAI22xp5_ASAP7_75t_L g1202 ( .A1(n_7), .A2(n_135), .B1(n_861), .B2(n_1044), .Y(n_1202) );
AOI22xp5_ASAP7_75t_L g1460 ( .A1(n_8), .A2(n_51), .B1(n_1435), .B2(n_1441), .Y(n_1460) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_9), .A2(n_248), .B1(n_328), .B2(n_1058), .Y(n_1190) );
OAI22xp33_ASAP7_75t_L g1198 ( .A1(n_9), .A2(n_248), .B1(n_1053), .B2(n_1109), .Y(n_1198) );
OAI211xp5_ASAP7_75t_L g780 ( .A1(n_10), .A2(n_411), .B(n_668), .C(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g795 ( .A(n_10), .Y(n_795) );
INVx1_ASAP7_75t_L g1005 ( .A(n_11), .Y(n_1005) );
INVx1_ASAP7_75t_L g519 ( .A(n_12), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_13), .A2(n_164), .B1(n_687), .B2(n_689), .Y(n_686) );
INVx1_ASAP7_75t_L g702 ( .A(n_13), .Y(n_702) );
INVx1_ASAP7_75t_L g1408 ( .A(n_14), .Y(n_1408) );
OAI211xp5_ASAP7_75t_L g1417 ( .A1(n_14), .A2(n_453), .B(n_1418), .C(n_1419), .Y(n_1417) );
OAI22xp33_ASAP7_75t_L g1107 ( .A1(n_15), .A2(n_154), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
OAI22xp33_ASAP7_75t_L g1111 ( .A1(n_15), .A2(n_154), .B1(n_328), .B2(n_788), .Y(n_1111) );
INVx1_ASAP7_75t_L g1387 ( .A(n_16), .Y(n_1387) );
CKINVDCx5p33_ASAP7_75t_R g1301 ( .A(n_17), .Y(n_1301) );
INVx2_ASAP7_75t_L g402 ( .A(n_18), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_19), .A2(n_311), .B1(n_609), .B2(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g624 ( .A(n_19), .Y(n_624) );
INVx1_ASAP7_75t_L g1152 ( .A(n_20), .Y(n_1152) );
INVx1_ASAP7_75t_L g1347 ( .A(n_21), .Y(n_1347) );
INVx1_ASAP7_75t_L g1021 ( .A(n_22), .Y(n_1021) );
AOI22xp5_ASAP7_75t_L g1474 ( .A1(n_23), .A2(n_201), .B1(n_1431), .B2(n_1438), .Y(n_1474) );
INVx1_ASAP7_75t_L g1393 ( .A(n_24), .Y(n_1393) );
OA222x2_ASAP7_75t_L g929 ( .A1(n_25), .A2(n_66), .B1(n_220), .B2(n_930), .C1(n_933), .C2(n_937), .Y(n_929) );
INVx1_ASAP7_75t_L g981 ( .A(n_25), .Y(n_981) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_26), .Y(n_321) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_26), .B(n_319), .Y(n_1432) );
AOI22xp5_ASAP7_75t_L g1459 ( .A1(n_27), .A2(n_185), .B1(n_1431), .B2(n_1438), .Y(n_1459) );
INVx1_ASAP7_75t_L g1271 ( .A(n_28), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_29), .A2(n_289), .B1(n_708), .B2(n_709), .Y(n_820) );
INVxp67_ASAP7_75t_SL g839 ( .A(n_29), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_30), .A2(n_191), .B1(n_585), .B2(n_587), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_30), .A2(n_237), .B1(n_640), .B2(n_642), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g1465 ( .A1(n_31), .A2(n_249), .B1(n_1431), .B2(n_1438), .Y(n_1465) );
INVx1_ASAP7_75t_L g545 ( .A(n_32), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g1305 ( .A(n_33), .Y(n_1305) );
INVx1_ASAP7_75t_L g1704 ( .A(n_34), .Y(n_1704) );
AOI22xp5_ASAP7_75t_L g1454 ( .A1(n_35), .A2(n_99), .B1(n_1431), .B2(n_1438), .Y(n_1454) );
INVx1_ASAP7_75t_L g739 ( .A(n_36), .Y(n_739) );
INVx1_ASAP7_75t_L g1015 ( .A(n_37), .Y(n_1015) );
INVx1_ASAP7_75t_L g1711 ( .A(n_38), .Y(n_1711) );
INVx1_ASAP7_75t_L g1083 ( .A(n_39), .Y(n_1083) );
CKINVDCx5p33_ASAP7_75t_R g950 ( .A(n_40), .Y(n_950) );
INVx1_ASAP7_75t_L g673 ( .A(n_41), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g711 ( .A1(n_41), .A2(n_712), .B(n_713), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g1452 ( .A1(n_42), .A2(n_166), .B1(n_1441), .B2(n_1453), .Y(n_1452) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_43), .A2(n_232), .B1(n_708), .B2(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_43), .A2(n_216), .B1(n_841), .B2(n_842), .Y(n_840) );
INVx1_ASAP7_75t_L g1103 ( .A(n_44), .Y(n_1103) );
OAI22xp33_ASAP7_75t_L g784 ( .A1(n_45), .A2(n_127), .B1(n_469), .B2(n_785), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_45), .A2(n_127), .B1(n_505), .B2(n_797), .Y(n_796) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_46), .Y(n_333) );
INVx1_ASAP7_75t_L g1079 ( .A(n_47), .Y(n_1079) );
OAI22xp33_ASAP7_75t_SL g813 ( .A1(n_48), .A2(n_223), .B1(n_814), .B2(n_815), .Y(n_813) );
INVx1_ASAP7_75t_L g856 ( .A(n_48), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_49), .A2(n_89), .B1(n_613), .B2(n_952), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_49), .A2(n_208), .B1(n_431), .B2(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g664 ( .A(n_50), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_50), .A2(n_277), .B1(n_695), .B2(n_697), .Y(n_694) );
XNOR2xp5_ASAP7_75t_L g1000 ( .A(n_51), .B(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1275 ( .A(n_52), .Y(n_1275) );
INVx1_ASAP7_75t_L g1208 ( .A(n_53), .Y(n_1208) );
AOI21xp33_ASAP7_75t_L g892 ( .A1(n_54), .A2(n_582), .B(n_893), .Y(n_892) );
AOI221xp5_ASAP7_75t_L g912 ( .A1(n_54), .A2(n_239), .B1(n_907), .B2(n_913), .C(n_916), .Y(n_912) );
XOR2x2_ASAP7_75t_L g1122 ( .A(n_55), .B(n_1123), .Y(n_1122) );
OAI222xp33_ASAP7_75t_L g870 ( .A1(n_56), .A2(n_64), .B1(n_70), .B2(n_521), .C1(n_871), .C2(n_872), .Y(n_870) );
OAI22xp33_ASAP7_75t_L g1315 ( .A1(n_57), .A2(n_104), .B1(n_328), .B2(n_788), .Y(n_1315) );
OAI22xp33_ASAP7_75t_L g1325 ( .A1(n_57), .A2(n_104), .B1(n_449), .B2(n_1053), .Y(n_1325) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_58), .A2(n_606), .B(n_607), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_58), .A2(n_191), .B1(n_626), .B2(n_629), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_59), .A2(n_214), .B1(n_1435), .B2(n_1441), .Y(n_1532) );
INVx1_ASAP7_75t_L g1051 ( .A(n_60), .Y(n_1051) );
OAI211xp5_ASAP7_75t_L g1065 ( .A1(n_60), .A2(n_790), .B(n_1066), .C(n_1067), .Y(n_1065) );
OAI22xp33_ASAP7_75t_L g1698 ( .A1(n_61), .A2(n_65), .B1(n_1699), .B2(n_1700), .Y(n_1698) );
OAI22xp33_ASAP7_75t_L g1735 ( .A1(n_61), .A2(n_65), .B1(n_1044), .B2(n_1416), .Y(n_1735) );
CKINVDCx5p33_ASAP7_75t_R g877 ( .A(n_62), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_63), .Y(n_572) );
OAI221xp5_ASAP7_75t_L g966 ( .A1(n_66), .A2(n_181), .B1(n_967), .B2(n_969), .C(n_971), .Y(n_966) );
INVx1_ASAP7_75t_L g944 ( .A(n_67), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_67), .A2(n_123), .B1(n_638), .B2(n_640), .Y(n_998) );
INVx1_ASAP7_75t_L g1720 ( .A(n_68), .Y(n_1720) );
XOR2x2_ASAP7_75t_L g1243 ( .A(n_69), .B(n_1244), .Y(n_1243) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_70), .A2(n_307), .B1(n_697), .B2(n_901), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g1437 ( .A1(n_71), .A2(n_167), .B1(n_1438), .B2(n_1441), .Y(n_1437) );
INVx1_ASAP7_75t_L g1340 ( .A(n_72), .Y(n_1340) );
INVx1_ASAP7_75t_L g1365 ( .A(n_73), .Y(n_1365) );
INVx1_ASAP7_75t_L g1248 ( .A(n_74), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_75), .A2(n_273), .B1(n_1431), .B2(n_1435), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_76), .A2(n_150), .B1(n_587), .B2(n_609), .Y(n_894) );
INVx1_ASAP7_75t_L g909 ( .A(n_76), .Y(n_909) );
INVx1_ASAP7_75t_L g1013 ( .A(n_77), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1655 ( .A1(n_78), .A2(n_244), .B1(n_846), .B2(n_855), .Y(n_1655) );
AOI221xp5_ASAP7_75t_L g1660 ( .A1(n_78), .A2(n_241), .B1(n_580), .B2(n_893), .C(n_1661), .Y(n_1660) );
AOI22xp5_ASAP7_75t_L g1477 ( .A1(n_79), .A2(n_148), .B1(n_1441), .B2(n_1450), .Y(n_1477) );
INVx1_ASAP7_75t_L g1650 ( .A(n_80), .Y(n_1650) );
AOI22xp33_ASAP7_75t_L g1662 ( .A1(n_80), .A2(n_269), .B1(n_587), .B2(n_1663), .Y(n_1662) );
XNOR2xp5_ASAP7_75t_L g734 ( .A(n_81), .B(n_735), .Y(n_734) );
OAI211xp5_ASAP7_75t_L g1191 ( .A1(n_82), .A2(n_890), .B(n_1192), .C(n_1196), .Y(n_1191) );
INVx1_ASAP7_75t_L g1201 ( .A(n_82), .Y(n_1201) );
INVx1_ASAP7_75t_L g746 ( .A(n_83), .Y(n_746) );
INVx1_ASAP7_75t_L g1080 ( .A(n_84), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1533 ( .A1(n_85), .A2(n_296), .B1(n_1431), .B2(n_1438), .Y(n_1533) );
OAI22xp33_ASAP7_75t_L g447 ( .A1(n_86), .A2(n_145), .B1(n_448), .B2(n_449), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g478 ( .A1(n_86), .A2(n_145), .B1(n_328), .B2(n_479), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g1696 ( .A1(n_87), .A2(n_136), .B1(n_1058), .B2(n_1697), .Y(n_1696) );
OAI22xp5_ASAP7_75t_L g1731 ( .A1(n_87), .A2(n_136), .B1(n_1372), .B2(n_1413), .Y(n_1731) );
OAI22xp33_ASAP7_75t_L g1403 ( .A1(n_88), .A2(n_96), .B1(n_788), .B2(n_1252), .Y(n_1403) );
OAI22xp33_ASAP7_75t_L g1412 ( .A1(n_88), .A2(n_96), .B1(n_1054), .B2(n_1413), .Y(n_1412) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_89), .A2(n_110), .B1(n_741), .B2(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g356 ( .A(n_90), .Y(n_356) );
INVx1_ASAP7_75t_L g685 ( .A(n_91), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_91), .A2(n_227), .B1(n_708), .B2(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g1641 ( .A(n_92), .Y(n_1641) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_93), .Y(n_568) );
INVx1_ASAP7_75t_L g319 ( .A(n_94), .Y(n_319) );
INVx1_ASAP7_75t_L g1011 ( .A(n_95), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_97), .A2(n_161), .B1(n_521), .B2(n_1154), .Y(n_1153) );
OAI211xp5_ASAP7_75t_L g1246 ( .A1(n_98), .A2(n_833), .B(n_1196), .C(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1259 ( .A(n_98), .Y(n_1259) );
INVx1_ASAP7_75t_L g1195 ( .A(n_100), .Y(n_1195) );
OAI211xp5_ASAP7_75t_L g1199 ( .A1(n_100), .A2(n_443), .B(n_668), .C(n_1200), .Y(n_1199) );
INVxp67_ASAP7_75t_SL g1144 ( .A(n_101), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_101), .A2(n_250), .B1(n_677), .B2(n_1170), .Y(n_1169) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_102), .A2(n_141), .B1(n_810), .B2(n_811), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_102), .B(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g1353 ( .A(n_103), .Y(n_1353) );
INVx1_ASAP7_75t_L g385 ( .A(n_105), .Y(n_385) );
INVx1_ASAP7_75t_L g1349 ( .A(n_106), .Y(n_1349) );
INVx1_ASAP7_75t_L g1351 ( .A(n_107), .Y(n_1351) );
OAI22xp5_ASAP7_75t_L g1368 ( .A1(n_108), .A2(n_120), .B1(n_506), .B2(n_1188), .Y(n_1368) );
OAI22xp33_ASAP7_75t_L g1376 ( .A1(n_108), .A2(n_120), .B1(n_1106), .B2(n_1255), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g1653 ( .A(n_109), .Y(n_1653) );
AOI221xp5_ASAP7_75t_L g1145 ( .A1(n_110), .A2(n_208), .B1(n_712), .B2(n_713), .C(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1280 ( .A(n_111), .Y(n_1280) );
OAI22xp5_ASAP7_75t_L g1409 ( .A1(n_112), .A2(n_267), .B1(n_505), .B2(n_1188), .Y(n_1409) );
OAI22xp5_ASAP7_75t_L g1415 ( .A1(n_112), .A2(n_267), .B1(n_469), .B2(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1407 ( .A(n_113), .Y(n_1407) );
INVx1_ASAP7_75t_L g1367 ( .A(n_114), .Y(n_1367) );
OAI211xp5_ASAP7_75t_L g1373 ( .A1(n_114), .A2(n_453), .B(n_1257), .C(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1341 ( .A(n_115), .Y(n_1341) );
INVx1_ASAP7_75t_L g1378 ( .A(n_116), .Y(n_1378) );
AOI22xp33_ASAP7_75t_SL g1464 ( .A1(n_116), .A2(n_196), .B1(n_1435), .B2(n_1441), .Y(n_1464) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_117), .A2(n_251), .B1(n_676), .B2(n_678), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_117), .A2(n_607), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g1649 ( .A(n_118), .Y(n_1649) );
AOI21xp33_ASAP7_75t_L g1671 ( .A1(n_118), .A2(n_893), .B(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1082 ( .A(n_119), .Y(n_1082) );
OAI211xp5_ASAP7_75t_L g1099 ( .A1(n_121), .A2(n_668), .B(n_1100), .C(n_1102), .Y(n_1099) );
INVx1_ASAP7_75t_L g1115 ( .A(n_121), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g1642 ( .A1(n_122), .A2(n_163), .B1(n_1643), .B2(n_1644), .Y(n_1642) );
OAI211xp5_ASAP7_75t_L g1658 ( .A1(n_122), .A2(n_1126), .B(n_1659), .C(n_1665), .Y(n_1658) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_123), .A2(n_168), .B1(n_613), .B2(n_952), .Y(n_951) );
AOI221xp5_ASAP7_75t_L g1129 ( .A1(n_124), .A2(n_250), .B1(n_1130), .B2(n_1131), .C(n_1132), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_124), .A2(n_211), .B1(n_1159), .B2(n_1161), .Y(n_1158) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_125), .A2(n_295), .B1(n_505), .B2(n_507), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1254 ( .A1(n_125), .A2(n_295), .B1(n_861), .B2(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1090 ( .A(n_126), .Y(n_1090) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_128), .A2(n_181), .B1(n_958), .B2(n_961), .Y(n_957) );
INVx1_ASAP7_75t_L g982 ( .A(n_128), .Y(n_982) );
INVx1_ASAP7_75t_L g363 ( .A(n_129), .Y(n_363) );
INVx1_ASAP7_75t_L g369 ( .A(n_130), .Y(n_369) );
OAI211xp5_ASAP7_75t_L g1316 ( .A1(n_131), .A2(n_1196), .B(n_1317), .C(n_1319), .Y(n_1316) );
INVx1_ASAP7_75t_L g1330 ( .A(n_131), .Y(n_1330) );
OAI22xp33_ASAP7_75t_L g1251 ( .A1(n_132), .A2(n_171), .B1(n_788), .B2(n_1252), .Y(n_1251) );
OAI22xp33_ASAP7_75t_L g1260 ( .A1(n_132), .A2(n_171), .B1(n_448), .B2(n_1054), .Y(n_1260) );
OAI22xp33_ASAP7_75t_L g1369 ( .A1(n_133), .A2(n_217), .B1(n_479), .B2(n_1252), .Y(n_1369) );
OAI22xp33_ASAP7_75t_L g1371 ( .A1(n_133), .A2(n_217), .B1(n_448), .B2(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1714 ( .A(n_134), .Y(n_1714) );
OAI221xp5_ASAP7_75t_L g830 ( .A1(n_137), .A2(n_291), .B1(n_831), .B2(n_832), .C(n_833), .Y(n_830) );
INVx1_ASAP7_75t_L g851 ( .A(n_137), .Y(n_851) );
INVx1_ASAP7_75t_L g818 ( .A(n_138), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_138), .A2(n_232), .B1(n_841), .B2(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g761 ( .A(n_139), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_140), .Y(n_822) );
INVx1_ASAP7_75t_L g854 ( .A(n_141), .Y(n_854) );
INVx1_ASAP7_75t_L g753 ( .A(n_142), .Y(n_753) );
OAI22xp33_ASAP7_75t_L g1052 ( .A1(n_143), .A2(n_228), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_143), .A2(n_228), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
INVx1_ASAP7_75t_L g1390 ( .A(n_144), .Y(n_1390) );
INVx1_ASAP7_75t_L g1193 ( .A(n_146), .Y(n_1193) );
INVx1_ASAP7_75t_L g1008 ( .A(n_147), .Y(n_1008) );
INVx1_ASAP7_75t_L g1017 ( .A(n_149), .Y(n_1017) );
INVxp67_ASAP7_75t_SL g917 ( .A(n_150), .Y(n_917) );
XOR2xp5_ASAP7_75t_L g1686 ( .A(n_151), .B(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g462 ( .A(n_152), .Y(n_462) );
INVx1_ASAP7_75t_L g1087 ( .A(n_153), .Y(n_1087) );
INVx1_ASAP7_75t_L g755 ( .A(n_155), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g777 ( .A1(n_156), .A2(n_300), .B1(n_449), .B2(n_778), .Y(n_777) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_156), .A2(n_300), .B1(n_328), .B2(n_788), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_157), .A2(n_179), .B1(n_785), .B2(n_1044), .Y(n_1043) );
OAI22xp33_ASAP7_75t_L g1059 ( .A1(n_157), .A2(n_179), .B1(n_1060), .B2(n_1062), .Y(n_1059) );
OAI211xp5_ASAP7_75t_L g1404 ( .A1(n_158), .A2(n_1217), .B(n_1405), .C(n_1406), .Y(n_1404) );
INVx1_ASAP7_75t_L g1420 ( .A(n_158), .Y(n_1420) );
INVx1_ASAP7_75t_L g744 ( .A(n_159), .Y(n_744) );
INVx1_ASAP7_75t_L g376 ( .A(n_160), .Y(n_376) );
OAI211xp5_ASAP7_75t_L g1125 ( .A1(n_161), .A2(n_1126), .B(n_1128), .C(n_1134), .Y(n_1125) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_162), .A2(n_298), .B1(n_578), .B2(n_580), .C(n_582), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_162), .A2(n_311), .B1(n_636), .B2(n_637), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_164), .A2(n_251), .B1(n_708), .B2(n_709), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g949 ( .A(n_165), .Y(n_949) );
INVx1_ASAP7_75t_L g803 ( .A(n_166), .Y(n_803) );
INVx1_ASAP7_75t_L g994 ( .A(n_168), .Y(n_994) );
INVx1_ASAP7_75t_L g1273 ( .A(n_169), .Y(n_1273) );
INVx1_ASAP7_75t_L g1249 ( .A(n_170), .Y(n_1249) );
OAI211xp5_ASAP7_75t_L g1256 ( .A1(n_170), .A2(n_453), .B(n_1257), .C(n_1258), .Y(n_1256) );
OAI22xp33_ASAP7_75t_L g1105 ( .A1(n_172), .A2(n_301), .B1(n_1044), .B2(n_1106), .Y(n_1105) );
OAI22xp33_ASAP7_75t_L g1112 ( .A1(n_172), .A2(n_301), .B1(n_1060), .B2(n_1062), .Y(n_1112) );
INVx1_ASAP7_75t_L g891 ( .A(n_173), .Y(n_891) );
AOI221x1_ASAP7_75t_SL g906 ( .A1(n_173), .A2(n_234), .B1(n_741), .B2(n_907), .C(n_908), .Y(n_906) );
INVx1_ASAP7_75t_L g1383 ( .A(n_174), .Y(n_1383) );
AOI221x1_ASAP7_75t_SL g939 ( .A1(n_175), .A2(n_230), .B1(n_940), .B2(n_942), .C(n_943), .Y(n_939) );
AOI21xp33_ASAP7_75t_L g996 ( .A1(n_175), .A2(n_915), .B(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g1135 ( .A(n_176), .Y(n_1135) );
OAI22xp33_ASAP7_75t_L g1175 ( .A1(n_176), .A2(n_275), .B1(n_1176), .B2(n_1177), .Y(n_1175) );
AOI21xp33_ASAP7_75t_L g898 ( .A1(n_177), .A2(n_606), .B(n_607), .Y(n_898) );
INVx1_ASAP7_75t_L g919 ( .A(n_177), .Y(n_919) );
OAI221xp5_ASAP7_75t_L g1138 ( .A1(n_178), .A2(n_231), .B1(n_1139), .B2(n_1140), .C(n_1141), .Y(n_1138) );
INVx1_ASAP7_75t_L g1172 ( .A(n_178), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_180), .B(n_1434), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_180), .B(n_270), .Y(n_1436) );
INVx2_ASAP7_75t_L g1440 ( .A(n_180), .Y(n_1440) );
INVx1_ASAP7_75t_L g1667 ( .A(n_182), .Y(n_1667) );
INVx1_ASAP7_75t_L g1694 ( .A(n_183), .Y(n_1694) );
AOI22xp5_ASAP7_75t_L g1448 ( .A1(n_184), .A2(n_224), .B1(n_1431), .B2(n_1441), .Y(n_1448) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_186), .A2(n_517), .B1(n_645), .B2(n_646), .Y(n_516) );
INVxp67_ASAP7_75t_L g646 ( .A(n_186), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g945 ( .A(n_187), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1449 ( .A1(n_188), .A2(n_192), .B1(n_1438), .B2(n_1450), .Y(n_1449) );
AOI22xp33_ASAP7_75t_SL g1651 ( .A1(n_189), .A2(n_241), .B1(n_846), .B2(n_855), .Y(n_1651) );
AOI22xp33_ASAP7_75t_SL g1673 ( .A1(n_189), .A2(n_244), .B1(n_591), .B2(n_826), .Y(n_1673) );
OAI211xp5_ASAP7_75t_L g1692 ( .A1(n_190), .A2(n_1066), .B(n_1094), .C(n_1693), .Y(n_1692) );
INVx1_ASAP7_75t_L g1734 ( .A(n_190), .Y(n_1734) );
XOR2x2_ASAP7_75t_L g1181 ( .A(n_192), .B(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g465 ( .A(n_193), .Y(n_465) );
OAI211xp5_ASAP7_75t_L g485 ( .A1(n_193), .A2(n_486), .B(n_488), .C(n_494), .Y(n_485) );
XOR2x2_ASAP7_75t_L g1289 ( .A(n_194), .B(n_1290), .Y(n_1289) );
OAI221xp5_ASAP7_75t_SL g554 ( .A1(n_195), .A2(n_265), .B1(n_555), .B2(n_561), .C(n_567), .Y(n_554) );
INVx1_ASAP7_75t_L g597 ( .A(n_195), .Y(n_597) );
INVx2_ASAP7_75t_L g401 ( .A(n_197), .Y(n_401) );
INVx1_ASAP7_75t_L g441 ( .A(n_197), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_197), .B(n_402), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g1478 ( .A1(n_198), .A2(n_304), .B1(n_1431), .B2(n_1438), .Y(n_1478) );
INVx1_ASAP7_75t_L g748 ( .A(n_199), .Y(n_748) );
INVx1_ASAP7_75t_L g1394 ( .A(n_200), .Y(n_1394) );
OAI22xp5_ASAP7_75t_L g1322 ( .A1(n_202), .A2(n_206), .B1(n_797), .B2(n_1323), .Y(n_1322) );
OAI22xp33_ASAP7_75t_L g1331 ( .A1(n_202), .A2(n_206), .B1(n_1106), .B2(n_1332), .Y(n_1331) );
CKINVDCx5p33_ASAP7_75t_R g1299 ( .A(n_203), .Y(n_1299) );
INVx1_ASAP7_75t_L g868 ( .A(n_204), .Y(n_868) );
INVx1_ASAP7_75t_L g1388 ( .A(n_205), .Y(n_1388) );
BUFx3_ASAP7_75t_L g408 ( .A(n_207), .Y(n_408) );
INVx1_ASAP7_75t_L g529 ( .A(n_209), .Y(n_529) );
INVx1_ASAP7_75t_L g1104 ( .A(n_210), .Y(n_1104) );
OAI211xp5_ASAP7_75t_L g1113 ( .A1(n_210), .A2(n_790), .B(n_1066), .C(n_1114), .Y(n_1113) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_211), .Y(n_1142) );
OAI22xp5_ASAP7_75t_SL g880 ( .A1(n_212), .A2(n_252), .B1(n_570), .B2(n_574), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g888 ( .A(n_212), .Y(n_888) );
INVx1_ASAP7_75t_L g1267 ( .A(n_213), .Y(n_1267) );
CKINVDCx5p33_ASAP7_75t_R g1295 ( .A(n_215), .Y(n_1295) );
AOI21xp33_ASAP7_75t_L g819 ( .A1(n_216), .A2(n_606), .B(n_607), .Y(n_819) );
INVx1_ASAP7_75t_L g1211 ( .A(n_218), .Y(n_1211) );
INVx1_ASAP7_75t_L g1710 ( .A(n_219), .Y(n_1710) );
INVx1_ASAP7_75t_L g972 ( .A(n_220), .Y(n_972) );
INVx1_ASAP7_75t_L g659 ( .A(n_221), .Y(n_659) );
INVx1_ASAP7_75t_L g1020 ( .A(n_222), .Y(n_1020) );
INVx1_ASAP7_75t_L g859 ( .A(n_223), .Y(n_859) );
BUFx3_ASAP7_75t_L g336 ( .A(n_225), .Y(n_336) );
INVx1_ASAP7_75t_L g482 ( .A(n_225), .Y(n_482) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_226), .A2(n_274), .B1(n_467), .B2(n_469), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_226), .A2(n_274), .B1(n_505), .B2(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g674 ( .A(n_227), .Y(n_674) );
XNOR2xp5_ASAP7_75t_L g1335 ( .A(n_229), .B(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g993 ( .A(n_230), .Y(n_993) );
INVx1_ASAP7_75t_L g1174 ( .A(n_231), .Y(n_1174) );
INVx1_ASAP7_75t_L g927 ( .A(n_233), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_234), .A2(n_239), .B1(n_587), .B2(n_609), .Y(n_899) );
INVx1_ASAP7_75t_L g1345 ( .A(n_235), .Y(n_1345) );
INVx1_ASAP7_75t_L g1221 ( .A(n_236), .Y(n_1221) );
INVx1_ASAP7_75t_L g604 ( .A(n_237), .Y(n_604) );
INVx1_ASAP7_75t_L g1695 ( .A(n_238), .Y(n_1695) );
OAI211xp5_ASAP7_75t_L g1732 ( .A1(n_238), .A2(n_668), .B(n_749), .C(n_1733), .Y(n_1732) );
INVx1_ASAP7_75t_L g1269 ( .A(n_240), .Y(n_1269) );
INVx1_ASAP7_75t_L g1666 ( .A(n_242), .Y(n_1666) );
CKINVDCx5p33_ASAP7_75t_R g1302 ( .A(n_243), .Y(n_1302) );
INVx1_ASAP7_75t_L g1715 ( .A(n_245), .Y(n_1715) );
INVx1_ASAP7_75t_L g1220 ( .A(n_246), .Y(n_1220) );
INVx1_ASAP7_75t_L g380 ( .A(n_247), .Y(n_380) );
INVx1_ASAP7_75t_L g884 ( .A(n_252), .Y(n_884) );
INVx1_ASAP7_75t_L g1216 ( .A(n_253), .Y(n_1216) );
INVx1_ASAP7_75t_L g410 ( .A(n_254), .Y(n_410) );
INVx1_ASAP7_75t_L g416 ( .A(n_254), .Y(n_416) );
INVx1_ASAP7_75t_L g783 ( .A(n_255), .Y(n_783) );
OAI211xp5_ASAP7_75t_L g789 ( .A1(n_255), .A2(n_790), .B(n_792), .C(n_794), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_256), .A2(n_648), .B1(n_649), .B2(n_729), .Y(n_647) );
INVxp67_ASAP7_75t_L g729 ( .A(n_256), .Y(n_729) );
INVx1_ASAP7_75t_L g1085 ( .A(n_257), .Y(n_1085) );
INVx1_ASAP7_75t_L g1227 ( .A(n_258), .Y(n_1227) );
CKINVDCx5p33_ASAP7_75t_R g1320 ( .A(n_259), .Y(n_1320) );
INVxp67_ASAP7_75t_SL g653 ( .A(n_260), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_260), .A2(n_299), .B1(n_717), .B2(n_718), .C(n_721), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g1297 ( .A(n_261), .Y(n_1297) );
INVx1_ASAP7_75t_L g386 ( .A(n_262), .Y(n_386) );
INVx1_ASAP7_75t_L g896 ( .A(n_263), .Y(n_896) );
INVx1_ASAP7_75t_L g1050 ( .A(n_264), .Y(n_1050) );
INVx1_ASAP7_75t_L g615 ( .A(n_265), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_266), .Y(n_661) );
AOI22xp5_ASAP7_75t_SL g1473 ( .A1(n_268), .A2(n_309), .B1(n_1441), .B2(n_1450), .Y(n_1473) );
INVx1_ASAP7_75t_L g1654 ( .A(n_269), .Y(n_1654) );
INVx1_ASAP7_75t_L g1434 ( .A(n_270), .Y(n_1434) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_270), .B(n_1440), .Y(n_1442) );
OAI211xp5_ASAP7_75t_SL g1045 ( .A1(n_271), .A2(n_668), .B(n_1046), .C(n_1048), .Y(n_1045) );
INVx1_ASAP7_75t_L g1072 ( .A(n_271), .Y(n_1072) );
CKINVDCx5p33_ASAP7_75t_R g1304 ( .A(n_272), .Y(n_1304) );
INVx1_ASAP7_75t_L g1136 ( .A(n_275), .Y(n_1136) );
INVx1_ASAP7_75t_L g1265 ( .A(n_276), .Y(n_1265) );
INVx1_ASAP7_75t_L g666 ( .A(n_277), .Y(n_666) );
INVx1_ASAP7_75t_L g828 ( .A(n_278), .Y(n_828) );
INVx1_ASAP7_75t_L g1321 ( .A(n_279), .Y(n_1321) );
OAI211xp5_ASAP7_75t_L g1326 ( .A1(n_279), .A2(n_453), .B(n_1327), .C(n_1329), .Y(n_1326) );
INVx1_ASAP7_75t_L g759 ( .A(n_280), .Y(n_759) );
CKINVDCx5p33_ASAP7_75t_R g683 ( .A(n_281), .Y(n_683) );
INVx1_ASAP7_75t_L g1226 ( .A(n_282), .Y(n_1226) );
INVx1_ASAP7_75t_L g1391 ( .A(n_283), .Y(n_1391) );
AOI21xp5_ASAP7_75t_SL g823 ( .A1(n_284), .A2(n_606), .B(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g838 ( .A(n_284), .Y(n_838) );
XNOR2xp5_ASAP7_75t_L g1074 ( .A(n_285), .B(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1089 ( .A(n_286), .Y(n_1089) );
INVx1_ASAP7_75t_L g353 ( .A(n_287), .Y(n_353) );
XOR2x2_ASAP7_75t_L g342 ( .A(n_288), .B(n_343), .Y(n_342) );
INVxp67_ASAP7_75t_L g844 ( .A(n_289), .Y(n_844) );
CKINVDCx5p33_ASAP7_75t_R g1294 ( .A(n_290), .Y(n_1294) );
INVxp67_ASAP7_75t_SL g858 ( .A(n_291), .Y(n_858) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_292), .Y(n_332) );
INVx1_ASAP7_75t_L g1706 ( .A(n_293), .Y(n_1706) );
INVx1_ASAP7_75t_L g1721 ( .A(n_294), .Y(n_1721) );
CKINVDCx5p33_ASAP7_75t_R g963 ( .A(n_297), .Y(n_963) );
INVx1_ASAP7_75t_L g623 ( .A(n_298), .Y(n_623) );
INVx1_ASAP7_75t_L g656 ( .A(n_299), .Y(n_656) );
INVx1_ASAP7_75t_L g1279 ( .A(n_302), .Y(n_1279) );
INVx1_ASAP7_75t_L g1218 ( .A(n_303), .Y(n_1218) );
INVx2_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
INVx1_ASAP7_75t_L g396 ( .A(n_305), .Y(n_396) );
INVx1_ASAP7_75t_L g440 ( .A(n_305), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g964 ( .A(n_306), .Y(n_964) );
INVx1_ASAP7_75t_L g879 ( .A(n_307), .Y(n_879) );
OAI22xp33_ASAP7_75t_SL g1656 ( .A1(n_308), .A2(n_310), .B1(n_561), .B2(n_876), .Y(n_1656) );
OAI221xp5_ASAP7_75t_L g1668 ( .A1(n_308), .A2(n_310), .B1(n_718), .B2(n_1669), .C(n_1670), .Y(n_1668) );
XNOR2xp5_ASAP7_75t_L g1638 ( .A(n_309), .B(n_1639), .Y(n_1638) );
AOI22xp33_ASAP7_75t_L g1682 ( .A1(n_309), .A2(n_1683), .B1(n_1685), .B2(n_1737), .Y(n_1682) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_337), .B(n_1424), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_322), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g1681 ( .A(n_316), .B(n_325), .Y(n_1681) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g1684 ( .A(n_318), .B(n_321), .Y(n_1684) );
INVx1_ASAP7_75t_L g1738 ( .A(n_318), .Y(n_1738) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g1740 ( .A(n_321), .B(n_1738), .Y(n_1740) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g511 ( .A(n_325), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g391 ( .A(n_326), .B(n_336), .Y(n_391) );
AND2x4_ASAP7_75t_L g583 ( .A(n_326), .B(n_335), .Y(n_583) );
INVxp67_ASAP7_75t_SL g1057 ( .A(n_327), .Y(n_1057) );
AND2x4_ASAP7_75t_SL g1680 ( .A(n_327), .B(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1697 ( .A(n_327), .Y(n_1697) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x6_ASAP7_75t_L g328 ( .A(n_329), .B(n_334), .Y(n_328) );
INVxp67_ASAP7_75t_L g355 ( .A(n_329), .Y(n_355) );
OR2x6_ASAP7_75t_L g506 ( .A(n_329), .B(n_481), .Y(n_506) );
BUFx4f_ASAP7_75t_L g764 ( .A(n_329), .Y(n_764) );
INVx1_ASAP7_75t_L g1039 ( .A(n_329), .Y(n_1039) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx3_ASAP7_75t_L g384 ( .A(n_330), .Y(n_384) );
BUFx4f_ASAP7_75t_L g1027 ( .A(n_330), .Y(n_1027) );
INVx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx2_ASAP7_75t_L g361 ( .A(n_332), .Y(n_361) );
INVx2_ASAP7_75t_L g368 ( .A(n_332), .Y(n_368) );
NAND2x1_ASAP7_75t_L g372 ( .A(n_332), .B(n_333), .Y(n_372) );
AND2x2_ASAP7_75t_L g483 ( .A(n_332), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g493 ( .A(n_332), .B(n_333), .Y(n_493) );
INVx1_ASAP7_75t_L g502 ( .A(n_332), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_333), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g367 ( .A(n_333), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g484 ( .A(n_333), .Y(n_484) );
BUFx2_ASAP7_75t_L g497 ( .A(n_333), .Y(n_497) );
INVx1_ASAP7_75t_L g537 ( .A(n_333), .Y(n_537) );
AND2x2_ASAP7_75t_L g588 ( .A(n_333), .B(n_361), .Y(n_588) );
OR2x6_ASAP7_75t_L g1252 ( .A(n_334), .B(n_384), .Y(n_1252) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g490 ( .A(n_335), .Y(n_490) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g496 ( .A(n_336), .Y(n_496) );
AND2x4_ASAP7_75t_L g500 ( .A(n_336), .B(n_501), .Y(n_500) );
XNOR2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_798), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AO22x2_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_731), .B2(n_732), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AO22x2_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_514), .B1(n_515), .B2(n_730), .Y(n_341) );
INVx1_ASAP7_75t_L g730 ( .A(n_342), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_446), .C(n_477), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_397), .Y(n_344) );
OAI33xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_352), .A3(n_362), .B1(n_373), .B2(n_381), .B3(n_389), .Y(n_345) );
OAI33xp33_ASAP7_75t_L g1306 ( .A1(n_346), .A2(n_389), .A3(n_1307), .B1(n_1308), .B2(n_1309), .B3(n_1312), .Y(n_1306) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g766 ( .A(n_348), .Y(n_766) );
INVx1_ASAP7_75t_L g1023 ( .A(n_348), .Y(n_1023) );
INVx2_ASAP7_75t_L g1206 ( .A(n_348), .Y(n_1206) );
INVx4_ASAP7_75t_L g1357 ( .A(n_348), .Y(n_1357) );
INVx2_ASAP7_75t_L g1398 ( .A(n_348), .Y(n_1398) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g619 ( .A(n_349), .Y(n_619) );
OR2x6_ASAP7_75t_L g1168 ( .A(n_349), .B(n_990), .Y(n_1168) );
BUFx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g728 ( .A(n_350), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_350), .B(n_602), .Y(n_956) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_356), .B2(n_357), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_353), .A2(n_376), .B1(n_404), .B2(n_411), .Y(n_403) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g442 ( .A1(n_356), .A2(n_380), .B1(n_404), .B2(n_443), .Y(n_442) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
INVx1_ASAP7_75t_L g765 ( .A(n_358), .Y(n_765) );
INVx2_ASAP7_75t_L g812 ( .A(n_358), .Y(n_812) );
INVx1_ASAP7_75t_L g1041 ( .A(n_358), .Y(n_1041) );
INVx4_ASAP7_75t_L g1214 ( .A(n_358), .Y(n_1214) );
INVx2_ASAP7_75t_L g1313 ( .A(n_358), .Y(n_1313) );
INVx8_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g509 ( .A(n_359), .B(n_496), .Y(n_509) );
BUFx2_ASAP7_75t_L g1143 ( .A(n_359), .Y(n_1143) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_369), .B2(n_370), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_363), .A2(n_385), .B1(n_419), .B2(n_425), .Y(n_418) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx4_ASAP7_75t_L g768 ( .A(n_365), .Y(n_768) );
INVx2_ASAP7_75t_L g770 ( .A(n_365), .Y(n_770) );
INVx2_ASAP7_75t_L g1096 ( .A(n_365), .Y(n_1096) );
INVx4_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g375 ( .A(n_367), .Y(n_375) );
BUFx3_ASAP7_75t_L g814 ( .A(n_367), .Y(n_814) );
INVx2_ASAP7_75t_L g1032 ( .A(n_367), .Y(n_1032) );
BUFx2_ASAP7_75t_L g1270 ( .A(n_367), .Y(n_1270) );
AND2x2_ASAP7_75t_L g536 ( .A(n_368), .B(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_368), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_369), .A2(n_386), .B1(n_430), .B2(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g791 ( .A(n_370), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_370), .A2(n_1270), .B1(n_1387), .B2(n_1390), .Y(n_1397) );
BUFx4f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx4_ASAP7_75t_L g487 ( .A(n_371), .Y(n_487) );
BUFx4f_ASAP7_75t_L g815 ( .A(n_371), .Y(n_815) );
BUFx6f_ASAP7_75t_L g833 ( .A(n_371), .Y(n_833) );
OR2x6_ASAP7_75t_L g953 ( .A(n_371), .B(n_954), .Y(n_953) );
BUFx4f_ASAP7_75t_L g1094 ( .A(n_371), .Y(n_1094) );
BUFx4f_ASAP7_75t_L g1217 ( .A(n_371), .Y(n_1217) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx3_ASAP7_75t_L g379 ( .A(n_372), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B1(n_377), .B2(n_380), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g948 ( .A1(n_374), .A2(n_815), .B1(n_949), .B2(n_950), .C(n_951), .Y(n_948) );
OAI22xp5_ASAP7_75t_SL g1308 ( .A1(n_374), .A2(n_833), .B1(n_1297), .B2(n_1301), .Y(n_1308) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g603 ( .A1(n_377), .A2(n_604), .B(n_605), .C(n_608), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_377), .A2(n_739), .B1(n_759), .B2(n_768), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_377), .A2(n_1011), .B1(n_1015), .B2(n_1029), .Y(n_1028) );
OAI22xp33_ASAP7_75t_L g1033 ( .A1(n_377), .A2(n_1008), .B1(n_1021), .B2(n_1034), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_377), .A2(n_1080), .B1(n_1090), .B2(n_1096), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1219 ( .A1(n_377), .A2(n_1031), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
INVx5_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
BUFx3_ASAP7_75t_L g703 ( .A(n_379), .Y(n_703) );
BUFx2_ASAP7_75t_SL g771 ( .A(n_379), .Y(n_771) );
OR2x2_ASAP7_75t_L g937 ( .A(n_379), .B(n_936), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_385), .B1(n_386), .B2(n_387), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g1141 ( .A1(n_382), .A2(n_1142), .B1(n_1143), .B2(n_1144), .C(n_1145), .Y(n_1141) );
OAI22xp33_ASAP7_75t_L g1307 ( .A1(n_382), .A2(n_387), .B1(n_1294), .B2(n_1304), .Y(n_1307) );
OAI22xp33_ASAP7_75t_L g1312 ( .A1(n_382), .A2(n_1299), .B1(n_1302), .B2(n_1313), .Y(n_1312) );
OAI22xp33_ASAP7_75t_L g1358 ( .A1(n_382), .A2(n_1214), .B1(n_1340), .B2(n_1351), .Y(n_1358) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
BUFx3_ASAP7_75t_L g773 ( .A(n_384), .Y(n_773) );
BUFx3_ASAP7_75t_L g810 ( .A(n_384), .Y(n_810) );
BUFx6f_ASAP7_75t_L g1266 ( .A(n_384), .Y(n_1266) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_387), .A2(n_1036), .B1(n_1083), .B2(n_1087), .Y(n_1097) );
OAI22xp33_ASAP7_75t_L g1278 ( .A1(n_387), .A2(n_764), .B1(n_1279), .B2(n_1280), .Y(n_1278) );
INVx5_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx6_ASAP7_75t_L g774 ( .A(n_388), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g947 ( .A1(n_389), .A2(n_948), .B(n_953), .Y(n_947) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g775 ( .A(n_390), .Y(n_775) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx4_ASAP7_75t_L g607 ( .A(n_391), .Y(n_607) );
INVx1_ASAP7_75t_SL g1132 ( .A(n_391), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_391), .B(n_392), .Y(n_1224) );
AND2x2_ASAP7_75t_SL g1277 ( .A(n_391), .B(n_394), .Y(n_1277) );
INVx4_ASAP7_75t_L g1661 ( .A(n_391), .Y(n_1661) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g399 ( .A(n_394), .B(n_400), .Y(n_399) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_394), .Y(n_476) );
OR2x2_ASAP7_75t_L g543 ( .A(n_394), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g513 ( .A(n_395), .Y(n_513) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI33xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_403), .A3(n_418), .B1(n_429), .B2(n_437), .B3(n_442), .Y(n_397) );
OAI33xp33_ASAP7_75t_L g1292 ( .A1(n_398), .A2(n_756), .A3(n_1293), .B1(n_1296), .B2(n_1300), .B3(n_1303), .Y(n_1292) );
BUFx8_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx4f_ASAP7_75t_L g630 ( .A(n_399), .Y(n_630) );
BUFx4f_ASAP7_75t_L g680 ( .A(n_399), .Y(n_680) );
BUFx2_ASAP7_75t_L g1282 ( .A(n_399), .Y(n_1282) );
BUFx2_ASAP7_75t_L g997 ( .A(n_400), .Y(n_997) );
NAND2xp33_ASAP7_75t_SL g400 ( .A(n_401), .B(n_402), .Y(n_400) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_401), .Y(n_474) );
INVx1_ASAP7_75t_L g526 ( .A(n_401), .Y(n_526) );
AND3x4_ASAP7_75t_L g923 ( .A(n_401), .B(n_460), .C(n_728), .Y(n_923) );
INVx3_ASAP7_75t_L g438 ( .A(n_402), .Y(n_438) );
BUFx3_ASAP7_75t_L g460 ( .A(n_402), .Y(n_460) );
OAI22xp33_ASAP7_75t_L g1293 ( .A1(n_404), .A2(n_749), .B1(n_1294), .B2(n_1295), .Y(n_1293) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g1007 ( .A(n_406), .Y(n_1007) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x4_ASAP7_75t_L g448 ( .A(n_407), .B(n_438), .Y(n_448) );
OR2x4_ASAP7_75t_L g468 ( .A(n_407), .B(n_451), .Y(n_468) );
INVx2_ASAP7_75t_L g540 ( .A(n_407), .Y(n_540) );
BUFx3_ASAP7_75t_L g754 ( .A(n_407), .Y(n_754) );
BUFx4f_ASAP7_75t_L g918 ( .A(n_407), .Y(n_918) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_408), .Y(n_417) );
INVx2_ASAP7_75t_L g424 ( .A(n_408), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_408), .B(n_416), .Y(n_428) );
AND2x4_ASAP7_75t_L g455 ( .A(n_408), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g524 ( .A(n_409), .Y(n_524) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g423 ( .A(n_410), .Y(n_423) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_SL g1101 ( .A(n_412), .Y(n_1101) );
INVxp67_ASAP7_75t_SL g1395 ( .A(n_412), .Y(n_1395) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g1047 ( .A(n_413), .Y(n_1047) );
BUFx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_414), .Y(n_445) );
BUFx3_ASAP7_75t_L g751 ( .A(n_414), .Y(n_751) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
BUFx2_ASAP7_75t_L g464 ( .A(n_415), .Y(n_464) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g456 ( .A(n_416), .Y(n_456) );
BUFx2_ASAP7_75t_L g461 ( .A(n_417), .Y(n_461) );
INVx2_ASAP7_75t_L g560 ( .A(n_417), .Y(n_560) );
AND2x4_ASAP7_75t_L g638 ( .A(n_417), .B(n_566), .Y(n_638) );
OAI221xp5_ASAP7_75t_L g843 ( .A1(n_419), .A2(n_425), .B1(n_822), .B2(n_844), .C(n_845), .Y(n_843) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g548 ( .A(n_420), .B(n_542), .Y(n_548) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g636 ( .A(n_421), .Y(n_636) );
BUFx2_ASAP7_75t_L g682 ( .A(n_421), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g1648 ( .A1(n_421), .A2(n_433), .B1(n_1649), .B2(n_1650), .C(n_1651), .Y(n_1648) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_422), .Y(n_432) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_422), .Y(n_743) );
BUFx8_ASAP7_75t_L g915 ( .A(n_422), .Y(n_915) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
AND2x4_ASAP7_75t_L g523 ( .A(n_424), .B(n_524), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g671 ( .A1(n_425), .A2(n_672), .B1(n_673), .B2(n_674), .C(n_675), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g835 ( .A1(n_425), .A2(n_836), .B1(n_838), .B2(n_839), .C(n_840), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_425), .A2(n_992), .B1(n_993), .B2(n_994), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g1300 ( .A1(n_425), .A2(n_758), .B1(n_1301), .B2(n_1302), .Y(n_1300) );
OAI221xp5_ASAP7_75t_L g1652 ( .A1(n_425), .A2(n_622), .B1(n_1653), .B2(n_1654), .C(n_1655), .Y(n_1652) );
CKINVDCx8_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g684 ( .A(n_426), .Y(n_684) );
INVx3_ASAP7_75t_L g1018 ( .A(n_426), .Y(n_1018) );
INVx3_ASAP7_75t_L g1233 ( .A(n_426), .Y(n_1233) );
INVx1_ASAP7_75t_L g1285 ( .A(n_426), .Y(n_1285) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g571 ( .A(n_427), .Y(n_571) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g436 ( .A(n_428), .Y(n_436) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g450 ( .A(n_432), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g622 ( .A(n_432), .Y(n_622) );
BUFx6f_ASAP7_75t_L g837 ( .A(n_432), .Y(n_837) );
INVx1_ASAP7_75t_L g1298 ( .A(n_432), .Y(n_1298) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_433), .A2(n_622), .B1(n_623), .B2(n_624), .C(n_625), .Y(n_621) );
OAI22xp33_ASAP7_75t_SL g738 ( .A1(n_433), .A2(n_739), .B1(n_740), .B2(n_744), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g1296 ( .A1(n_433), .A2(n_1297), .B1(n_1298), .B2(n_1299), .Y(n_1296) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OR2x6_ASAP7_75t_L g471 ( .A(n_436), .B(n_438), .Y(n_471) );
BUFx3_ASAP7_75t_L g760 ( .A(n_436), .Y(n_760) );
INVx3_ASAP7_75t_L g644 ( .A(n_437), .Y(n_644) );
INVx3_ASAP7_75t_L g1718 ( .A(n_437), .Y(n_1718) );
NAND3x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .C(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g451 ( .A(n_438), .Y(n_451) );
AND2x4_ASAP7_75t_L g454 ( .A(n_438), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g525 ( .A(n_438), .B(n_526), .Y(n_525) );
NAND2x1p5_ASAP7_75t_L g990 ( .A(n_438), .B(n_441), .Y(n_990) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g558 ( .A(n_440), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_440), .B(n_535), .Y(n_936) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g911 ( .A(n_444), .Y(n_911) );
INVx2_ASAP7_75t_L g988 ( .A(n_444), .Y(n_988) );
INVx1_ASAP7_75t_L g1328 ( .A(n_444), .Y(n_1328) );
INVx4_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g574 ( .A(n_445), .B(n_543), .Y(n_574) );
INVx3_ASAP7_75t_L g921 ( .A(n_445), .Y(n_921) );
BUFx6f_ASAP7_75t_L g1352 ( .A(n_445), .Y(n_1352) );
OAI31xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_452), .A3(n_466), .B(n_472), .Y(n_446) );
INVx2_ASAP7_75t_SL g665 ( .A(n_448), .Y(n_665) );
INVx1_ASAP7_75t_L g779 ( .A(n_448), .Y(n_779) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_448), .Y(n_1108) );
INVx2_ASAP7_75t_SL g1414 ( .A(n_448), .Y(n_1414) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_450), .A2(n_652), .B1(n_653), .B2(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g1054 ( .A(n_450), .Y(n_1054) );
INVx1_ASAP7_75t_L g1109 ( .A(n_450), .Y(n_1109) );
INVx2_ASAP7_75t_L g1372 ( .A(n_450), .Y(n_1372) );
CKINVDCx8_ASAP7_75t_R g453 ( .A(n_454), .Y(n_453) );
CKINVDCx8_ASAP7_75t_R g668 ( .A(n_454), .Y(n_668) );
OAI31xp33_ASAP7_75t_L g848 ( .A1(n_454), .A2(n_849), .A3(n_860), .B(n_862), .Y(n_848) );
BUFx2_ASAP7_75t_L g629 ( .A(n_455), .Y(n_629) );
BUFx2_ASAP7_75t_L g633 ( .A(n_455), .Y(n_633) );
INVx2_ASAP7_75t_L g643 ( .A(n_455), .Y(n_643) );
BUFx2_ASAP7_75t_L g662 ( .A(n_455), .Y(n_662) );
BUFx2_ASAP7_75t_L g846 ( .A(n_455), .Y(n_846) );
BUFx3_ASAP7_75t_L g852 ( .A(n_455), .Y(n_852) );
BUFx2_ASAP7_75t_L g1161 ( .A(n_455), .Y(n_1161) );
INVx1_ASAP7_75t_L g566 ( .A(n_456), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_462), .B1(n_463), .B2(n_465), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_458), .A2(n_463), .B1(n_858), .B2(n_859), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_458), .A2(n_463), .B1(n_1248), .B2(n_1259), .Y(n_1258) );
AOI22xp33_ASAP7_75t_SL g1329 ( .A1(n_458), .A2(n_463), .B1(n_1320), .B2(n_1330), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g1374 ( .A1(n_458), .A2(n_463), .B1(n_1365), .B2(n_1375), .Y(n_1374) );
AOI22xp33_ASAP7_75t_SL g1419 ( .A1(n_458), .A2(n_463), .B1(n_1407), .B2(n_1420), .Y(n_1419) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
AND2x4_ASAP7_75t_L g463 ( .A(n_459), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g658 ( .A(n_459), .B(n_461), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g849 ( .A1(n_459), .A2(n_850), .B(n_853), .C(n_857), .Y(n_849) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_462), .A2(n_495), .B1(n_498), .B2(n_503), .Y(n_494) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_463), .Y(n_660) );
BUFx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g667 ( .A(n_468), .Y(n_667) );
BUFx2_ASAP7_75t_L g785 ( .A(n_468), .Y(n_785) );
BUFx2_ASAP7_75t_L g861 ( .A(n_468), .Y(n_861) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g654 ( .A(n_471), .Y(n_654) );
BUFx3_ASAP7_75t_L g1044 ( .A(n_471), .Y(n_1044) );
INVx1_ASAP7_75t_L g1333 ( .A(n_471), .Y(n_1333) );
OAI31xp33_ASAP7_75t_L g776 ( .A1(n_472), .A2(n_777), .A3(n_780), .B(n_784), .Y(n_776) );
OAI31xp33_ASAP7_75t_L g1042 ( .A1(n_472), .A2(n_1043), .A3(n_1045), .B(n_1052), .Y(n_1042) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
AND2x4_ASAP7_75t_L g669 ( .A(n_473), .B(n_475), .Y(n_669) );
AND2x2_ASAP7_75t_L g862 ( .A(n_473), .B(n_475), .Y(n_862) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_473), .B(n_475), .Y(n_1261) );
AND2x2_ASAP7_75t_SL g1736 ( .A(n_473), .B(n_475), .Y(n_1736) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI31xp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_485), .A3(n_504), .B(n_510), .Y(n_477) );
INVx4_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g788 ( .A(n_480), .Y(n_788) );
INVx3_ASAP7_75t_SL g1058 ( .A(n_480), .Y(n_1058) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_483), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_483), .Y(n_552) );
INVx2_ASAP7_75t_L g706 ( .A(n_483), .Y(n_706) );
BUFx3_ASAP7_75t_L g893 ( .A(n_483), .Y(n_893) );
NAND2xp5_ASAP7_75t_SL g885 ( .A(n_486), .B(n_886), .Y(n_885) );
OAI22xp5_ASAP7_75t_SL g1268 ( .A1(n_486), .A2(n_1269), .B1(n_1270), .B2(n_1271), .Y(n_1268) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g890 ( .A(n_487), .Y(n_890) );
INVx2_ASAP7_75t_L g897 ( .A(n_487), .Y(n_897) );
INVx2_ASAP7_75t_L g1274 ( .A(n_487), .Y(n_1274) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g1405 ( .A(n_489), .Y(n_1405) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AND2x2_ASAP7_75t_L g793 ( .A(n_490), .B(n_581), .Y(n_793) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g599 ( .A(n_492), .Y(n_599) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_493), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_495), .A2(n_498), .B1(n_782), .B2(n_795), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_495), .A2(n_1070), .B1(n_1320), .B2(n_1321), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_495), .A2(n_1365), .B1(n_1366), .B2(n_1367), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_495), .A2(n_1366), .B1(n_1407), .B2(n_1408), .Y(n_1406) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
AND2x4_ASAP7_75t_L g1069 ( .A(n_496), .B(n_497), .Y(n_1069) );
INVx1_ASAP7_75t_L g596 ( .A(n_497), .Y(n_596) );
BUFx2_ASAP7_75t_L g887 ( .A(n_497), .Y(n_887) );
INVx1_ASAP7_75t_L g960 ( .A(n_497), .Y(n_960) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g1071 ( .A(n_500), .Y(n_1071) );
BUFx3_ASAP7_75t_L g1194 ( .A(n_500), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_500), .A2(n_1069), .B1(n_1248), .B2(n_1249), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_501), .B(n_602), .Y(n_723) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g1061 ( .A(n_506), .Y(n_1061) );
BUFx2_ASAP7_75t_L g1323 ( .A(n_506), .Y(n_1323) );
HB1xp67_ASAP7_75t_L g1699 ( .A(n_506), .Y(n_1699) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g797 ( .A(n_508), .Y(n_797) );
INVx1_ASAP7_75t_L g1700 ( .A(n_508), .Y(n_1700) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g1064 ( .A(n_509), .Y(n_1064) );
INVx1_ASAP7_75t_L g1189 ( .A(n_509), .Y(n_1189) );
OAI31xp33_ASAP7_75t_L g786 ( .A1(n_510), .A2(n_787), .A3(n_789), .B(n_796), .Y(n_786) );
OAI31xp33_ASAP7_75t_L g1314 ( .A1(n_510), .A2(n_1315), .A3(n_1316), .B(n_1322), .Y(n_1314) );
BUFx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_SL g1073 ( .A(n_511), .Y(n_1073) );
INVx1_ASAP7_75t_L g1183 ( .A(n_511), .Y(n_1183) );
OAI31xp33_ASAP7_75t_L g1362 ( .A1(n_511), .A2(n_1363), .A3(n_1368), .B(n_1369), .Y(n_1362) );
BUFx2_ASAP7_75t_L g1410 ( .A(n_511), .Y(n_1410) );
OAI31xp33_ASAP7_75t_L g1691 ( .A1(n_511), .A2(n_1692), .A3(n_1696), .B(n_1698), .Y(n_1691) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVxp67_ASAP7_75t_L g527 ( .A(n_513), .Y(n_527) );
INVx1_ASAP7_75t_L g533 ( .A(n_513), .Y(n_533) );
OR2x2_ASAP7_75t_L g961 ( .A(n_513), .B(n_723), .Y(n_961) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
XOR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_647), .Y(n_515) );
INVx1_ASAP7_75t_L g645 ( .A(n_517), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .C(n_553), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_519), .A2(n_612), .B1(n_615), .B2(n_616), .Y(n_611) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OR2x6_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
OR2x2_ASAP7_75t_L g1644 ( .A(n_522), .B(n_527), .Y(n_1644) );
NAND2x1p5_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
BUFx3_ASAP7_75t_L g628 ( .A(n_523), .Y(n_628) );
INVx8_ASAP7_75t_L g641 ( .A(n_523), .Y(n_641) );
BUFx3_ASAP7_75t_L g677 ( .A(n_523), .Y(n_677) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_523), .Y(n_977) );
AND2x4_ASAP7_75t_L g557 ( .A(n_525), .B(n_558), .Y(n_557) );
AND2x6_ASAP7_75t_L g968 ( .A(n_525), .B(n_559), .Y(n_968) );
AND2x2_ASAP7_75t_L g970 ( .A(n_525), .B(n_565), .Y(n_970) );
INVx1_ASAP7_75t_L g974 ( .A(n_525), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B1(n_545), .B2(n_546), .Y(n_528) );
INVxp67_ASAP7_75t_L g871 ( .A(n_530), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_538), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_532), .A2(n_550), .B1(n_963), .B2(n_964), .Y(n_962) );
AND2x4_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
AND2x4_ASAP7_75t_L g550 ( .A(n_533), .B(n_551), .Y(n_550) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_534), .Y(n_696) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x2_ASAP7_75t_L g551 ( .A(n_535), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g612 ( .A(n_535), .B(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_SL g617 ( .A(n_535), .B(n_581), .Y(n_617) );
AND2x4_ASAP7_75t_L g700 ( .A(n_535), .B(n_552), .Y(n_700) );
BUFx2_ASAP7_75t_L g816 ( .A(n_535), .Y(n_816) );
AND2x4_ASAP7_75t_L g1127 ( .A(n_535), .B(n_709), .Y(n_1127) );
INVx3_ASAP7_75t_L g586 ( .A(n_536), .Y(n_586) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_536), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_536), .B(n_602), .Y(n_717) );
OR2x6_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_539), .B(n_541), .Y(n_1176) );
INVx2_ASAP7_75t_SL g1239 ( .A(n_539), .Y(n_1239) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
INVx3_ASAP7_75t_L g747 ( .A(n_540), .Y(n_747) );
INVxp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g570 ( .A(n_543), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g1179 ( .A(n_543), .Y(n_1179) );
INVx1_ASAP7_75t_L g985 ( .A(n_544), .Y(n_985) );
INVx1_ASAP7_75t_L g872 ( .A(n_546), .Y(n_872) );
NAND2x1_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g579 ( .A(n_552), .Y(n_579) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_552), .Y(n_606) );
NOR3xp33_ASAP7_75t_SL g553 ( .A(n_554), .B(n_575), .C(n_620), .Y(n_553) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_SL g556 ( .A(n_557), .B(n_559), .Y(n_556) );
AND2x4_ASAP7_75t_SL g562 ( .A(n_557), .B(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g632 ( .A(n_557), .B(n_633), .Y(n_632) );
NAND2x1_ASAP7_75t_L g876 ( .A(n_557), .B(n_559), .Y(n_876) );
AND2x4_ASAP7_75t_L g878 ( .A(n_557), .B(n_563), .Y(n_878) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_557), .B(n_559), .Y(n_1173) );
OR2x2_ASAP7_75t_L g932 ( .A(n_558), .B(n_717), .Y(n_932) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_572), .B2(n_573), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_568), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g1151 ( .A(n_570), .B(n_932), .Y(n_1151) );
BUFx3_ASAP7_75t_L g1348 ( .A(n_571), .Y(n_1348) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_572), .A2(n_593), .B1(n_595), .B2(n_597), .C(n_598), .Y(n_592) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g1154 ( .A(n_574), .B(n_961), .Y(n_1154) );
AND2x4_ASAP7_75t_L g1643 ( .A(n_574), .B(n_961), .Y(n_1643) );
AOI31xp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_603), .A3(n_611), .B(n_618), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_584), .B(n_589), .Y(n_576) );
INVx2_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
BUFx2_ASAP7_75t_L g942 ( .A(n_580), .Y(n_942) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x6_ASAP7_75t_L g724 ( .A(n_581), .B(n_602), .Y(n_724) );
BUFx3_ASAP7_75t_L g1130 ( .A(n_581), .Y(n_1130) );
INVx1_ASAP7_75t_L g1147 ( .A(n_581), .Y(n_1147) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g713 ( .A(n_583), .Y(n_713) );
INVx1_ASAP7_75t_L g824 ( .A(n_583), .Y(n_824) );
INVx2_ASAP7_75t_L g1672 ( .A(n_583), .Y(n_1672) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_SL g591 ( .A(n_586), .Y(n_591) );
INVx1_ASAP7_75t_L g609 ( .A(n_586), .Y(n_609) );
INVx2_ASAP7_75t_L g952 ( .A(n_586), .Y(n_952) );
BUFx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx3_ASAP7_75t_L g610 ( .A(n_588), .Y(n_610) );
INVx2_ASAP7_75t_L g614 ( .A(n_588), .Y(n_614) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_588), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B(n_600), .Y(n_589) );
INVx1_ASAP7_75t_L g832 ( .A(n_593), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_593), .A2(n_877), .B1(n_887), .B2(n_888), .Y(n_886) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g831 ( .A(n_595), .Y(n_831) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2x1_ASAP7_75t_L g719 ( .A(n_596), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_SL g827 ( .A1(n_601), .A2(n_828), .B(n_829), .C(n_830), .Y(n_827) );
A2O1A1Ixp33_ASAP7_75t_L g883 ( .A1(n_601), .A2(n_829), .B(n_884), .C(n_885), .Y(n_883) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g720 ( .A(n_602), .Y(n_720) );
INVx2_ASAP7_75t_L g697 ( .A(n_612), .Y(n_697) );
AND2x4_ASAP7_75t_L g934 ( .A(n_613), .B(n_935), .Y(n_934) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g826 ( .A(n_614), .Y(n_826) );
AOI211xp5_ASAP7_75t_SL g715 ( .A1(n_616), .A2(n_659), .B(n_716), .C(n_724), .Y(n_715) );
BUFx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g903 ( .A(n_617), .Y(n_903) );
OAI31xp67_ASAP7_75t_L g965 ( .A1(n_618), .A2(n_966), .A3(n_975), .B(n_986), .Y(n_965) );
INVx2_ASAP7_75t_L g1674 ( .A(n_618), .Y(n_1674) );
BUFx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI211xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_630), .B(n_631), .C(n_634), .Y(n_620) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_629), .A2(n_907), .B1(n_981), .B2(n_982), .Y(n_980) );
OAI33xp33_ASAP7_75t_L g1003 ( .A1(n_630), .A2(n_691), .A3(n_1004), .B1(n_1010), .B2(n_1014), .B3(n_1019), .Y(n_1003) );
OAI33xp33_ASAP7_75t_L g1077 ( .A1(n_630), .A2(n_691), .A3(n_1078), .B1(n_1081), .B2(n_1084), .B3(n_1088), .Y(n_1077) );
OAI33xp33_ASAP7_75t_L g1228 ( .A1(n_630), .A2(n_691), .A3(n_1229), .B1(n_1232), .B2(n_1234), .B3(n_1237), .Y(n_1228) );
INVx2_ASAP7_75t_SL g1180 ( .A(n_631), .Y(n_1180) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_632), .A2(n_644), .B1(n_906), .B2(n_912), .C(n_922), .Y(n_905) );
HB1xp67_ASAP7_75t_L g1646 ( .A(n_632), .Y(n_1646) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_639), .C(n_644), .Y(n_634) );
INVx1_ASAP7_75t_L g672 ( .A(n_636), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_637), .A2(n_828), .B1(n_851), .B2(n_852), .Y(n_850) );
BUFx12f_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx3_ASAP7_75t_L g907 ( .A(n_638), .Y(n_907) );
INVx5_ASAP7_75t_L g1164 ( .A(n_638), .Y(n_1164) );
BUFx3_ASAP7_75t_L g1166 ( .A(n_638), .Y(n_1166) );
INVx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_641), .Y(n_841) );
INVx8_ASAP7_75t_L g855 ( .A(n_641), .Y(n_855) );
INVx2_ASAP7_75t_L g1677 ( .A(n_641), .Y(n_1677) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g678 ( .A(n_643), .Y(n_678) );
INVx2_ASAP7_75t_L g842 ( .A(n_643), .Y(n_842) );
INVx1_ASAP7_75t_L g1170 ( .A(n_643), .Y(n_1170) );
INVx2_ASAP7_75t_L g691 ( .A(n_644), .Y(n_691) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_644), .Y(n_756) );
INVx2_ASAP7_75t_L g847 ( .A(n_644), .Y(n_847) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_669), .B(n_670), .C(n_692), .Y(n_649) );
NAND4xp25_ASAP7_75t_L g650 ( .A(n_651), .B(n_655), .C(n_663), .D(n_668), .Y(n_650) );
INVx2_ASAP7_75t_L g1255 ( .A(n_654), .Y(n_1255) );
AOI222xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_659), .B2(n_660), .C1(n_661), .C2(n_662), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_657), .A2(n_660), .B1(n_782), .B2(n_783), .Y(n_781) );
BUFx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx3_ASAP7_75t_L g1049 ( .A(n_658), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_660), .A2(n_1049), .B1(n_1050), .B2(n_1051), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_660), .A2(n_1049), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_660), .A2(n_1049), .B1(n_1193), .B2(n_1201), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1733 ( .A1(n_660), .A2(n_1049), .B1(n_1694), .B2(n_1734), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_661), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g690 ( .A(n_662), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_666), .B2(n_667), .Y(n_663) );
INVx2_ASAP7_75t_L g1053 ( .A(n_665), .Y(n_1053) );
INVx2_ASAP7_75t_L g1106 ( .A(n_667), .Y(n_1106) );
INVx1_ASAP7_75t_L g1416 ( .A(n_667), .Y(n_1416) );
OAI31xp33_ASAP7_75t_L g1098 ( .A1(n_669), .A2(n_1099), .A3(n_1105), .B(n_1107), .Y(n_1098) );
CKINVDCx14_ASAP7_75t_R g1203 ( .A(n_669), .Y(n_1203) );
OAI31xp33_ASAP7_75t_L g1324 ( .A1(n_669), .A2(n_1325), .A3(n_1326), .B(n_1331), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_679), .B1(n_681), .B2(n_691), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_672), .A2(n_1216), .B1(n_1226), .B2(n_1233), .Y(n_1232) );
BUFx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g688 ( .A(n_677), .Y(n_688) );
INVx2_ASAP7_75t_SL g1160 ( .A(n_677), .Y(n_1160) );
OAI33xp33_ASAP7_75t_L g737 ( .A1(n_679), .A2(n_738), .A3(n_745), .B1(n_752), .B2(n_756), .B3(n_757), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g834 ( .A1(n_679), .A2(n_835), .B1(n_843), .B2(n_847), .Y(n_834) );
OAI33xp33_ASAP7_75t_L g1702 ( .A1(n_679), .A2(n_1703), .A3(n_1709), .B1(n_1712), .B2(n_1716), .B3(n_1719), .Y(n_1702) );
BUFx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI22xp5_ASAP7_75t_SL g1647 ( .A1(n_680), .A2(n_847), .B1(n_1648), .B2(n_1652), .Y(n_1647) );
OAI221xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_684), .B2(n_685), .C(n_686), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g1284 ( .A1(n_682), .A2(n_1269), .B1(n_1279), .B2(n_1285), .Y(n_1284) );
OAI22xp5_ASAP7_75t_L g1343 ( .A1(n_682), .A2(n_684), .B1(n_1344), .B2(n_1345), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_682), .A2(n_1347), .B1(n_1348), .B2(n_1349), .Y(n_1346) );
OAI22xp5_ASAP7_75t_L g1386 ( .A1(n_682), .A2(n_1285), .B1(n_1387), .B2(n_1388), .Y(n_1386) );
OAI211xp5_ASAP7_75t_SL g710 ( .A1(n_683), .A2(n_703), .B(n_711), .C(n_714), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_684), .A2(n_1218), .B1(n_1227), .B2(n_1235), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_684), .A2(n_1271), .B1(n_1280), .B2(n_1287), .Y(n_1286) );
OAI22xp5_ASAP7_75t_L g1389 ( .A1(n_684), .A2(n_1287), .B1(n_1390), .B2(n_1391), .Y(n_1389) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_715), .B(n_725), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_698), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_696), .A2(n_1135), .B1(n_1136), .B2(n_1137), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1665 ( .A1(n_696), .A2(n_700), .B1(n_1666), .B2(n_1667), .Y(n_1665) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
HB1xp67_ASAP7_75t_L g1137 ( .A(n_700), .Y(n_1137) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_704), .C(n_707), .Y(n_701) );
INVx1_ASAP7_75t_L g1318 ( .A(n_703), .Y(n_1318) );
OAI22xp5_ASAP7_75t_L g1359 ( .A1(n_703), .A2(n_1270), .B1(n_1344), .B2(n_1347), .Y(n_1359) );
OAI22xp5_ASAP7_75t_L g1360 ( .A1(n_703), .A2(n_1270), .B1(n_1341), .B2(n_1353), .Y(n_1360) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g712 ( .A(n_706), .Y(n_712) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_708), .Y(n_829) );
INVx3_ASAP7_75t_L g1664 ( .A(n_708), .Y(n_1664) );
INVx2_ASAP7_75t_L g941 ( .A(n_712), .Y(n_941) );
BUFx2_ASAP7_75t_L g1140 ( .A(n_718), .Y(n_1140) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI21xp5_ASAP7_75t_SL g1128 ( .A1(n_724), .A2(n_1129), .B(n_1133), .Y(n_1128) );
AOI21xp5_ASAP7_75t_L g1659 ( .A1(n_724), .A2(n_1660), .B(n_1662), .Y(n_1659) );
INVx1_ASAP7_75t_L g1148 ( .A(n_725), .Y(n_1148) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_726), .Y(n_904) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_727), .Y(n_806) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_776), .C(n_786), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_762), .Y(n_736) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g1012 ( .A(n_741), .Y(n_1012) );
INVx8_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
BUFx3_ASAP7_75t_L g758 ( .A(n_742), .Y(n_758) );
INVx5_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_743), .A2(n_854), .B1(n_855), .B2(n_856), .Y(n_853) );
INVx3_ASAP7_75t_L g979 ( .A(n_743), .Y(n_979) );
HB1xp67_ASAP7_75t_L g1236 ( .A(n_743), .Y(n_1236) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_744), .A2(n_761), .B1(n_773), .B2(n_774), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_745) );
OAI22xp33_ASAP7_75t_L g763 ( .A1(n_746), .A2(n_753), .B1(n_764), .B2(n_765), .Y(n_763) );
BUFx4f_ASAP7_75t_SL g910 ( .A(n_747), .Y(n_910) );
OAI22xp33_ASAP7_75t_L g1283 ( .A1(n_747), .A2(n_920), .B1(n_1265), .B2(n_1273), .Y(n_1283) );
OAI22xp33_ASAP7_75t_L g1288 ( .A1(n_747), .A2(n_751), .B1(n_1267), .B2(n_1275), .Y(n_1288) );
OAI22xp33_ASAP7_75t_L g1350 ( .A1(n_747), .A2(n_1351), .B1(n_1352), .B2(n_1353), .Y(n_1350) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_748), .A2(n_755), .B1(n_770), .B2(n_771), .Y(n_769) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_749), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_752) );
OAI22xp33_ASAP7_75t_L g1088 ( .A1(n_749), .A2(n_1006), .B1(n_1089), .B2(n_1090), .Y(n_1088) );
OAI22xp33_ASAP7_75t_L g1229 ( .A1(n_749), .A2(n_1208), .B1(n_1220), .B2(n_1230), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1719 ( .A1(n_749), .A2(n_1705), .B1(n_1720), .B2(n_1721), .Y(n_1719) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g1418 ( .A(n_750), .Y(n_1418) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx6f_ASAP7_75t_L g1009 ( .A(n_751), .Y(n_1009) );
OAI221xp5_ASAP7_75t_L g987 ( .A1(n_754), .A2(n_945), .B1(n_950), .B2(n_988), .C(n_989), .Y(n_987) );
OAI22xp33_ASAP7_75t_L g1392 ( .A1(n_754), .A2(n_1393), .B1(n_1394), .B2(n_1395), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_760), .A2(n_1011), .B1(n_1012), .B2(n_1013), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_760), .A2(n_1012), .B1(n_1082), .B2(n_1083), .Y(n_1081) );
OAI33xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_766), .A3(n_767), .B1(n_769), .B2(n_772), .B3(n_775), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g1361 ( .A1(n_764), .A2(n_1143), .B1(n_1345), .B2(n_1349), .Y(n_1361) );
OAI22xp5_ASAP7_75t_L g1400 ( .A1(n_764), .A2(n_1143), .B1(n_1388), .B2(n_1391), .Y(n_1400) );
INVx1_ASAP7_75t_L g946 ( .A(n_766), .Y(n_946) );
OAI33xp33_ASAP7_75t_L g1722 ( .A1(n_766), .A2(n_1222), .A3(n_1723), .B1(n_1727), .B2(n_1728), .B3(n_1729), .Y(n_1722) );
OAI22xp5_ASAP7_75t_L g1272 ( .A1(n_768), .A2(n_1273), .B1(n_1274), .B2(n_1275), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g1401 ( .A1(n_768), .A2(n_1274), .B1(n_1384), .B2(n_1394), .Y(n_1401) );
OAI22xp33_ASAP7_75t_L g1024 ( .A1(n_774), .A2(n_1005), .B1(n_1020), .B2(n_1025), .Y(n_1024) );
OAI22xp33_ASAP7_75t_L g1092 ( .A1(n_774), .A2(n_1025), .B1(n_1079), .B2(n_1089), .Y(n_1092) );
OAI33xp33_ASAP7_75t_L g1022 ( .A1(n_775), .A2(n_1023), .A3(n_1024), .B1(n_1028), .B2(n_1033), .B3(n_1035), .Y(n_1022) );
OAI33xp33_ASAP7_75t_L g1091 ( .A1(n_775), .A2(n_1023), .A3(n_1092), .B1(n_1093), .B2(n_1095), .B3(n_1097), .Y(n_1091) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g1066 ( .A(n_793), .Y(n_1066) );
INVx3_ASAP7_75t_L g1196 ( .A(n_793), .Y(n_1196) );
XOR2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_1118), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_863), .B1(n_1116), .B2(n_1117), .Y(n_799) );
INVx1_ASAP7_75t_L g1116 ( .A(n_800), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
XNOR2x1_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_848), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_807), .B(n_834), .Y(n_805) );
NAND4xp25_ASAP7_75t_L g807 ( .A(n_808), .B(n_817), .C(n_821), .D(n_827), .Y(n_807) );
OAI21xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_813), .B(n_816), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_810), .A2(n_811), .B1(n_944), .B2(n_945), .Y(n_943) );
INVx1_ASAP7_75t_L g1210 ( .A(n_810), .Y(n_1210) );
BUFx6f_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_814), .Y(n_1034) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_814), .A2(n_1082), .B1(n_1085), .B2(n_1094), .Y(n_1093) );
OAI211xp5_ASAP7_75t_SL g817 ( .A1(n_815), .A2(n_818), .B(n_819), .C(n_820), .Y(n_817) );
OAI211xp5_ASAP7_75t_SL g821 ( .A1(n_815), .A2(n_822), .B(n_823), .C(n_825), .Y(n_821) );
INVx2_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
INVx2_ASAP7_75t_L g992 ( .A(n_837), .Y(n_992) );
A2O1A1Ixp33_ASAP7_75t_L g971 ( .A1(n_841), .A2(n_852), .B(n_972), .C(n_973), .Y(n_971) );
INVx1_ASAP7_75t_L g1117 ( .A(n_863), .Y(n_1117) );
XNOR2xp5_ASAP7_75t_L g863 ( .A(n_864), .B(n_999), .Y(n_863) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_866), .B1(n_924), .B2(n_925), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_867), .Y(n_866) );
XNOR2x1_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
NOR2x1_ASAP7_75t_L g869 ( .A(n_870), .B(n_873), .Y(n_869) );
NAND3xp33_ASAP7_75t_SL g873 ( .A(n_874), .B(n_881), .C(n_905), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_877), .B1(n_878), .B2(n_879), .C(n_880), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_878), .A2(n_1172), .B1(n_1173), .B2(n_1174), .Y(n_1171) );
OAI21xp5_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_900), .B(n_904), .Y(n_881) );
NAND3xp33_ASAP7_75t_L g882 ( .A(n_883), .B(n_889), .C(n_895), .Y(n_882) );
OAI211xp5_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_891), .B(n_892), .C(n_894), .Y(n_889) );
OAI211xp5_ASAP7_75t_L g1670 ( .A1(n_890), .A2(n_1653), .B(n_1671), .C(n_1673), .Y(n_1670) );
OAI211xp5_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_897), .B(n_898), .C(n_899), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_896), .A2(n_909), .B1(n_910), .B2(n_911), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g1309 ( .A1(n_897), .A2(n_1295), .B1(n_1305), .B2(n_1310), .Y(n_1309) );
INVx2_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g1139 ( .A(n_902), .Y(n_1139) );
INVx2_ASAP7_75t_L g1669 ( .A(n_902), .Y(n_1669) );
INVx4_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g1339 ( .A1(n_910), .A2(n_1340), .B1(n_1341), .B2(n_1342), .Y(n_1339) );
OAI22xp33_ASAP7_75t_L g1382 ( .A1(n_910), .A2(n_1383), .B1(n_1384), .B2(n_1385), .Y(n_1382) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_SL g914 ( .A(n_915), .Y(n_914) );
INVx3_ASAP7_75t_L g1086 ( .A(n_915), .Y(n_1086) );
AND2x4_ASAP7_75t_L g1178 ( .A(n_915), .B(n_1179), .Y(n_1178) );
INVx2_ASAP7_75t_SL g1287 ( .A(n_915), .Y(n_1287) );
INVx3_ASAP7_75t_L g1713 ( .A(n_915), .Y(n_1713) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_918), .B1(n_919), .B2(n_920), .Y(n_916) );
INVx1_ASAP7_75t_L g1231 ( .A(n_918), .Y(n_1231) );
OAI211xp5_ASAP7_75t_L g995 ( .A1(n_920), .A2(n_949), .B(n_996), .C(n_998), .Y(n_995) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
BUFx3_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
AOI33xp33_ASAP7_75t_L g1157 ( .A1(n_923), .A2(n_1158), .A3(n_1162), .B1(n_1165), .B2(n_1167), .B3(n_1169), .Y(n_1157) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
XNOR2x1_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .Y(n_926) );
NAND4xp75_ASAP7_75t_L g928 ( .A(n_929), .B(n_938), .C(n_962), .D(n_965), .Y(n_928) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
AOI211x1_ASAP7_75t_L g938 ( .A1(n_939), .A2(n_946), .B(n_947), .C(n_957), .Y(n_938) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx2_ASAP7_75t_L g1131 ( .A(n_941), .Y(n_1131) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
NAND2x2_ASAP7_75t_L g958 ( .A(n_955), .B(n_959), .Y(n_958) );
INVx2_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx2_ASAP7_75t_SL g959 ( .A(n_960), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_963), .A2(n_964), .B1(n_977), .B2(n_978), .Y(n_976) );
INVx4_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx2_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
AOI21xp33_ASAP7_75t_L g975 ( .A1(n_976), .A2(n_980), .B(n_983), .Y(n_975) );
INVx2_ASAP7_75t_L g1016 ( .A(n_978), .Y(n_1016) );
INVx2_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
OAI21xp5_ASAP7_75t_SL g986 ( .A1(n_987), .A2(n_991), .B(n_995), .Y(n_986) );
HB1xp67_ASAP7_75t_L g1257 ( .A(n_988), .Y(n_1257) );
INVx3_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
XOR2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1074), .Y(n_999) );
AND3x1_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1042), .C(n_1055), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1022), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1004 ( .A1(n_1005), .A2(n_1006), .B1(n_1008), .B2(n_1009), .Y(n_1004) );
OAI22xp33_ASAP7_75t_L g1019 ( .A1(n_1006), .A2(n_1009), .B1(n_1020), .B2(n_1021), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g1078 ( .A1(n_1006), .A2(n_1009), .B1(n_1079), .B2(n_1080), .Y(n_1078) );
OAI22xp33_ASAP7_75t_L g1303 ( .A1(n_1006), .A2(n_1101), .B1(n_1304), .B2(n_1305), .Y(n_1303) );
INVx2_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
OAI22xp33_ASAP7_75t_L g1237 ( .A1(n_1009), .A2(n_1211), .B1(n_1221), .B2(n_1238), .Y(n_1237) );
OAI22xp5_ASAP7_75t_L g1709 ( .A1(n_1012), .A2(n_1233), .B1(n_1710), .B2(n_1711), .Y(n_1709) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_1013), .A2(n_1017), .B1(n_1036), .B2(n_1040), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_1015), .A2(n_1016), .B1(n_1017), .B2(n_1018), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_1018), .A2(n_1085), .B1(n_1086), .B2(n_1087), .Y(n_1084) );
INVx2_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
BUFx6f_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx3_ASAP7_75t_L g1726 ( .A(n_1027), .Y(n_1726) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1215 ( .A1(n_1031), .A2(n_1216), .B1(n_1217), .B2(n_1218), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g1727 ( .A1(n_1031), .A2(n_1217), .B1(n_1710), .B2(n_1714), .Y(n_1727) );
OAI22xp5_ASAP7_75t_L g1728 ( .A1(n_1031), .A2(n_1217), .B1(n_1706), .B2(n_1721), .Y(n_1728) );
INVx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
BUFx2_ASAP7_75t_L g1311 ( .A(n_1032), .Y(n_1311) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
BUFx3_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVxp67_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1047), .Y(n_1342) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1047), .Y(n_1385) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_1050), .A2(n_1068), .B1(n_1070), .B2(n_1072), .Y(n_1067) );
OAI31xp33_ASAP7_75t_SL g1055 ( .A1(n_1056), .A2(n_1059), .A3(n_1065), .B(n_1073), .Y(n_1055) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx2_ASAP7_75t_SL g1063 ( .A(n_1064), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_1068), .A2(n_1070), .B1(n_1103), .B2(n_1115), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_1068), .A2(n_1193), .B1(n_1194), .B2(n_1195), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g1693 ( .A1(n_1068), .A2(n_1194), .B1(n_1694), .B2(n_1695), .Y(n_1693) );
BUFx3_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx2_ASAP7_75t_L g1366 ( .A(n_1071), .Y(n_1366) );
OAI31xp33_ASAP7_75t_L g1110 ( .A1(n_1073), .A2(n_1111), .A3(n_1112), .B(n_1113), .Y(n_1110) );
OAI31xp33_ASAP7_75t_L g1245 ( .A1(n_1073), .A2(n_1246), .A3(n_1250), .B(n_1251), .Y(n_1245) );
AND3x1_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1098), .C(n_1110), .Y(n_1075) );
NOR2xp33_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1091), .Y(n_1076) );
HB1xp67_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
OA22x2_ASAP7_75t_L g1118 ( .A1(n_1119), .A2(n_1240), .B1(n_1241), .B2(n_1423), .Y(n_1118) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1119), .Y(n_1423) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
XNOR2xp5_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1181), .Y(n_1121) );
NAND3xp33_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1149), .C(n_1155), .Y(n_1123) );
OAI21xp33_ASAP7_75t_L g1124 ( .A1(n_1125), .A2(n_1138), .B(n_1148), .Y(n_1124) );
INVx2_ASAP7_75t_SL g1126 ( .A(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
AOI21xp33_ASAP7_75t_SL g1149 ( .A1(n_1150), .A2(n_1152), .B(n_1153), .Y(n_1149) );
AOI21xp5_ASAP7_75t_L g1640 ( .A1(n_1150), .A2(n_1641), .B(n_1642), .Y(n_1640) );
INVx8_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
NOR3xp33_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1175), .C(n_1180), .Y(n_1155) );
NAND2xp5_ASAP7_75t_SL g1156 ( .A(n_1157), .B(n_1171), .Y(n_1156) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
OAI33xp33_ASAP7_75t_L g1281 ( .A1(n_1168), .A2(n_1282), .A3(n_1283), .B1(n_1284), .B2(n_1286), .B3(n_1288), .Y(n_1281) );
OAI33xp33_ASAP7_75t_L g1338 ( .A1(n_1168), .A2(n_1282), .A3(n_1339), .B1(n_1343), .B2(n_1346), .B3(n_1350), .Y(n_1338) );
OAI33xp33_ASAP7_75t_L g1381 ( .A1(n_1168), .A2(n_1282), .A3(n_1382), .B1(n_1386), .B2(n_1389), .B3(n_1392), .Y(n_1381) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1675 ( .A1(n_1178), .A2(n_1666), .B1(n_1667), .B2(n_1676), .Y(n_1675) );
AND2x4_ASAP7_75t_L g1676 ( .A(n_1179), .B(n_1677), .Y(n_1676) );
OAI221xp5_ASAP7_75t_L g1182 ( .A1(n_1183), .A2(n_1184), .B1(n_1197), .B2(n_1203), .C(n_1204), .Y(n_1182) );
NOR3xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1190), .C(n_1191), .Y(n_1184) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx2_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
NOR3xp33_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1199), .C(n_1202), .Y(n_1197) );
NOR2xp33_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1228), .Y(n_1204) );
OAI33xp33_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1207), .A3(n_1215), .B1(n_1219), .B2(n_1222), .B3(n_1225), .Y(n_1205) );
OAI33xp33_ASAP7_75t_L g1263 ( .A1(n_1206), .A2(n_1264), .A3(n_1268), .B1(n_1272), .B2(n_1276), .B3(n_1278), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1207 ( .A1(n_1208), .A2(n_1209), .B1(n_1211), .B2(n_1212), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1225 ( .A1(n_1209), .A2(n_1212), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1723 ( .A1(n_1212), .A2(n_1704), .B1(n_1720), .B2(n_1724), .Y(n_1723) );
OAI22xp5_ASAP7_75t_L g1729 ( .A1(n_1212), .A2(n_1711), .B1(n_1715), .B2(n_1724), .Y(n_1729) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
OAI22xp33_ASAP7_75t_L g1264 ( .A1(n_1214), .A2(n_1265), .B1(n_1266), .B2(n_1267), .Y(n_1264) );
OAI22xp33_ASAP7_75t_L g1399 ( .A1(n_1214), .A2(n_1266), .B1(n_1383), .B2(n_1393), .Y(n_1399) );
INVx2_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1712 ( .A1(n_1233), .A2(n_1713), .B1(n_1714), .B2(n_1715), .Y(n_1712) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1239), .Y(n_1705) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
AOI22xp5_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1334), .B1(n_1421), .B2(n_1422), .Y(n_1241) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1242), .Y(n_1421) );
XNOR2xp5_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1289), .Y(n_1242) );
NAND3xp33_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1253), .C(n_1262), .Y(n_1244) );
OAI31xp33_ASAP7_75t_L g1253 ( .A1(n_1254), .A2(n_1256), .A3(n_1260), .B(n_1261), .Y(n_1253) );
OAI31xp33_ASAP7_75t_L g1370 ( .A1(n_1261), .A2(n_1371), .A3(n_1373), .B(n_1376), .Y(n_1370) );
OAI31xp33_ASAP7_75t_SL g1411 ( .A1(n_1261), .A2(n_1412), .A3(n_1415), .B(n_1417), .Y(n_1411) );
NOR2xp33_ASAP7_75t_SL g1262 ( .A(n_1263), .B(n_1281), .Y(n_1262) );
OAI33xp33_ASAP7_75t_L g1354 ( .A1(n_1276), .A2(n_1355), .A3(n_1358), .B1(n_1359), .B2(n_1360), .B3(n_1361), .Y(n_1354) );
OAI33xp33_ASAP7_75t_L g1396 ( .A1(n_1276), .A2(n_1397), .A3(n_1398), .B1(n_1399), .B2(n_1400), .B3(n_1401), .Y(n_1396) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
NAND3xp33_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1314), .C(n_1324), .Y(n_1290) );
NOR2xp33_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1306), .Y(n_1291) );
INVx4_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
HB1xp67_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1334), .Y(n_1422) );
XOR2xp5_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1377), .Y(n_1334) );
NAND3xp33_ASAP7_75t_L g1336 ( .A(n_1337), .B(n_1362), .C(n_1370), .Y(n_1336) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1354), .Y(n_1337) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1352), .Y(n_1708) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
INVx2_ASAP7_75t_SL g1356 ( .A(n_1357), .Y(n_1356) );
XNOR2xp5_ASAP7_75t_L g1377 ( .A(n_1378), .B(n_1379), .Y(n_1377) );
AND3x1_ASAP7_75t_L g1379 ( .A(n_1380), .B(n_1402), .C(n_1411), .Y(n_1379) );
NOR2xp33_ASAP7_75t_SL g1380 ( .A(n_1381), .B(n_1396), .Y(n_1380) );
OAI31xp33_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1404), .A3(n_1409), .B(n_1410), .Y(n_1402) );
INVx2_ASAP7_75t_SL g1413 ( .A(n_1414), .Y(n_1413) );
OAI221xp5_ASAP7_75t_L g1424 ( .A1(n_1425), .A2(n_1632), .B1(n_1635), .B2(n_1678), .C(n_1682), .Y(n_1424) );
AOI211xp5_ASAP7_75t_L g1425 ( .A1(n_1426), .A2(n_1546), .B(n_1592), .C(n_1616), .Y(n_1425) );
OAI211xp5_ASAP7_75t_L g1426 ( .A1(n_1427), .A2(n_1443), .B(n_1488), .C(n_1534), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1566 ( .A(n_1427), .B(n_1567), .Y(n_1566) );
OAI211xp5_ASAP7_75t_L g1616 ( .A1(n_1427), .A2(n_1617), .B(n_1619), .C(n_1625), .Y(n_1616) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
OAI221xp5_ASAP7_75t_L g1518 ( .A1(n_1428), .A2(n_1519), .B1(n_1525), .B2(n_1528), .C(n_1530), .Y(n_1518) );
OAI32xp33_ASAP7_75t_L g1584 ( .A1(n_1428), .A2(n_1489), .A3(n_1506), .B1(n_1541), .B2(n_1585), .Y(n_1584) );
OAI221xp5_ASAP7_75t_L g1592 ( .A1(n_1428), .A2(n_1517), .B1(n_1593), .B2(n_1600), .C(n_1602), .Y(n_1592) );
INVx3_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
INVx3_ASAP7_75t_L g1512 ( .A(n_1429), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1429), .B(n_1516), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1529 ( .A(n_1429), .B(n_1462), .Y(n_1529) );
OR2x2_ASAP7_75t_L g1551 ( .A(n_1429), .B(n_1484), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1429), .B(n_1475), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1608 ( .A(n_1429), .B(n_1500), .Y(n_1608) );
NAND2xp5_ASAP7_75t_L g1615 ( .A(n_1429), .B(n_1484), .Y(n_1615) );
NOR2xp33_ASAP7_75t_L g1620 ( .A(n_1429), .B(n_1621), .Y(n_1620) );
AND2x4_ASAP7_75t_SL g1429 ( .A(n_1430), .B(n_1437), .Y(n_1429) );
AND2x6_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1433), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1435 ( .A(n_1432), .B(n_1436), .Y(n_1435) );
AND2x4_ASAP7_75t_L g1438 ( .A(n_1432), .B(n_1439), .Y(n_1438) );
AND2x6_ASAP7_75t_L g1441 ( .A(n_1432), .B(n_1442), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1432), .B(n_1436), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1432), .B(n_1436), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1434), .B(n_1440), .Y(n_1439) );
INVx2_ASAP7_75t_L g1634 ( .A(n_1441), .Y(n_1634) );
OAI21xp5_ASAP7_75t_L g1737 ( .A1(n_1442), .A2(n_1738), .B(n_1739), .Y(n_1737) );
AOI221xp5_ASAP7_75t_L g1443 ( .A1(n_1444), .A2(n_1455), .B1(n_1466), .B2(n_1483), .C(n_1485), .Y(n_1443) );
A2O1A1Ixp33_ASAP7_75t_SL g1513 ( .A1(n_1444), .A2(n_1494), .B(n_1514), .C(n_1515), .Y(n_1513) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1444), .Y(n_1544) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1451), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
OR2x2_ASAP7_75t_L g1506 ( .A(n_1446), .B(n_1451), .Y(n_1506) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1470 ( .A(n_1447), .B(n_1471), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1447), .B(n_1471), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1447), .B(n_1472), .Y(n_1497) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1447), .Y(n_1509) );
NOR2xp33_ASAP7_75t_L g1521 ( .A(n_1447), .B(n_1451), .Y(n_1521) );
NAND2xp5_ASAP7_75t_L g1447 ( .A(n_1448), .B(n_1449), .Y(n_1447) );
NOR2xp33_ASAP7_75t_L g1468 ( .A(n_1451), .B(n_1458), .Y(n_1468) );
CKINVDCx5p33_ASAP7_75t_R g1482 ( .A(n_1451), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1451), .B(n_1458), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1524 ( .A(n_1451), .B(n_1481), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_1451), .B(n_1497), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1578 ( .A(n_1451), .B(n_1509), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1598 ( .A(n_1451), .B(n_1599), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1454), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_1452), .B(n_1454), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1461), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1456), .B(n_1508), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1456), .B(n_1521), .Y(n_1520) );
OR2x2_ASAP7_75t_L g1561 ( .A(n_1456), .B(n_1524), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1456), .B(n_1500), .Y(n_1591) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1456), .B(n_1489), .Y(n_1626) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1457), .B(n_1480), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_1457), .B(n_1486), .Y(n_1535) );
NOR2xp33_ASAP7_75t_L g1539 ( .A(n_1457), .B(n_1506), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_1457), .B(n_1489), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1457), .B(n_1553), .Y(n_1552) );
NAND2xp5_ASAP7_75t_L g1556 ( .A(n_1457), .B(n_1496), .Y(n_1556) );
NAND2xp5_ASAP7_75t_L g1564 ( .A(n_1457), .B(n_1491), .Y(n_1564) );
INVx3_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
INVx2_ASAP7_75t_L g1494 ( .A(n_1458), .Y(n_1494) );
NAND2xp5_ASAP7_75t_L g1579 ( .A(n_1458), .B(n_1462), .Y(n_1579) );
OR2x2_ASAP7_75t_L g1621 ( .A(n_1458), .B(n_1491), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1460), .Y(n_1458) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1462), .Y(n_1536) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1462), .B(n_1601), .Y(n_1600) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
OR2x2_ASAP7_75t_L g1483 ( .A(n_1463), .B(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1463), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_1463), .B(n_1484), .Y(n_1500) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1463), .Y(n_1517) );
NAND2xp5_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1465), .Y(n_1463) );
OAI32xp33_ASAP7_75t_L g1466 ( .A1(n_1467), .A2(n_1469), .A3(n_1475), .B1(n_1476), .B2(n_1479), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1468), .B(n_1486), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1469), .B(n_1527), .Y(n_1526) );
NAND2xp5_ASAP7_75t_SL g1541 ( .A(n_1469), .B(n_1494), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1469), .B(n_1482), .Y(n_1583) );
OAI21xp5_ASAP7_75t_L g1588 ( .A1(n_1469), .A2(n_1589), .B(n_1591), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1469), .B(n_1487), .Y(n_1595) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1471), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_1471), .B(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1472), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1474), .Y(n_1472) );
OAI21xp33_ASAP7_75t_L g1537 ( .A1(n_1475), .A2(n_1538), .B(n_1540), .Y(n_1537) );
AOI221xp5_ASAP7_75t_L g1625 ( .A1(n_1475), .A2(n_1507), .B1(n_1626), .B2(n_1627), .C(n_1628), .Y(n_1625) );
INVx2_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
AOI22xp33_ASAP7_75t_L g1519 ( .A1(n_1476), .A2(n_1520), .B1(n_1522), .B2(n_1523), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1522 ( .A(n_1476), .B(n_1491), .Y(n_1522) );
CKINVDCx6p67_ASAP7_75t_R g1570 ( .A(n_1476), .Y(n_1570) );
AND2x4_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1478), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1477), .B(n_1478), .Y(n_1484) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1482), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1482), .B(n_1497), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1501 ( .A(n_1482), .B(n_1502), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1482), .B(n_1508), .Y(n_1507) );
OR2x2_ASAP7_75t_L g1540 ( .A(n_1482), .B(n_1541), .Y(n_1540) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1482), .B(n_1605), .Y(n_1604) );
OR2x2_ASAP7_75t_L g1511 ( .A(n_1483), .B(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1483), .Y(n_1586) );
OR2x2_ASAP7_75t_L g1490 ( .A(n_1484), .B(n_1491), .Y(n_1490) );
AOI21xp33_ASAP7_75t_L g1559 ( .A1(n_1484), .A2(n_1530), .B(n_1560), .Y(n_1559) );
NAND2xp5_ASAP7_75t_SL g1575 ( .A(n_1484), .B(n_1576), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1484), .B(n_1512), .Y(n_1631) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1485), .Y(n_1571) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1485), .B(n_1516), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1485), .B(n_1517), .Y(n_1627) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1486), .B(n_1487), .Y(n_1485) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1486), .Y(n_1502) );
AOI211xp5_ASAP7_75t_L g1488 ( .A1(n_1489), .A2(n_1492), .B(n_1498), .C(n_1518), .Y(n_1488) );
INVx2_ASAP7_75t_SL g1489 ( .A(n_1490), .Y(n_1489) );
NOR2xp33_ASAP7_75t_L g1573 ( .A(n_1490), .B(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
OR2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1495), .Y(n_1493) );
INVx2_ASAP7_75t_L g1505 ( .A(n_1494), .Y(n_1505) );
NAND2xp5_ASAP7_75t_SL g1558 ( .A(n_1494), .B(n_1522), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1612 ( .A(n_1494), .B(n_1578), .Y(n_1612) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1497), .Y(n_1607) );
OAI211xp5_ASAP7_75t_L g1498 ( .A1(n_1499), .A2(n_1501), .B(n_1503), .C(n_1513), .Y(n_1498) );
CKINVDCx14_ASAP7_75t_R g1499 ( .A(n_1500), .Y(n_1499) );
NOR2xp33_ASAP7_75t_L g1548 ( .A(n_1501), .B(n_1511), .Y(n_1548) );
OR2x2_ASAP7_75t_L g1590 ( .A(n_1502), .B(n_1527), .Y(n_1590) );
OAI21xp5_ASAP7_75t_L g1503 ( .A1(n_1504), .A2(n_1507), .B(n_1510), .Y(n_1503) );
NOR2xp33_ASAP7_75t_L g1504 ( .A(n_1505), .B(n_1506), .Y(n_1504) );
AOI311xp33_ASAP7_75t_L g1580 ( .A1(n_1505), .A2(n_1550), .A3(n_1581), .B(n_1584), .C(n_1587), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1505), .B(n_1507), .Y(n_1614) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1507), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1508), .B(n_1527), .Y(n_1553) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1508), .Y(n_1606) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
NAND2xp5_ASAP7_75t_L g1585 ( .A(n_1512), .B(n_1586), .Y(n_1585) );
AOI221xp5_ASAP7_75t_L g1554 ( .A1(n_1515), .A2(n_1555), .B1(n_1557), .B2(n_1566), .C(n_1568), .Y(n_1554) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1516), .Y(n_1542) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
AOI21xp5_ASAP7_75t_L g1628 ( .A1(n_1525), .A2(n_1629), .B(n_1630), .Y(n_1628) );
CKINVDCx5p33_ASAP7_75t_R g1525 ( .A(n_1526), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1527), .B(n_1535), .Y(n_1603) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1530), .Y(n_1567) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1533), .Y(n_1531) );
AOI221xp5_ASAP7_75t_L g1534 ( .A1(n_1535), .A2(n_1536), .B1(n_1537), .B2(n_1542), .C(n_1543), .Y(n_1534) );
INVxp33_ASAP7_75t_SL g1538 ( .A(n_1539), .Y(n_1538) );
OAI31xp33_ASAP7_75t_L g1610 ( .A1(n_1542), .A2(n_1560), .A3(n_1589), .B(n_1611), .Y(n_1610) );
NOR2xp33_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1545), .Y(n_1543) );
OAI211xp5_ASAP7_75t_L g1557 ( .A1(n_1544), .A2(n_1558), .B(n_1559), .C(n_1562), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1581 ( .A(n_1544), .B(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1545), .Y(n_1622) );
NAND3xp33_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1554), .C(n_1580), .Y(n_1546) );
NOR2xp33_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1549), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1550), .B(n_1552), .Y(n_1549) );
AOI22xp33_ASAP7_75t_SL g1593 ( .A1(n_1550), .A2(n_1594), .B1(n_1596), .B2(n_1597), .Y(n_1593) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1553), .Y(n_1624) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
NAND2xp5_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1565), .Y(n_1562) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
OAI211xp5_ASAP7_75t_L g1568 ( .A1(n_1569), .A2(n_1571), .B(n_1572), .C(n_1575), .Y(n_1568) );
CKINVDCx6p67_ASAP7_75t_R g1569 ( .A(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
INVxp33_ASAP7_75t_SL g1629 ( .A(n_1576), .Y(n_1629) );
NOR2xp33_ASAP7_75t_L g1576 ( .A(n_1577), .B(n_1579), .Y(n_1576) );
CKINVDCx14_ASAP7_75t_R g1577 ( .A(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
INVxp67_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1590), .B(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
O2A1O1Ixp33_ASAP7_75t_L g1602 ( .A1(n_1603), .A2(n_1604), .B(n_1608), .C(n_1609), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1605 ( .A(n_1606), .B(n_1607), .Y(n_1605) );
AOI21xp5_ASAP7_75t_L g1609 ( .A1(n_1610), .A2(n_1613), .B(n_1615), .Y(n_1609) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
OAI21xp33_ASAP7_75t_L g1619 ( .A1(n_1620), .A2(n_1622), .B(n_1623), .Y(n_1619) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
CKINVDCx20_ASAP7_75t_R g1632 ( .A(n_1633), .Y(n_1632) );
CKINVDCx20_ASAP7_75t_R g1633 ( .A(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
HB1xp67_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
AND4x1_ASAP7_75t_L g1639 ( .A(n_1640), .B(n_1645), .C(n_1657), .D(n_1675), .Y(n_1639) );
NOR3xp33_ASAP7_75t_L g1645 ( .A(n_1646), .B(n_1647), .C(n_1656), .Y(n_1645) );
OAI21xp5_ASAP7_75t_L g1657 ( .A1(n_1658), .A2(n_1668), .B(n_1674), .Y(n_1657) );
INVx2_ASAP7_75t_SL g1663 ( .A(n_1664), .Y(n_1663) );
INVx2_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
BUFx3_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
HB1xp67_ASAP7_75t_SL g1683 ( .A(n_1684), .Y(n_1683) );
INVxp33_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
HB1xp67_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
NAND3xp33_ASAP7_75t_L g1690 ( .A(n_1691), .B(n_1701), .C(n_1730), .Y(n_1690) );
NOR2xp33_ASAP7_75t_SL g1701 ( .A(n_1702), .B(n_1722), .Y(n_1701) );
OAI22xp5_ASAP7_75t_L g1703 ( .A1(n_1704), .A2(n_1705), .B1(n_1706), .B2(n_1707), .Y(n_1703) );
INVx2_ASAP7_75t_SL g1707 ( .A(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1717), .Y(n_1716) );
BUFx2_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
INVx2_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
INVx2_ASAP7_75t_SL g1725 ( .A(n_1726), .Y(n_1725) );
OAI31xp33_ASAP7_75t_L g1730 ( .A1(n_1731), .A2(n_1732), .A3(n_1735), .B(n_1736), .Y(n_1730) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1740), .Y(n_1739) );
endmodule