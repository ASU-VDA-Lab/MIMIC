module real_aes_877_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_0), .B(n_159), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_1), .A2(n_141), .B(n_192), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_2), .A2(n_464), .B1(n_469), .B2(n_814), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_3), .B(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_4), .A2(n_11), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_4), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_5), .B(n_149), .Y(n_205) );
INVx1_ASAP7_75t_L g146 ( .A(n_6), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_7), .B(n_149), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_8), .A2(n_121), .B1(n_445), .B2(n_446), .Y(n_120) );
INVxp67_ASAP7_75t_L g446 ( .A(n_8), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_8), .B(n_136), .Y(n_505) );
INVx1_ASAP7_75t_L g533 ( .A(n_9), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_10), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_11), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_12), .Y(n_548) );
NAND2xp33_ASAP7_75t_L g186 ( .A(n_13), .B(n_153), .Y(n_186) );
INVx2_ASAP7_75t_L g138 ( .A(n_14), .Y(n_138) );
AOI221x1_ASAP7_75t_L g228 ( .A1(n_15), .A2(n_28), .B1(n_141), .B2(n_159), .C(n_229), .Y(n_228) );
AND3x1_ASAP7_75t_L g109 ( .A(n_16), .B(n_41), .C(n_110), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_16), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_17), .B(n_159), .Y(n_182) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_18), .A2(n_180), .B(n_181), .Y(n_179) );
INVx1_ASAP7_75t_L g514 ( .A(n_19), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_20), .B(n_172), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_21), .B(n_149), .Y(n_148) );
AO21x1_ASAP7_75t_L g200 ( .A1(n_22), .A2(n_159), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g108 ( .A(n_23), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_24), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g512 ( .A(n_25), .Y(n_512) );
INVx1_ASAP7_75t_SL g498 ( .A(n_26), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_27), .B(n_160), .Y(n_592) );
INVxp33_ASAP7_75t_L g823 ( .A(n_29), .Y(n_823) );
NAND2x1_ASAP7_75t_L g214 ( .A(n_30), .B(n_149), .Y(n_214) );
AOI33xp33_ASAP7_75t_L g560 ( .A1(n_31), .A2(n_56), .A3(n_488), .B1(n_495), .B2(n_561), .B3(n_562), .Y(n_560) );
NAND2x1_ASAP7_75t_L g168 ( .A(n_32), .B(n_153), .Y(n_168) );
INVx1_ASAP7_75t_L g542 ( .A(n_33), .Y(n_542) );
OR2x2_ASAP7_75t_L g137 ( .A(n_34), .B(n_90), .Y(n_137) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_34), .A2(n_90), .B(n_138), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_35), .B(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_36), .B(n_153), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_37), .B(n_149), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_38), .B(n_153), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_39), .A2(n_141), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g142 ( .A(n_40), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g157 ( .A(n_40), .B(n_146), .Y(n_157) );
INVx1_ASAP7_75t_L g494 ( .A(n_40), .Y(n_494) );
OR2x6_ASAP7_75t_L g452 ( .A(n_41), .B(n_453), .Y(n_452) );
XNOR2xp5_ASAP7_75t_L g465 ( .A(n_42), .B(n_466), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_43), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_44), .B(n_159), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_45), .B(n_486), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_46), .A2(n_136), .B1(n_176), .B2(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_47), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_48), .B(n_160), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_49), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_50), .B(n_153), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_51), .B(n_180), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_52), .B(n_160), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_53), .A2(n_141), .B(n_167), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_54), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_55), .B(n_153), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_57), .B(n_160), .Y(n_572) );
INVx1_ASAP7_75t_L g145 ( .A(n_58), .Y(n_145) );
INVx1_ASAP7_75t_L g155 ( .A(n_58), .Y(n_155) );
AND2x2_ASAP7_75t_L g573 ( .A(n_59), .B(n_172), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_60), .A2(n_77), .B1(n_486), .B2(n_492), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_61), .B(n_486), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_62), .B(n_149), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_63), .B(n_176), .Y(n_550) );
AOI21xp5_ASAP7_75t_SL g522 ( .A1(n_64), .A2(n_492), .B(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_65), .A2(n_141), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g508 ( .A(n_66), .Y(n_508) );
AO21x1_ASAP7_75t_L g202 ( .A1(n_67), .A2(n_141), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_68), .B(n_159), .Y(n_190) );
INVx1_ASAP7_75t_L g571 ( .A(n_69), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_70), .B(n_159), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_71), .A2(n_492), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g251 ( .A(n_72), .B(n_173), .Y(n_251) );
INVx1_ASAP7_75t_L g143 ( .A(n_73), .Y(n_143) );
INVx1_ASAP7_75t_L g151 ( .A(n_73), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_74), .A2(n_100), .B1(n_467), .B2(n_468), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_74), .Y(n_467) );
AND2x2_ASAP7_75t_L g174 ( .A(n_75), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_76), .B(n_486), .Y(n_563) );
AND2x2_ASAP7_75t_L g501 ( .A(n_78), .B(n_175), .Y(n_501) );
INVx1_ASAP7_75t_L g509 ( .A(n_79), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_80), .A2(n_492), .B(n_497), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g590 ( .A1(n_81), .A2(n_492), .B(n_555), .C(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_82), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g454 ( .A(n_82), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_83), .B(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g188 ( .A(n_84), .B(n_175), .Y(n_188) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_85), .B(n_175), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_86), .A2(n_492), .B1(n_558), .B2(n_559), .Y(n_557) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_87), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_87), .Y(n_123) );
XNOR2xp5_ASAP7_75t_L g464 ( .A(n_88), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g201 ( .A(n_89), .B(n_136), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_91), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g218 ( .A(n_92), .B(n_175), .Y(n_218) );
INVx1_ASAP7_75t_L g524 ( .A(n_93), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_94), .B(n_149), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_95), .A2(n_141), .B(n_147), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_96), .B(n_153), .Y(n_230) );
AND2x2_ASAP7_75t_L g564 ( .A(n_97), .B(n_175), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_98), .B(n_149), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_99), .A2(n_540), .B(n_541), .C(n_543), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_100), .Y(n_468) );
BUFx2_ASAP7_75t_L g118 ( .A(n_101), .Y(n_118) );
BUFx2_ASAP7_75t_SL g461 ( .A(n_101), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_102), .A2(n_141), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_103), .B(n_160), .Y(n_525) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_113), .B(n_822), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_105), .B(n_823), .Y(n_822) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_109), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_108), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OA22x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B1(n_458), .B2(n_462), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_447), .B(n_455), .Y(n_119) );
INVx1_ASAP7_75t_L g445 ( .A(n_121), .Y(n_445) );
XNOR2x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_128), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_128), .A2(n_470), .B1(n_474), .B2(n_477), .Y(n_469) );
INVx2_ASAP7_75t_L g819 ( .A(n_128), .Y(n_819) );
OR2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_343), .Y(n_128) );
NAND3xp33_ASAP7_75t_SL g129 ( .A(n_130), .B(n_255), .C(n_310), .Y(n_129) );
AOI221xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_195), .B1(n_219), .B2(n_223), .C(n_233), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_178), .Y(n_131) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_132), .B(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g254 ( .A(n_132), .Y(n_254) );
AND2x2_ASAP7_75t_L g299 ( .A(n_132), .B(n_236), .Y(n_299) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_163), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g287 ( .A(n_134), .Y(n_287) );
INVx1_ASAP7_75t_L g297 ( .A(n_134), .Y(n_297) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_139), .B(n_161), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_135), .B(n_162), .Y(n_161) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_135), .A2(n_139), .B(n_161), .Y(n_261) );
INVx1_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_136), .A2(n_182), .B(n_183), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_136), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_136), .B(n_156), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_136), .A2(n_522), .B(n_526), .Y(n_521) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_137), .B(n_138), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_158), .Y(n_139) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
BUFx3_ASAP7_75t_L g490 ( .A(n_142), .Y(n_490) );
AND2x6_ASAP7_75t_L g153 ( .A(n_143), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g496 ( .A(n_143), .Y(n_496) );
AND2x4_ASAP7_75t_L g492 ( .A(n_144), .B(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g149 ( .A(n_145), .B(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g488 ( .A(n_145), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_146), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_152), .B(n_156), .Y(n_147) );
INVxp67_ASAP7_75t_L g515 ( .A(n_149), .Y(n_515) );
AND2x4_ASAP7_75t_L g160 ( .A(n_150), .B(n_154), .Y(n_160) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVxp67_ASAP7_75t_L g513 ( .A(n_153), .Y(n_513) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_156), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_156), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_156), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_156), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_156), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_156), .A2(n_230), .B(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_156), .A2(n_248), .B(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_SL g497 ( .A1(n_156), .A2(n_498), .B(n_499), .C(n_500), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_156), .A2(n_499), .B(n_524), .C(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_156), .A2(n_499), .B(n_533), .C(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g558 ( .A(n_156), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_156), .A2(n_499), .B(n_571), .C(n_572), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_156), .A2(n_592), .B(n_593), .Y(n_591) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g159 ( .A(n_157), .B(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_157), .Y(n_543) );
INVx1_ASAP7_75t_L g510 ( .A(n_160), .Y(n_510) );
OR2x2_ASAP7_75t_L g276 ( .A(n_163), .B(n_179), .Y(n_276) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_163), .B(n_222), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_163), .B(n_187), .Y(n_320) );
INVx2_ASAP7_75t_L g329 ( .A(n_163), .Y(n_329) );
AND2x2_ASAP7_75t_L g350 ( .A(n_163), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g434 ( .A(n_163), .B(n_253), .Y(n_434) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g262 ( .A(n_164), .B(n_187), .Y(n_262) );
AND2x2_ASAP7_75t_L g395 ( .A(n_164), .B(n_222), .Y(n_395) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_164), .Y(n_421) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_171), .B(n_174), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_170), .Y(n_165) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_171), .A2(n_484), .B(n_501), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_172), .A2(n_190), .B(n_191), .Y(n_189) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_172), .A2(n_228), .B(n_232), .Y(n_227) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_172), .A2(n_228), .B(n_232), .Y(n_239) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx3_ASAP7_75t_L g217 ( .A(n_175), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_175), .A2(n_217), .B1(n_539), .B2(n_544), .Y(n_538) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_176), .B(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx4f_ASAP7_75t_L g180 ( .A(n_177), .Y(n_180) );
AND2x4_ASAP7_75t_L g349 ( .A(n_178), .B(n_350), .Y(n_349) );
AOI321xp33_ASAP7_75t_L g363 ( .A1(n_178), .A2(n_292), .A3(n_293), .B1(n_325), .B2(n_364), .C(n_367), .Y(n_363) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_187), .Y(n_178) );
BUFx3_ASAP7_75t_L g220 ( .A(n_179), .Y(n_220) );
INVx2_ASAP7_75t_L g253 ( .A(n_179), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_179), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g286 ( .A(n_179), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g319 ( .A(n_179), .Y(n_319) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_180), .A2(n_531), .B(n_535), .Y(n_530) );
INVx2_ASAP7_75t_SL g555 ( .A(n_180), .Y(n_555) );
INVx5_ASAP7_75t_L g222 ( .A(n_187), .Y(n_222) );
NOR2x1_ASAP7_75t_SL g271 ( .A(n_187), .B(n_261), .Y(n_271) );
BUFx2_ASAP7_75t_L g366 ( .A(n_187), .Y(n_366) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
INVxp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_208), .Y(n_196) );
NOR2xp33_ASAP7_75t_SL g264 ( .A(n_197), .B(n_265), .Y(n_264) );
NOR4xp25_ASAP7_75t_L g367 ( .A(n_197), .B(n_361), .C(n_365), .D(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g405 ( .A(n_197), .Y(n_405) );
AND2x2_ASAP7_75t_L g439 ( .A(n_197), .B(n_379), .Y(n_439) );
BUFx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g240 ( .A(n_198), .Y(n_240) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g294 ( .A(n_199), .Y(n_294) );
OAI21x1_ASAP7_75t_SL g199 ( .A1(n_200), .A2(n_202), .B(n_206), .Y(n_199) );
INVx1_ASAP7_75t_L g207 ( .A(n_201), .Y(n_207) );
AOI33xp33_ASAP7_75t_L g435 ( .A1(n_208), .A2(n_237), .A3(n_268), .B1(n_284), .B2(n_390), .B3(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g225 ( .A(n_209), .B(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g235 ( .A(n_209), .B(n_236), .Y(n_235) );
BUFx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g242 ( .A(n_210), .Y(n_242) );
INVxp67_ASAP7_75t_L g323 ( .A(n_210), .Y(n_323) );
AND2x2_ASAP7_75t_L g379 ( .A(n_210), .B(n_244), .Y(n_379) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_217), .B(n_218), .Y(n_210) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_211), .A2(n_217), .B(n_218), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_216), .Y(n_211) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_217), .A2(n_245), .B(n_251), .Y(n_244) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_217), .A2(n_245), .B(n_251), .Y(n_280) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_217), .A2(n_567), .B(n_573), .Y(n_566) );
AO21x2_ASAP7_75t_L g604 ( .A1(n_217), .A2(n_567), .B(n_573), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_219), .A2(n_401), .B(n_402), .Y(n_400) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
AND2x2_ASAP7_75t_L g388 ( .A(n_220), .B(n_262), .Y(n_388) );
AND3x2_ASAP7_75t_L g390 ( .A(n_220), .B(n_274), .C(n_329), .Y(n_390) );
INVx3_ASAP7_75t_SL g342 ( .A(n_221), .Y(n_342) );
INVx4_ASAP7_75t_L g236 ( .A(n_222), .Y(n_236) );
AND2x2_ASAP7_75t_L g274 ( .A(n_222), .B(n_261), .Y(n_274) );
INVxp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
BUFx2_ASAP7_75t_L g268 ( .A(n_226), .Y(n_268) );
AND2x4_ASAP7_75t_L g293 ( .A(n_226), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g356 ( .A(n_226), .B(n_244), .Y(n_356) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g326 ( .A(n_227), .Y(n_326) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_227), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_R g233 ( .A1(n_234), .A2(n_237), .B(n_241), .C(n_252), .Y(n_233) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g285 ( .A(n_236), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_236), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_236), .B(n_253), .Y(n_414) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g396 ( .A(n_238), .B(n_386), .Y(n_396) );
AND2x2_ASAP7_75t_SL g238 ( .A(n_239), .B(n_240), .Y(n_238) );
AND2x2_ASAP7_75t_L g243 ( .A(n_239), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g265 ( .A(n_239), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g281 ( .A(n_239), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g314 ( .A(n_239), .B(n_294), .Y(n_314) );
AND2x4_ASAP7_75t_L g279 ( .A(n_240), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g303 ( .A(n_240), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g341 ( .A(n_240), .B(n_266), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g269 ( .A(n_242), .B(n_266), .Y(n_269) );
AND2x2_ASAP7_75t_L g284 ( .A(n_242), .B(n_244), .Y(n_284) );
BUFx2_ASAP7_75t_L g340 ( .A(n_242), .Y(n_340) );
AND2x2_ASAP7_75t_L g354 ( .A(n_242), .B(n_265), .Y(n_354) );
INVx2_ASAP7_75t_L g266 ( .A(n_244), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_246), .B(n_250), .Y(n_245) );
OAI22xp33_ASAP7_75t_L g302 ( .A1(n_252), .A2(n_303), .B1(n_305), .B2(n_309), .Y(n_302) );
INVx2_ASAP7_75t_SL g333 ( .A(n_252), .Y(n_333) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_L g308 ( .A(n_253), .B(n_261), .Y(n_308) );
INVx1_ASAP7_75t_L g415 ( .A(n_254), .Y(n_415) );
NOR3xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_288), .C(n_302), .Y(n_255) );
OAI221xp5_ASAP7_75t_SL g256 ( .A1(n_257), .A2(n_263), .B1(n_267), .B2(n_270), .C(n_272), .Y(n_256) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g316 ( .A(n_260), .Y(n_316) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_260), .Y(n_444) );
INVx1_ASAP7_75t_L g407 ( .A(n_262), .Y(n_407) );
AND2x2_ASAP7_75t_SL g417 ( .A(n_262), .B(n_286), .Y(n_417) );
INVxp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_266), .B(n_294), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OR2x2_ASAP7_75t_L g300 ( .A(n_268), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g378 ( .A(n_268), .Y(n_378) );
AND2x2_ASAP7_75t_L g313 ( .A(n_269), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g359 ( .A(n_271), .B(n_319), .Y(n_359) );
AND2x2_ASAP7_75t_L g436 ( .A(n_271), .B(n_434), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_277), .B1(n_284), .B2(n_285), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g295 ( .A(n_276), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx2_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
AND2x4_ASAP7_75t_L g325 ( .A(n_279), .B(n_326), .Y(n_325) );
OAI21xp33_ASAP7_75t_SL g355 ( .A1(n_279), .A2(n_356), .B(n_357), .Y(n_355) );
AND2x2_ASAP7_75t_L g382 ( .A(n_279), .B(n_340), .Y(n_382) );
INVx2_ASAP7_75t_L g304 ( .A(n_280), .Y(n_304) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_280), .Y(n_337) );
INVx1_ASAP7_75t_SL g361 ( .A(n_281), .Y(n_361) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g292 ( .A(n_283), .Y(n_292) );
AND2x4_ASAP7_75t_SL g386 ( .A(n_283), .B(n_304), .Y(n_386) );
AND2x2_ASAP7_75t_L g383 ( .A(n_286), .B(n_329), .Y(n_383) );
AND2x2_ASAP7_75t_L g409 ( .A(n_286), .B(n_395), .Y(n_409) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_287), .Y(n_331) );
INVx1_ASAP7_75t_L g351 ( .A(n_287), .Y(n_351) );
OAI22xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_295), .B1(n_298), .B2(n_300), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_293), .B(n_304), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_293), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g432 ( .A(n_293), .Y(n_432) );
INVx2_ASAP7_75t_SL g357 ( .A(n_295), .Y(n_357) );
AND2x2_ASAP7_75t_L g369 ( .A(n_297), .B(n_329), .Y(n_369) );
INVx2_ASAP7_75t_L g375 ( .A(n_297), .Y(n_375) );
INVxp33_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g334 ( .A(n_300), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_303), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g425 ( .A(n_303), .Y(n_425) );
INVx1_ASAP7_75t_L g353 ( .A(n_305), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_306), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g364 ( .A(n_308), .B(n_365), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_308), .A2(n_438), .B1(n_439), .B2(n_440), .Y(n_437) );
NOR3xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_332), .C(n_335), .Y(n_310) );
OAI221xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B1(n_317), .B2(n_321), .C(n_324), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g430 ( .A(n_315), .Y(n_430) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g399 ( .A(n_316), .B(n_365), .Y(n_399) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g330 ( .A(n_319), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g401 ( .A(n_321), .Y(n_401) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g398 ( .A(n_322), .Y(n_398) );
INVx1_ASAP7_75t_L g404 ( .A(n_323), .Y(n_404) );
OR2x2_ASAP7_75t_L g427 ( .A(n_323), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_SL g336 ( .A(n_326), .Y(n_336) );
AND2x2_ASAP7_75t_L g406 ( .A(n_326), .B(n_386), .Y(n_406) );
AND2x2_ASAP7_75t_SL g438 ( .A(n_326), .B(n_339), .Y(n_438) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g443 ( .A(n_329), .Y(n_443) );
INVx1_ASAP7_75t_L g393 ( .A(n_331), .Y(n_393) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B(n_338), .C(n_342), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_336), .B(n_386), .Y(n_410) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_339), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AND2x2_ASAP7_75t_L g347 ( .A(n_341), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g428 ( .A(n_341), .Y(n_428) );
NAND4xp75_ASAP7_75t_L g343 ( .A(n_344), .B(n_400), .C(n_416), .D(n_437), .Y(n_343) );
NOR3x1_ASAP7_75t_L g344 ( .A(n_345), .B(n_362), .C(n_384), .Y(n_344) );
NAND4xp75_ASAP7_75t_L g345 ( .A(n_346), .B(n_352), .C(n_355), .D(n_358), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_347), .B(n_349), .Y(n_346) );
AND2x2_ASAP7_75t_L g397 ( .A(n_348), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g422 ( .A(n_349), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_SL g411 ( .A(n_354), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_370), .Y(n_362) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_366), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_376), .B(n_380), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI322xp33_ASAP7_75t_L g402 ( .A1(n_374), .A2(n_403), .A3(n_407), .B1(n_408), .B2(n_410), .C1(n_411), .C2(n_412), .Y(n_402) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_375), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_378), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_379), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B(n_389), .C(n_391), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_396), .B1(n_397), .B2(n_399), .Y(n_391) );
NOR2xp33_ASAP7_75t_SL g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B(n_406), .Y(n_403) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_409), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_413), .B(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g419 ( .A(n_414), .B(n_420), .Y(n_419) );
O2A1O1Ixp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B(n_423), .C(n_426), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI221xp5_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_429), .B1(n_431), .B2(n_433), .C(n_435), .Y(n_426) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g457 ( .A(n_449), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
AND2x6_ASAP7_75t_SL g473 ( .A(n_450), .B(n_452), .Y(n_473) );
OR2x6_ASAP7_75t_SL g476 ( .A(n_450), .B(n_451), .Y(n_476) );
OR2x2_ASAP7_75t_L g815 ( .A(n_450), .B(n_452), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_455), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
CKINVDCx11_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
CKINVDCx8_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_463), .B(n_816), .Y(n_462) );
INVx1_ASAP7_75t_L g817 ( .A(n_464), .Y(n_817) );
CKINVDCx6p67_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
INVx4_ASAP7_75t_SL g820 ( .A(n_471), .Y(n_820) );
INVx3_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
CKINVDCx11_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
OAI22x1_ASAP7_75t_L g818 ( .A1(n_476), .A2(n_819), .B1(n_820), .B2(n_821), .Y(n_818) );
INVx1_ASAP7_75t_L g821 ( .A(n_477), .Y(n_821) );
OR3x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_679), .C(n_750), .Y(n_477) );
NAND3x1_ASAP7_75t_SL g478 ( .A(n_479), .B(n_606), .C(n_628), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_596), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_527), .B1(n_574), .B2(n_578), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_481), .A2(n_782), .B1(n_783), .B2(n_785), .Y(n_781) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_502), .Y(n_481) );
AND2x2_ASAP7_75t_L g597 ( .A(n_482), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_482), .B(n_644), .Y(n_663) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g581 ( .A(n_483), .Y(n_581) );
AND2x2_ASAP7_75t_L g631 ( .A(n_483), .B(n_504), .Y(n_631) );
INVx1_ASAP7_75t_L g670 ( .A(n_483), .Y(n_670) );
OR2x2_ASAP7_75t_L g707 ( .A(n_483), .B(n_519), .Y(n_707) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_483), .Y(n_719) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_483), .Y(n_743) );
AND2x2_ASAP7_75t_L g800 ( .A(n_483), .B(n_627), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_491), .Y(n_484) );
INVx1_ASAP7_75t_L g551 ( .A(n_486), .Y(n_551) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g587 ( .A(n_487), .Y(n_587) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
OR2x6_ASAP7_75t_L g499 ( .A(n_488), .B(n_496), .Y(n_499) );
INVxp33_ASAP7_75t_L g561 ( .A(n_488), .Y(n_561) );
INVx1_ASAP7_75t_L g588 ( .A(n_490), .Y(n_588) );
INVxp67_ASAP7_75t_L g549 ( .A(n_492), .Y(n_549) );
NOR2x1p5_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g562 ( .A(n_495), .Y(n_562) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_499), .A2(n_508), .B1(n_509), .B2(n_510), .Y(n_507) );
INVxp67_ASAP7_75t_L g540 ( .A(n_499), .Y(n_540) );
INVx2_ASAP7_75t_L g594 ( .A(n_499), .Y(n_594) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_517), .Y(n_502) );
INVx1_ASAP7_75t_L g675 ( .A(n_503), .Y(n_675) );
AND2x2_ASAP7_75t_L g701 ( .A(n_503), .B(n_519), .Y(n_701) );
NAND2x1_ASAP7_75t_L g717 ( .A(n_503), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g598 ( .A(n_504), .B(n_584), .Y(n_598) );
INVx3_ASAP7_75t_L g627 ( .A(n_504), .Y(n_627) );
NOR2x1_ASAP7_75t_SL g746 ( .A(n_504), .B(n_519), .Y(n_746) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_511), .B(n_516), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_510), .B(n_542), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B1(n_514), .B2(n_515), .Y(n_511) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_517), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g625 ( .A(n_518), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g595 ( .A(n_519), .Y(n_595) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_519), .Y(n_640) );
AND2x2_ASAP7_75t_L g712 ( .A(n_519), .B(n_584), .Y(n_712) );
AND2x4_ASAP7_75t_L g729 ( .A(n_519), .B(n_673), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_519), .B(n_671), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_519), .B(n_580), .Y(n_805) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_527), .A2(n_622), .B1(n_693), .B2(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_552), .Y(n_527) );
INVx2_ASAP7_75t_L g695 ( .A(n_528), .Y(n_695) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_536), .Y(n_528) );
BUFx3_ASAP7_75t_L g685 ( .A(n_529), .Y(n_685) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_530), .B(n_554), .Y(n_577) );
INVx2_ASAP7_75t_L g601 ( .A(n_530), .Y(n_601) );
INVx1_ASAP7_75t_L g613 ( .A(n_530), .Y(n_613) );
AND2x4_ASAP7_75t_L g620 ( .A(n_530), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g637 ( .A(n_530), .B(n_537), .Y(n_637) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_530), .Y(n_651) );
INVxp67_ASAP7_75t_L g659 ( .A(n_530), .Y(n_659) );
AND2x2_ASAP7_75t_L g688 ( .A(n_536), .B(n_604), .Y(n_688) );
AND2x2_ASAP7_75t_L g704 ( .A(n_536), .B(n_605), .Y(n_704) );
NOR2xp67_ASAP7_75t_L g791 ( .A(n_536), .B(n_604), .Y(n_791) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g600 ( .A(n_537), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g611 ( .A(n_537), .Y(n_611) );
INVx1_ASAP7_75t_L g624 ( .A(n_537), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_537), .B(n_566), .Y(n_661) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_545), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_549), .B1(n_550), .B2(n_551), .Y(n_545) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g784 ( .A(n_552), .Y(n_784) );
AND2x4_ASAP7_75t_L g552 ( .A(n_553), .B(n_565), .Y(n_552) );
AND2x2_ASAP7_75t_L g658 ( .A(n_553), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g687 ( .A(n_553), .Y(n_687) );
AND2x2_ASAP7_75t_L g789 ( .A(n_553), .B(n_604), .Y(n_789) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_554), .B(n_566), .Y(n_649) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B(n_564), .Y(n_554) );
AO21x2_ASAP7_75t_L g605 ( .A1(n_555), .A2(n_556), .B(n_564), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_557), .B(n_563), .Y(n_556) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx3_ASAP7_75t_L g575 ( .A(n_565), .Y(n_575) );
NAND2x1p5_ASAP7_75t_L g764 ( .A(n_565), .B(n_685), .Y(n_764) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_566), .Y(n_678) );
AND2x2_ASAP7_75t_L g705 ( .A(n_566), .B(n_651), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AND2x2_ASAP7_75t_L g619 ( .A(n_575), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g635 ( .A(n_575), .Y(n_635) );
AND2x2_ASAP7_75t_L g723 ( .A(n_575), .B(n_600), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_575), .B(n_743), .Y(n_748) );
AND2x2_ASAP7_75t_L g758 ( .A(n_575), .B(n_637), .Y(n_758) );
OR2x2_ASAP7_75t_L g795 ( .A(n_575), .B(n_695), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_576), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g755 ( .A(n_576), .B(n_611), .Y(n_755) );
AND2x2_ASAP7_75t_L g771 ( .A(n_576), .B(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g765 ( .A(n_577), .B(n_661), .Y(n_765) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
INVx1_ASAP7_75t_L g647 ( .A(n_579), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_579), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g745 ( .A(n_579), .B(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_579), .B(n_626), .Y(n_770) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_580), .Y(n_617) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_581), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_582), .A2(n_615), .B1(n_633), .B2(n_636), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_582), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_SL g749 ( .A(n_582), .Y(n_749) );
AND2x4_ASAP7_75t_SL g582 ( .A(n_583), .B(n_595), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g626 ( .A(n_584), .B(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g646 ( .A(n_584), .Y(n_646) );
INVx1_ASAP7_75t_L g673 ( .A(n_584), .Y(n_673) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .Y(n_584) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .C(n_589), .Y(n_586) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_595), .Y(n_615) );
AND2x4_ASAP7_75t_L g672 ( .A(n_595), .B(n_673), .Y(n_672) );
NOR2x1_ASAP7_75t_L g733 ( .A(n_595), .B(n_702), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
AND2x2_ASAP7_75t_L g697 ( .A(n_597), .B(n_640), .Y(n_697) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_597), .A2(n_778), .B(n_779), .Y(n_777) );
INVx2_ASAP7_75t_L g655 ( .A(n_598), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_599), .A2(n_709), .B1(n_713), .B2(n_716), .Y(n_708) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_600), .Y(n_666) );
AND2x2_ASAP7_75t_L g676 ( .A(n_600), .B(n_677), .Y(n_676) );
INVx3_ASAP7_75t_L g715 ( .A(n_600), .Y(n_715) );
NAND2x1_ASAP7_75t_SL g740 ( .A(n_600), .B(n_609), .Y(n_740) );
AND2x2_ASAP7_75t_L g636 ( .A(n_602), .B(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NOR2x1_ASAP7_75t_L g612 ( .A(n_604), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g609 ( .A(n_605), .Y(n_609) );
INVx2_ASAP7_75t_L g621 ( .A(n_605), .Y(n_621) );
AOI21xp5_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_614), .B(n_618), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_609), .B(n_803), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_610), .A2(n_699), .B1(n_703), .B2(n_706), .Y(n_698) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
BUFx2_ASAP7_75t_L g803 ( .A(n_611), .Y(n_803) );
INVx1_ASAP7_75t_SL g810 ( .A(n_611), .Y(n_810) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_612), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OA21x2_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B(n_625), .Y(n_618) );
AND2x2_ASAP7_75t_L g622 ( .A(n_620), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g664 ( .A(n_620), .B(n_660), .Y(n_664) );
AND2x2_ASAP7_75t_L g779 ( .A(n_620), .B(n_677), .Y(n_779) );
AND2x2_ASAP7_75t_L g782 ( .A(n_620), .B(n_688), .Y(n_782) );
AND2x4_ASAP7_75t_L g790 ( .A(n_620), .B(n_791), .Y(n_790) );
OAI21xp33_ASAP7_75t_L g744 ( .A1(n_622), .A2(n_745), .B(n_747), .Y(n_744) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g772 ( .A(n_624), .Y(n_772) );
AND2x2_ASAP7_75t_L g788 ( .A(n_624), .B(n_789), .Y(n_788) );
INVx4_ASAP7_75t_L g702 ( .A(n_626), .Y(n_702) );
INVx1_ASAP7_75t_L g671 ( .A(n_627), .Y(n_671) );
AND2x2_ASAP7_75t_L g693 ( .A(n_627), .B(n_646), .Y(n_693) );
NOR2x1_ASAP7_75t_L g628 ( .A(n_629), .B(n_652), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B(n_638), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g639 ( .A(n_631), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_SL g792 ( .A(n_631), .B(n_644), .Y(n_792) );
AND2x2_ASAP7_75t_L g813 ( .A(n_631), .B(n_729), .Y(n_813) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g739 ( .A(n_636), .Y(n_739) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_641), .B(n_648), .Y(n_638) );
OR2x6_ASAP7_75t_L g691 ( .A(n_640), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_647), .Y(n_642) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
OR2x2_ASAP7_75t_L g714 ( .A(n_649), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g811 ( .A(n_649), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_650), .B(n_784), .Y(n_783) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_665), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_656), .B1(n_662), .B2(n_664), .Y(n_653) );
OR2x2_ASAP7_75t_L g725 ( .A(n_655), .B(n_726), .Y(n_725) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_657), .Y(n_682) );
NAND2x1p5_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVx1_ASAP7_75t_L g731 ( .A(n_660), .Y(n_731) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_674), .B2(n_676), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_672), .Y(n_668) );
AND2x4_ASAP7_75t_SL g669 ( .A(n_670), .B(n_671), .Y(n_669) );
AND2x2_ASAP7_75t_L g674 ( .A(n_672), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g735 ( .A(n_675), .B(n_729), .Y(n_735) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_680), .B(n_720), .Y(n_679) );
NOR2xp67_ASAP7_75t_L g680 ( .A(n_681), .B(n_694), .Y(n_680) );
AOI21xp33_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_683), .B(n_689), .Y(n_681) );
OR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
INVx3_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2x1p5_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI22xp33_ASAP7_75t_SL g759 ( .A1(n_691), .A2(n_760), .B1(n_762), .B2(n_765), .Y(n_759) );
NOR2x1_ASAP7_75t_L g706 ( .A(n_692), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g742 ( .A(n_693), .B(n_743), .Y(n_742) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B(n_698), .C(n_708), .Y(n_694) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp33_ASAP7_75t_SL g699 ( .A(n_700), .B(n_702), .Y(n_699) );
INVxp33_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g711 ( .A(n_702), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_703), .A2(n_723), .B1(n_724), .B2(n_727), .C(n_730), .Y(n_722) );
AND2x4_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g763 ( .A(n_704), .Y(n_763) );
INVx2_ASAP7_75t_SL g761 ( .A(n_707), .Y(n_761) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
NAND2x1_ASAP7_75t_L g760 ( .A(n_711), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g757 ( .A(n_717), .Y(n_757) );
INVx1_ASAP7_75t_L g786 ( .A(n_718), .Y(n_786) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NOR2x1_ASAP7_75t_L g720 ( .A(n_721), .B(n_736), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_734), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g775 ( .A(n_726), .Y(n_775) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g796 ( .A(n_729), .B(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g801 ( .A(n_729), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVxp33_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g754 ( .A(n_733), .Y(n_754) );
OAI21xp5_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_741), .B(n_744), .Y(n_736) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
BUFx2_ASAP7_75t_L g797 ( .A(n_743), .Y(n_797) );
AND2x2_ASAP7_75t_L g785 ( .A(n_746), .B(n_786), .Y(n_785) );
NOR2xp33_ASAP7_75t_R g747 ( .A(n_748), .B(n_749), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_766), .C(n_793), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_759), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_753), .B(n_756), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
OR2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_780), .Y(n_766) );
NAND2xp5_ASAP7_75t_SL g767 ( .A(n_768), .B(n_777), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_769), .A2(n_771), .B1(n_773), .B2(n_774), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NOR2x1_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVxp67_ASAP7_75t_SL g778 ( .A(n_776), .Y(n_778) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_781), .B(n_787), .Y(n_780) );
OAI21xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_790), .B(n_792), .Y(n_787) );
INVx1_ASAP7_75t_L g806 ( .A(n_790), .Y(n_806) );
AOI211xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_796), .B(n_798), .C(n_807), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_802), .B1(n_804), .B2(n_806), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_812), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVxp67_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
endmodule