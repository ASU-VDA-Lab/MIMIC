module fake_jpeg_21401_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_40),
.Y(n_48)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_44),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_25),
.B(n_23),
.C(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_48),
.Y(n_78)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_20),
.B1(n_16),
.B2(n_21),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_16),
.B1(n_20),
.B2(n_19),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_36),
.B1(n_44),
.B2(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_20),
.B1(n_19),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_65),
.A2(n_35),
.B1(n_17),
.B2(n_28),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_69),
.A2(n_47),
.B1(n_37),
.B2(n_21),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_75),
.A2(n_97),
.B1(n_32),
.B2(n_42),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_76),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_79),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_47),
.B1(n_37),
.B2(n_30),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_51),
.B(n_25),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_54),
.B(n_44),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_31),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_92),
.A2(n_100),
.B(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_18),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_18),
.Y(n_98)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_49),
.A2(n_68),
.B(n_30),
.C(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_49),
.B(n_28),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_56),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_110),
.B1(n_32),
.B2(n_42),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_31),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_18),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_18),
.Y(n_107)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_18),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_17),
.B(n_27),
.Y(n_117)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_24),
.B1(n_27),
.B2(n_41),
.Y(n_116)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx2_ASAP7_75t_SL g113 ( 
.A(n_111),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_87),
.B(n_104),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_99),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_117),
.A2(n_86),
.B1(n_96),
.B2(n_94),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_78),
.B(n_32),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_97),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_122),
.A2(n_136),
.B1(n_83),
.B2(n_82),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_96),
.B1(n_94),
.B2(n_90),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_139),
.B(n_104),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_32),
.B1(n_29),
.B2(n_13),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_77),
.A2(n_29),
.B(n_31),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_143),
.B(n_147),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_149),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_158),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_73),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_92),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_148),
.B(n_160),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_92),
.C(n_103),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_151),
.C(n_126),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_73),
.C(n_84),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_74),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_152),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_100),
.B1(n_84),
.B2(n_106),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_154),
.B1(n_165),
.B2(n_115),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_110),
.B1(n_88),
.B2(n_102),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_80),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_167),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_29),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_120),
.B(n_80),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_125),
.B1(n_113),
.B2(n_132),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_163),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_120),
.B(n_80),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_88),
.B1(n_42),
.B2(n_45),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_170),
.B1(n_115),
.B2(n_121),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_45),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_90),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_172),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_45),
.B1(n_111),
.B2(n_33),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_114),
.B(n_29),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_82),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_184),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_116),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_188),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_135),
.C(n_130),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_186),
.A2(n_146),
.B1(n_29),
.B2(n_34),
.Y(n_224)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_157),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_156),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_167),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_172),
.B1(n_165),
.B2(n_137),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_116),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_116),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_116),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_33),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_146),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_201),
.B(n_132),
.Y(n_211)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_135),
.B1(n_126),
.B2(n_139),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_162),
.B1(n_153),
.B2(n_121),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_205),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_158),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_209),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_194),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_210),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_142),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_220),
.B1(n_227),
.B2(n_197),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_151),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_204),
.C(n_184),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_219),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_137),
.B1(n_132),
.B2(n_117),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_221),
.A2(n_224),
.B1(n_189),
.B2(n_198),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_180),
.A2(n_33),
.B(n_26),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_226),
.Y(n_236)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

NOR2x1_ASAP7_75t_R g228 ( 
.A(n_200),
.B(n_26),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_221),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_174),
.B(n_26),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_175),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_26),
.Y(n_230)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_1),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_182),
.B1(n_181),
.B2(n_199),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_179),
.B(n_1),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_239),
.A2(n_227),
.B1(n_230),
.B2(n_220),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_248),
.C(n_249),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_243),
.B1(n_253),
.B2(n_258),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_229),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_235),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_246),
.B(n_257),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_175),
.C(n_177),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_195),
.C(n_180),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_215),
.A2(n_191),
.B1(n_181),
.B2(n_182),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_193),
.C(n_178),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_201),
.C(n_190),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_222),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_215),
.A2(n_187),
.B1(n_192),
.B2(n_202),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_244),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_261),
.B(n_236),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_214),
.C(n_207),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_275),
.C(n_276),
.Y(n_283)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_234),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_271),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_218),
.B(n_228),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_274),
.B1(n_255),
.B2(n_241),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_245),
.B(n_206),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_247),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_231),
.B1(n_206),
.B2(n_213),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_213),
.C(n_232),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_248),
.C(n_256),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_225),
.C(n_224),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_278),
.C(n_242),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_237),
.B(n_236),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_284),
.B(n_290),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_251),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_293),
.B1(n_268),
.B2(n_264),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_288),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_238),
.C(n_176),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_291),
.C(n_294),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_262),
.A2(n_176),
.B(n_226),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_7),
.C(n_14),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_5),
.C(n_11),
.Y(n_294)
);

FAx1_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_268),
.CI(n_271),
.CON(n_296),
.SN(n_296)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_304),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_275),
.C(n_261),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_303),
.C(n_308),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_270),
.Y(n_301)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_259),
.C(n_6),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_5),
.C(n_11),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_5),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_306),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_292),
.B(n_10),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_11),
.C(n_15),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_308),
.B(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_310),
.B(n_318),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_280),
.B(n_287),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_297),
.Y(n_324)
);

INVx11_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_303),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_296),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_15),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_314),
.A2(n_298),
.B(n_311),
.Y(n_320)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_321),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_307),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_324),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_297),
.C(n_307),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_318),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_322),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_331),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_319),
.B(n_316),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_328),
.C(n_326),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_329),
.B(n_309),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_315),
.Y(n_336)
);


endmodule