module fake_jpeg_12102_n_585 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_585);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_585;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_60),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_63),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_62),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_65),
.Y(n_128)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_70),
.Y(n_170)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_72),
.B(n_120),
.Y(n_154)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_74),
.B(n_85),
.Y(n_132)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_77),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_78),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_79),
.Y(n_200)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_82),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_83),
.Y(n_209)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_84),
.Y(n_191)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_27),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_87),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_29),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

BUFx24_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

CKINVDCx6p67_ASAP7_75t_R g161 ( 
.A(n_89),
.Y(n_161)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_90),
.Y(n_194)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_91),
.Y(n_193)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_27),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_95),
.B(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_27),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_103),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_29),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_104),
.Y(n_210)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_105),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_29),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_119),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_25),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_115),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_19),
.B(n_15),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_125),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_28),
.B(n_1),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_117),
.B(n_118),
.Y(n_199)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_28),
.Y(n_118)
);

INVx2_ASAP7_75t_R g119 ( 
.A(n_29),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_39),
.B(n_52),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_30),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_122),
.B(n_124),
.Y(n_206)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_41),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_40),
.Y(n_176)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_39),
.B(n_15),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_52),
.B(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_126),
.B(n_4),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_41),
.B1(n_55),
.B2(n_53),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_130),
.A2(n_143),
.B1(n_151),
.B2(n_165),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_45),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_135),
.B(n_176),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_63),
.A2(n_50),
.B1(n_46),
.B2(n_42),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_142),
.A2(n_180),
.B1(n_128),
.B2(n_127),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_34),
.B1(n_54),
.B2(n_37),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_60),
.A2(n_55),
.B1(n_41),
.B2(n_46),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_145),
.A2(n_148),
.B1(n_150),
.B2(n_157),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_60),
.A2(n_55),
.B1(n_46),
.B2(n_42),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_82),
.A2(n_50),
.B1(n_26),
.B2(n_45),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_106),
.A2(n_40),
.B1(n_56),
.B2(n_38),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_82),
.A2(n_50),
.B1(n_26),
.B2(n_45),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_112),
.A2(n_45),
.B1(n_53),
.B2(n_49),
.Y(n_158)
);

AO22x1_ASAP7_75t_L g214 ( 
.A1(n_158),
.A2(n_187),
.B1(n_189),
.B2(n_9),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_117),
.A2(n_23),
.B1(n_54),
.B2(n_37),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_89),
.A2(n_45),
.B1(n_49),
.B2(n_48),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_166),
.A2(n_168),
.B1(n_195),
.B2(n_78),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_84),
.B(n_34),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_167),
.B(n_188),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_89),
.A2(n_38),
.B1(n_56),
.B2(n_48),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_97),
.B(n_58),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_174),
.B(n_196),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_109),
.A2(n_58),
.B1(n_32),
.B2(n_24),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_90),
.B(n_2),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_9),
.Y(n_219)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_92),
.Y(n_183)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_73),
.A2(n_32),
.B1(n_24),
.B2(n_23),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_110),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_97),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_59),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_77),
.B(n_4),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_205),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_88),
.B(n_7),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_70),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_113),
.B(n_121),
.Y(n_205)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_93),
.B(n_8),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_212),
.Y(n_236)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_123),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_211),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_99),
.B(n_8),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_136),
.B(n_9),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_213),
.B(n_216),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_214),
.A2(n_245),
.B(n_262),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_169),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_135),
.B(n_9),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_218),
.B(n_226),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_219),
.B(n_231),
.Y(n_310)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_220),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_221),
.Y(n_315)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_222),
.Y(n_288)
);

BUFx8_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_223),
.Y(n_331)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_225),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_155),
.B(n_10),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_151),
.A2(n_79),
.B1(n_101),
.B2(n_100),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_227),
.A2(n_209),
.B1(n_170),
.B2(n_198),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_133),
.B(n_67),
.C(n_98),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_228),
.B(n_249),
.C(n_260),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_230),
.B(n_242),
.Y(n_293)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_130),
.A2(n_83),
.B1(n_104),
.B2(n_12),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_233),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_191),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_238),
.Y(n_287)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_235),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_129),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_244),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_131),
.B(n_10),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_129),
.Y(n_244)
);

OR2x4_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_14),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_145),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_247),
.B(n_254),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_140),
.Y(n_248)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_11),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_176),
.B(n_11),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_250),
.B(n_255),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_154),
.B(n_11),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_251),
.B(n_269),
.Y(n_314)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_138),
.Y(n_252)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_252),
.Y(n_320)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_253),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_186),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_141),
.B(n_11),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_144),
.B(n_12),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_256),
.B(n_261),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_211),
.A2(n_127),
.B1(n_207),
.B2(n_172),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_257),
.Y(n_297)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_177),
.Y(n_258)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_140),
.Y(n_259)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_259),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_156),
.B(n_152),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_168),
.B(n_173),
.Y(n_261)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_204),
.Y(n_263)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_137),
.B(n_173),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_264),
.B(n_267),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_184),
.B(n_183),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_282),
.C(n_163),
.Y(n_318)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_139),
.Y(n_266)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_266),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_137),
.B(n_166),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_153),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_284),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_161),
.B(n_193),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_161),
.A2(n_148),
.B(n_150),
.C(n_157),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_270),
.B(n_279),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_149),
.A2(n_160),
.B1(n_159),
.B2(n_190),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_271),
.A2(n_273),
.B1(n_278),
.B2(n_285),
.Y(n_336)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_170),
.Y(n_272)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_149),
.A2(n_160),
.B1(n_159),
.B2(n_190),
.Y(n_273)
);

OR2x2_ASAP7_75t_SL g275 ( 
.A(n_147),
.B(n_172),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_163),
.C(n_146),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_193),
.B(n_139),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_276),
.B(n_283),
.Y(n_324)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_153),
.Y(n_277)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_171),
.A2(n_210),
.B1(n_192),
.B2(n_200),
.Y(n_278)
);

AO22x1_ASAP7_75t_SL g279 ( 
.A1(n_195),
.A2(n_179),
.B1(n_210),
.B2(n_192),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_178),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_186),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_128),
.B(n_179),
.C(n_185),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_147),
.B(n_146),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_185),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_171),
.B(n_200),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_285),
.B(n_231),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_260),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_295),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_260),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_296),
.A2(n_341),
.B(n_268),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_265),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_303),
.B(n_298),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_304),
.A2(n_308),
.B1(n_329),
.B2(n_331),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_229),
.A2(n_198),
.B1(n_209),
.B2(n_178),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_308),
.A2(n_329),
.B1(n_332),
.B2(n_304),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_274),
.B(n_163),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_316),
.B(n_321),
.Y(n_364)
);

INVx8_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_317),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_223),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_216),
.B(n_134),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_319),
.B(n_322),
.C(n_340),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_249),
.B(n_134),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_217),
.B(n_244),
.C(n_228),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_237),
.A2(n_227),
.B1(n_247),
.B2(n_261),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_237),
.A2(n_231),
.B1(n_217),
.B2(n_265),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_226),
.B(n_236),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_333),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_336),
.A2(n_315),
.B1(n_335),
.B2(n_289),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_230),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_217),
.B(n_213),
.C(n_218),
.Y(n_340)
);

AOI32xp33_ASAP7_75t_L g341 ( 
.A1(n_267),
.A2(n_250),
.A3(n_264),
.B1(n_255),
.B2(n_256),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_343),
.B(n_344),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_219),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_287),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_345),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_338),
.A2(n_231),
.B1(n_219),
.B2(n_282),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_346),
.A2(n_349),
.B1(n_354),
.B2(n_358),
.Y(n_396)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_309),
.Y(n_347)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_347),
.Y(n_398)
);

OAI32xp33_ASAP7_75t_L g348 ( 
.A1(n_328),
.A2(n_232),
.A3(n_270),
.B1(n_214),
.B2(n_275),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_348),
.B(n_351),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_310),
.A2(n_279),
.B1(n_215),
.B2(n_284),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_335),
.A2(n_280),
.B(n_279),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_350),
.A2(n_355),
.B(n_375),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_239),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_352),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_362),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_296),
.A2(n_223),
.B(n_245),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_239),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_356),
.B(n_363),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_310),
.A2(n_272),
.B1(n_259),
.B2(n_240),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_325),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_366),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_305),
.B(n_263),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_361),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_312),
.B(n_290),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_310),
.A2(n_258),
.B1(n_280),
.B2(n_246),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_365),
.A2(n_326),
.B1(n_327),
.B2(n_337),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_325),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_324),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_367),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_312),
.B(n_246),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_372),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_301),
.A2(n_277),
.B(n_253),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_371),
.A2(n_379),
.B(n_380),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_290),
.B(n_292),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_373),
.A2(n_381),
.B1(n_382),
.B2(n_299),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_330),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_374),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_305),
.B(n_319),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_376),
.B(n_378),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_325),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_377),
.A2(n_384),
.B(n_359),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_292),
.B(n_293),
.Y(n_378)
);

INVx2_ASAP7_75t_R g379 ( 
.A(n_309),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_315),
.A2(n_322),
.B(n_314),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_318),
.A2(n_297),
.B1(n_340),
.B2(n_311),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_302),
.Y(n_383)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_383),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_331),
.A2(n_339),
.B(n_326),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_351),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_387),
.B(n_412),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_370),
.B(n_311),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_391),
.B(n_372),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_375),
.A2(n_306),
.B(n_320),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_395),
.A2(n_417),
.B(n_355),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_397),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_299),
.C(n_320),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_418),
.C(n_353),
.Y(n_434)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_401),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_373),
.A2(n_336),
.B1(n_339),
.B2(n_330),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_402),
.A2(n_414),
.B(n_384),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_403),
.A2(n_406),
.B1(n_409),
.B2(n_291),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_404),
.A2(n_349),
.B1(n_343),
.B2(n_361),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_354),
.A2(n_323),
.B1(n_337),
.B2(n_306),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_346),
.A2(n_323),
.B1(n_307),
.B2(n_288),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_383),
.Y(n_410)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_410),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_368),
.B(n_288),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_381),
.A2(n_291),
.B1(n_300),
.B2(n_307),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_376),
.Y(n_415)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_356),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_345),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_375),
.A2(n_355),
.B(n_361),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_300),
.C(n_327),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_420),
.A2(n_429),
.B1(n_396),
.B2(n_409),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_342),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_421),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_363),
.Y(n_422)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_422),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_423),
.A2(n_435),
.B(n_448),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_425),
.B(n_393),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_394),
.B(n_342),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_426),
.Y(n_475)
);

A2O1A1O1Ixp25_ASAP7_75t_L g427 ( 
.A1(n_417),
.A2(n_362),
.B(n_380),
.C(n_378),
.D(n_344),
.Y(n_427)
);

NOR3xp33_ASAP7_75t_L g470 ( 
.A(n_427),
.B(n_431),
.C(n_395),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_382),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_434),
.C(n_439),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_404),
.A2(n_350),
.B1(n_369),
.B2(n_358),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_412),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_445),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_437),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_413),
.A2(n_353),
.B(n_377),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_436),
.Y(n_463)
);

OAI32xp33_ASAP7_75t_L g437 ( 
.A1(n_399),
.A2(n_364),
.A3(n_348),
.B1(n_366),
.B2(n_365),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_389),
.B(n_353),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_392),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_389),
.B(n_357),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_447),
.C(n_450),
.Y(n_467)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_443),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_394),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_419),
.Y(n_446)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_446),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_400),
.B(n_371),
.C(n_364),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_413),
.A2(n_379),
.B(n_347),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_411),
.B(n_286),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_398),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_451),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_453),
.A2(n_457),
.B1(n_405),
.B2(n_433),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_429),
.A2(n_396),
.B1(n_406),
.B2(n_386),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_454),
.A2(n_461),
.B1(n_443),
.B2(n_449),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_420),
.A2(n_386),
.B1(n_399),
.B2(n_407),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_407),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_459),
.B(n_469),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_448),
.A2(n_386),
.B1(n_416),
.B2(n_387),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_428),
.B(n_418),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_471),
.C(n_477),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_286),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_470),
.B(n_478),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_434),
.B(n_411),
.C(n_413),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_424),
.B(n_408),
.Y(n_473)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_473),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_426),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_421),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_425),
.B(n_393),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_426),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_422),
.B(n_405),
.Y(n_479)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_479),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_480),
.B(n_439),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_442),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_481),
.B(n_493),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_483),
.B(n_452),
.Y(n_509)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_484),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_456),
.Y(n_486)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_486),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_487),
.A2(n_455),
.B1(n_461),
.B2(n_403),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_462),
.A2(n_449),
.B(n_458),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_488),
.A2(n_472),
.B(n_427),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_452),
.B(n_447),
.C(n_435),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_467),
.C(n_477),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_438),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_495),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_462),
.A2(n_421),
.B(n_423),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_491),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_390),
.Y(n_493)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_476),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_497),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_473),
.B(n_405),
.Y(n_497)
);

CKINVDCx14_ASAP7_75t_R g498 ( 
.A(n_479),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_498),
.A2(n_502),
.B1(n_503),
.B2(n_401),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_467),
.B(n_390),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_504),
.Y(n_512)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_463),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_501),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_453),
.A2(n_402),
.B1(n_414),
.B2(n_437),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_436),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_465),
.B(n_430),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_505),
.B(n_457),
.Y(n_506)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_506),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_499),
.A2(n_472),
.B1(n_465),
.B2(n_454),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_508),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_509),
.B(n_519),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_515),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_513),
.B(n_516),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_514),
.A2(n_522),
.B1(n_523),
.B2(n_501),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_482),
.B(n_480),
.C(n_455),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_482),
.B(n_468),
.C(n_463),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_481),
.B(n_468),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_489),
.B(n_440),
.C(n_410),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_488),
.C(n_491),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_487),
.A2(n_502),
.B1(n_494),
.B2(n_504),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_507),
.A2(n_484),
.B1(n_494),
.B2(n_490),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_526),
.B(n_533),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_527),
.B(n_529),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_500),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_SL g530 ( 
.A(n_520),
.B(n_492),
.Y(n_530)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_530),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_485),
.Y(n_532)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_532),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_519),
.B(n_493),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_534),
.A2(n_538),
.B1(n_525),
.B2(n_388),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_513),
.B(n_483),
.C(n_495),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_535),
.B(n_524),
.C(n_515),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_507),
.A2(n_496),
.B(n_388),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_536),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_518),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_541),
.B(n_528),
.C(n_526),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_531),
.B(n_512),
.C(n_524),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_543),
.B(n_544),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_527),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_540),
.A2(n_517),
.B1(n_511),
.B2(n_523),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_549),
.B(n_550),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_537),
.A2(n_525),
.B1(n_510),
.B2(n_512),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_529),
.B(n_509),
.C(n_514),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_551),
.B(n_553),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_552),
.B(n_441),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_540),
.A2(n_460),
.B1(n_464),
.B2(n_451),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_548),
.Y(n_554)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_554),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_542),
.A2(n_539),
.B(n_535),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_555),
.A2(n_547),
.B(n_392),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_545),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_557),
.B(n_558),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_546),
.B(n_533),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_561),
.B(n_562),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_541),
.C(n_551),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_563),
.B(n_564),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_546),
.B(n_528),
.C(n_460),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_563),
.B(n_464),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_565),
.B(n_571),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_556),
.B(n_549),
.Y(n_566)
);

AO21x1_ASAP7_75t_L g577 ( 
.A1(n_566),
.A2(n_570),
.B(n_398),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_569),
.A2(n_562),
.B(n_564),
.Y(n_575)
);

AOI21xp33_ASAP7_75t_L g570 ( 
.A1(n_560),
.A2(n_547),
.B(n_392),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_568),
.B(n_554),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_573),
.B(n_574),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_575),
.B(n_576),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_567),
.B(n_559),
.C(n_558),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_577),
.B(n_572),
.C(n_571),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_579),
.A2(n_580),
.B(n_578),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_581),
.A2(n_582),
.B(n_379),
.Y(n_583)
);

OAI211xp5_ASAP7_75t_SL g582 ( 
.A1(n_578),
.A2(n_379),
.B(n_360),
.C(n_374),
.Y(n_582)
);

OAI221xp5_ASAP7_75t_SL g584 ( 
.A1(n_583),
.A2(n_360),
.B1(n_374),
.B2(n_294),
.C(n_317),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_584),
.B(n_360),
.Y(n_585)
);


endmodule