module fake_jpeg_19672_n_163 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_163);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_34),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_37),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_20),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_44),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_23),
.B1(n_30),
.B2(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_53),
.B1(n_67),
.B2(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_60),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_23),
.B1(n_30),
.B2(n_21),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_16),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_1),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_15),
.B(n_25),
.C(n_16),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_34),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_65),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_17),
.B1(n_28),
.B2(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_17),
.B1(n_28),
.B2(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_86),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_75),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_38),
.B1(n_29),
.B2(n_28),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_93),
.B1(n_48),
.B2(n_46),
.Y(n_99)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_65),
.B(n_62),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_54),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_14),
.B1(n_20),
.B2(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_13),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_101),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_49),
.B1(n_46),
.B2(n_48),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_103),
.B(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_108),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_75),
.B1(n_76),
.B2(n_86),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_85),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_73),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_50),
.Y(n_108)
);

OAI21x1_ASAP7_75t_R g110 ( 
.A1(n_92),
.A2(n_57),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_70),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_84),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_74),
.C(n_87),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_126),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_118),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_121),
.B(n_122),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_97),
.B1(n_111),
.B2(n_106),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_120),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_81),
.B(n_79),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_89),
.B1(n_82),
.B2(n_47),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVx2_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_98),
.B1(n_52),
.B2(n_87),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_71),
.B1(n_47),
.B2(n_50),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_106),
.B1(n_109),
.B2(n_103),
.Y(n_130)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_119),
.B1(n_124),
.B2(n_112),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_131),
.B1(n_57),
.B2(n_11),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_110),
.B1(n_100),
.B2(n_107),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_98),
.B(n_110),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_122),
.B(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_9),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_121),
.Y(n_138)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_146),
.B1(n_128),
.B2(n_137),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_145),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_141),
.Y(n_148)
);

AO221x1_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_77),
.B1(n_126),
.B2(n_57),
.C(n_113),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_134),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_144),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_127),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_129),
.B(n_135),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_146),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_134),
.C(n_140),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_149),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_138),
.B1(n_143),
.B2(n_139),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_153),
.B(n_156),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_155),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_149),
.Y(n_155)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_152),
.B(n_148),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_155),
.C(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_151),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_160),
.A2(n_161),
.B(n_159),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_158),
.Y(n_163)
);


endmodule