module fake_jpeg_12130_n_64 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_5),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_26),
.B1(n_14),
.B2(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_37),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_35),
.B1(n_38),
.B2(n_9),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_23),
.B1(n_18),
.B2(n_13),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2x1_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_14),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_31),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_44),
.C(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_0),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_29),
.B1(n_30),
.B2(n_9),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_36),
.B1(n_33),
.B2(n_11),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_50),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_3),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_45),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_51),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_48),
.C(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_7),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_55),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_53),
.B(n_56),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_7),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_61),
.B(n_8),
.Y(n_64)
);


endmodule