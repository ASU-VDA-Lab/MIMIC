module fake_netlist_1_6100_n_525 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_525);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_525;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_44), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_67), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_69), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_10), .Y(n_79) );
NOR2xp67_ASAP7_75t_L g80 ( .A(n_64), .B(n_28), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_65), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_17), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_22), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_6), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_18), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_71), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_0), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_5), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_50), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_70), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_60), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_63), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_11), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_36), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_57), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_13), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_12), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_52), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_49), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_48), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_38), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_30), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_2), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_1), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_5), .B(n_32), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_51), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_54), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_10), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_15), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_73), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_55), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_0), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_62), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_41), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_81), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_81), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_84), .A2(n_109), .B1(n_79), .B2(n_111), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_84), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_82), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_82), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_93), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_85), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_114), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_77), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_83), .B(n_3), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_97), .B(n_4), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_109), .B(n_4), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_94), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_97), .B(n_6), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_91), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_94), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_108), .B(n_7), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
BUFx3_ASAP7_75t_L g136 ( .A(n_131), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_121), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_121), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_131), .B(n_108), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_124), .B(n_78), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_121), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_121), .Y(n_142) );
INVx4_ASAP7_75t_SL g143 ( .A(n_131), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_117), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_121), .Y(n_146) );
BUFx4f_ASAP7_75t_L g147 ( .A(n_115), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_125), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_125), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_124), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_122), .B(n_87), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_126), .A2(n_103), .B1(n_96), .B2(n_104), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_115), .B(n_78), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_129), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_129), .Y(n_155) );
BUFx10_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_133), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_117), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_133), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_148), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_153), .B(n_126), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_156), .B(n_116), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_156), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_156), .B(n_119), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_156), .B(n_119), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_140), .B(n_120), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_147), .B(n_120), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_139), .A2(n_134), .B1(n_127), .B2(n_118), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_147), .B(n_123), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g172 ( .A1(n_147), .A2(n_135), .B(n_132), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_150), .B(n_86), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_136), .A2(n_135), .B(n_132), .Y(n_175) );
OAI22xp33_ASAP7_75t_L g176 ( .A1(n_145), .A2(n_128), .B1(n_130), .B2(n_123), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_151), .B(n_130), .Y(n_177) );
O2A1O1Ixp5_ASAP7_75t_L g178 ( .A1(n_150), .A2(n_134), .B(n_127), .C(n_89), .Y(n_178) );
AOI22x1_ASAP7_75t_L g179 ( .A1(n_137), .A2(n_114), .B1(n_95), .B2(n_99), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_158), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_151), .B(n_113), .Y(n_182) );
OR2x2_ASAP7_75t_L g183 ( .A(n_152), .B(n_112), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_150), .B(n_113), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_136), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_144), .B(n_86), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_152), .B(n_87), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_150), .B(n_90), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_144), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_143), .Y(n_190) );
NOR3xp33_ASAP7_75t_SL g191 ( .A(n_181), .B(n_90), .C(n_101), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_169), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
OR2x6_ASAP7_75t_L g194 ( .A(n_164), .B(n_144), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_189), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_173), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_177), .B(n_162), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_172), .B(n_143), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_163), .A2(n_139), .B(n_159), .Y(n_199) );
NOR2xp33_ASAP7_75t_R g200 ( .A(n_181), .B(n_101), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_163), .B(n_143), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_172), .B(n_143), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_164), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_182), .B(n_139), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_165), .A2(n_139), .B1(n_155), .B2(n_159), .Y(n_205) );
INVx4_ASAP7_75t_L g206 ( .A(n_164), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_173), .Y(n_207) );
AO32x1_ASAP7_75t_L g208 ( .A1(n_160), .A2(n_95), .A3(n_76), .B1(n_92), .B2(n_102), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_173), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_170), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_166), .B(n_155), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_178), .A2(n_149), .B(n_157), .C(n_154), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_175), .A2(n_149), .B(n_157), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_164), .B(n_107), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_176), .B(n_107), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
NAND2xp33_ASAP7_75t_SL g217 ( .A(n_164), .B(n_105), .Y(n_217) );
BUFx4f_ASAP7_75t_L g218 ( .A(n_185), .Y(n_218) );
INVx6_ASAP7_75t_L g219 ( .A(n_189), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_185), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_184), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_203), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_212), .A2(n_190), .B(n_180), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_216), .A2(n_197), .B(n_217), .C(n_199), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_201), .A2(n_184), .B(n_188), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_221), .B(n_170), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_217), .A2(n_183), .B1(n_186), .B2(n_187), .Y(n_227) );
NOR2x1_ASAP7_75t_SL g228 ( .A(n_194), .B(n_189), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_211), .A2(n_183), .B1(n_185), .B2(n_187), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_192), .A2(n_190), .B(n_180), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_204), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_196), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_210), .B(n_174), .Y(n_233) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_195), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_203), .Y(n_235) );
CKINVDCx12_ASAP7_75t_R g236 ( .A(n_194), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_193), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_205), .A2(n_179), .B1(n_105), .B2(n_88), .Y(n_238) );
BUFx8_ASAP7_75t_L g239 ( .A(n_207), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_200), .Y(n_240) );
AOI221x1_ASAP7_75t_L g241 ( .A1(n_213), .A2(n_98), .B1(n_100), .B2(n_110), .C(n_88), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_196), .A2(n_160), .B(n_161), .Y(n_242) );
NAND3xp33_ASAP7_75t_SL g243 ( .A(n_210), .B(n_106), .C(n_142), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_198), .A2(n_154), .B(n_148), .C(n_80), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_207), .A2(n_161), .B(n_168), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_215), .B(n_168), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_198), .B(n_168), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_237), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_224), .A2(n_194), .B(n_220), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_232), .Y(n_250) );
OAI211xp5_ASAP7_75t_SL g251 ( .A1(n_233), .A2(n_191), .B(n_214), .C(n_138), .Y(n_251) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_244), .A2(n_179), .B(n_138), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_242), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_224), .A2(n_194), .B(n_220), .Y(n_254) );
OR2x6_ASAP7_75t_L g255 ( .A(n_222), .B(n_206), .Y(n_255) );
HB1xp67_ASAP7_75t_SL g256 ( .A(n_240), .Y(n_256) );
NAND3xp33_ASAP7_75t_L g257 ( .A(n_244), .B(n_202), .C(n_203), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_239), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_243), .A2(n_202), .B1(n_219), .B2(n_218), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_246), .A2(n_209), .B(n_218), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_231), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_227), .B(n_209), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_229), .A2(n_142), .B(n_141), .C(n_137), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_236), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_226), .B(n_206), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_239), .B(n_206), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_222), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_245), .A2(n_141), .B(n_146), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_230), .Y(n_269) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_249), .A2(n_223), .B(n_225), .Y(n_270) );
OAI31xp33_ASAP7_75t_L g271 ( .A1(n_261), .A2(n_238), .A3(n_246), .B(n_234), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_255), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_250), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_255), .Y(n_274) );
AND2x6_ASAP7_75t_L g275 ( .A(n_269), .B(n_247), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_261), .B(n_235), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_254), .A2(n_247), .B(n_218), .C(n_235), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g278 ( .A1(n_248), .A2(n_154), .B1(n_148), .B2(n_222), .C(n_146), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_250), .B(n_222), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_248), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_251), .A2(n_219), .B1(n_154), .B2(n_148), .Y(n_281) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_257), .A2(n_208), .B(n_228), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_269), .B(n_241), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g284 ( .A1(n_262), .A2(n_154), .B1(n_168), .B2(n_208), .C(n_11), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_265), .B(n_154), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_267), .B(n_7), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_267), .B(n_8), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_255), .B(n_8), .Y(n_288) );
OR2x6_ASAP7_75t_L g289 ( .A(n_255), .B(n_219), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_253), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_290), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_280), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_272), .B(n_257), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_280), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_273), .B(n_255), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_290), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_279), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_279), .B(n_252), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_290), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_273), .B(n_266), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_274), .B(n_264), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_276), .B(n_252), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_274), .B(n_252), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_272), .B(n_252), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_272), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_272), .B(n_260), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_270), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_270), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_288), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_283), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_283), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_288), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_270), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_289), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_282), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_289), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_298), .B(n_282), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_298), .B(n_282), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_303), .B(n_270), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_301), .B(n_271), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_303), .B(n_287), .Y(n_324) );
INVx5_ASAP7_75t_SL g325 ( .A(n_293), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_304), .B(n_287), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_301), .B(n_300), .Y(n_327) );
BUFx6f_ASAP7_75t_SL g328 ( .A(n_318), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_311), .B(n_285), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_304), .B(n_286), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_292), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_291), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_307), .B(n_286), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_300), .B(n_271), .Y(n_334) );
NOR2xp67_ASAP7_75t_L g335 ( .A(n_316), .B(n_285), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_292), .B(n_275), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_294), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_307), .B(n_275), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_294), .B(n_275), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_291), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_305), .B(n_275), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_291), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_305), .B(n_275), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_296), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_293), .B(n_275), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_295), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_310), .A2(n_275), .B1(n_259), .B2(n_289), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_311), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_313), .B(n_275), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_302), .B(n_277), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_312), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_296), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_312), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_318), .B(n_253), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_296), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_306), .B(n_260), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_302), .B(n_289), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_295), .Y(n_358) );
NOR2x1p5_ASAP7_75t_L g359 ( .A(n_318), .B(n_258), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_299), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_321), .B(n_293), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_331), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_337), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_337), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_322), .B(n_315), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_321), .B(n_293), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_346), .B(n_327), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_348), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_358), .B(n_317), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_324), .B(n_317), .Y(n_371) );
INVx2_ASAP7_75t_SL g372 ( .A(n_359), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_332), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_348), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_351), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_332), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_351), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_324), .B(n_316), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_319), .B(n_314), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_334), .B(n_323), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_329), .B(n_314), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_335), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_319), .B(n_314), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_353), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_320), .B(n_309), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_320), .B(n_309), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_332), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_329), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_355), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_357), .B(n_256), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_326), .B(n_309), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_350), .B(n_315), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_359), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g395 ( .A(n_335), .B(n_306), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_355), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_326), .B(n_308), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_333), .B(n_308), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_330), .B(n_299), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_330), .B(n_299), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_333), .B(n_289), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_341), .B(n_284), .Y(n_402) );
INVxp33_ASAP7_75t_L g403 ( .A(n_354), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_349), .Y(n_404) );
NAND2xp33_ASAP7_75t_SL g405 ( .A(n_328), .B(n_281), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_356), .B(n_9), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_347), .A2(n_278), .B1(n_219), .B2(n_268), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_360), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_360), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_341), .B(n_278), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_362), .Y(n_411) );
NAND2x1_ASAP7_75t_SL g412 ( .A(n_382), .B(n_345), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_368), .B(n_342), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_379), .B(n_325), .Y(n_414) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_395), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_368), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_371), .B(n_342), .Y(n_417) );
NOR2xp33_ASAP7_75t_SL g418 ( .A(n_372), .B(n_328), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_373), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_399), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_373), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_393), .A2(n_345), .B1(n_338), .B2(n_328), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_376), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_380), .B(n_356), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_389), .B(n_339), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_366), .Y(n_426) );
NOR2x1_ASAP7_75t_L g427 ( .A(n_391), .B(n_345), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_405), .A2(n_354), .B(n_336), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_379), .B(n_325), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_399), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_376), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_363), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_383), .B(n_325), .Y(n_433) );
INVxp67_ASAP7_75t_SL g434 ( .A(n_395), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_383), .B(n_325), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_364), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_394), .B(n_328), .Y(n_437) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_395), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_386), .B(n_338), .Y(n_439) );
OA21x2_ASAP7_75t_L g440 ( .A1(n_388), .A2(n_342), .B(n_352), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_386), .B(n_352), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_365), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_369), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_374), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_387), .B(n_352), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_372), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_371), .B(n_344), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_387), .B(n_344), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_361), .B(n_325), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_392), .B(n_344), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_378), .B(n_340), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_361), .B(n_343), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_378), .B(n_340), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_392), .B(n_340), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_420), .B(n_398), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_426), .A2(n_404), .B1(n_367), .B2(n_406), .C(n_375), .Y(n_456) );
AOI31xp33_ASAP7_75t_L g457 ( .A1(n_415), .A2(n_403), .A3(n_405), .B(n_401), .Y(n_457) );
NOR2x1_ASAP7_75t_L g458 ( .A(n_427), .B(n_409), .Y(n_458) );
AOI211xp5_ASAP7_75t_L g459 ( .A1(n_437), .A2(n_401), .B(n_403), .C(n_402), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_416), .B(n_397), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_424), .A2(n_367), .B1(n_397), .B2(n_402), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_411), .Y(n_462) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_413), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_411), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_430), .A2(n_384), .B1(n_377), .B2(n_385), .C(n_400), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_446), .A2(n_407), .B1(n_400), .B2(n_345), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_413), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_432), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_412), .A2(n_410), .B(n_370), .C(n_343), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_417), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_452), .B(n_410), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_446), .A2(n_381), .B1(n_370), .B2(n_354), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_441), .B(n_381), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_425), .B(n_408), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_434), .A2(n_396), .B1(n_390), .B2(n_388), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_436), .A2(n_263), .B1(n_12), .B2(n_13), .C(n_14), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_418), .A2(n_268), .B1(n_208), .B2(n_15), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_445), .B(n_9), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_452), .B(n_14), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_442), .B(n_16), .Y(n_480) );
O2A1O1Ixp5_ASAP7_75t_L g481 ( .A1(n_438), .A2(n_208), .B(n_16), .C(n_20), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_443), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_457), .A2(n_428), .B(n_440), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_456), .A2(n_439), .B1(n_454), .B2(n_450), .C(n_448), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_466), .A2(n_429), .B1(n_414), .B2(n_433), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_457), .A2(n_453), .B(n_451), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_465), .A2(n_429), .B1(n_414), .B2(n_433), .C(n_435), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_462), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_469), .A2(n_412), .B(n_449), .C(n_422), .Y(n_490) );
OAI21xp33_ASAP7_75t_SL g491 ( .A1(n_463), .A2(n_449), .B(n_435), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_458), .B(n_453), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_479), .A2(n_451), .B1(n_447), .B2(n_417), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_471), .B(n_447), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_464), .Y(n_495) );
AOI221x1_ASAP7_75t_L g496 ( .A1(n_480), .A2(n_431), .B1(n_423), .B2(n_421), .C(n_419), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_468), .Y(n_497) );
AOI21xp33_ASAP7_75t_SL g498 ( .A1(n_472), .A2(n_440), .B(n_431), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g499 ( .A1(n_482), .A2(n_423), .B1(n_421), .B2(n_419), .C(n_440), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_459), .A2(n_19), .B(n_21), .C(n_23), .Y(n_500) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_498), .A2(n_475), .B1(n_470), .B2(n_461), .C(n_483), .Y(n_501) );
OAI211xp5_ASAP7_75t_L g502 ( .A1(n_491), .A2(n_478), .B(n_476), .C(n_477), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_490), .B(n_481), .C(n_470), .D(n_474), .Y(n_503) );
OAI221xp5_ASAP7_75t_SL g504 ( .A1(n_488), .A2(n_455), .B1(n_467), .B2(n_473), .C(n_460), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g505 ( .A1(n_485), .A2(n_168), .B1(n_25), .B2(n_26), .C(n_27), .Y(n_505) );
AOI221xp5_ASAP7_75t_L g506 ( .A1(n_487), .A2(n_24), .B1(n_29), .B2(n_31), .C(n_33), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_486), .A2(n_34), .B1(n_35), .B2(n_37), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_493), .A2(n_39), .B1(n_40), .B2(n_42), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_497), .Y(n_509) );
OAI211xp5_ASAP7_75t_L g510 ( .A1(n_501), .A2(n_484), .B(n_500), .C(n_496), .Y(n_510) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_505), .B(n_484), .C(n_499), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_504), .B(n_492), .Y(n_512) );
OR5x1_ASAP7_75t_L g513 ( .A(n_503), .B(n_489), .C(n_495), .D(n_494), .E(n_47), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_502), .B(n_43), .C(n_45), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g515 ( .A(n_510), .B(n_506), .C(n_508), .Y(n_515) );
NOR2x2_ASAP7_75t_L g516 ( .A(n_513), .B(n_507), .Y(n_516) );
XNOR2x1_ASAP7_75t_SL g517 ( .A(n_514), .B(n_509), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_517), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_515), .Y(n_519) );
XNOR2xp5_ASAP7_75t_L g520 ( .A(n_519), .B(n_511), .Y(n_520) );
OAI22x1_ASAP7_75t_L g521 ( .A1(n_520), .A2(n_518), .B1(n_512), .B2(n_516), .Y(n_521) );
AOI222xp33_ASAP7_75t_SL g522 ( .A1(n_521), .A2(n_518), .B1(n_53), .B2(n_56), .C1(n_58), .C2(n_59), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_522), .A2(n_46), .B(n_61), .Y(n_523) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_523), .A2(n_66), .B(n_68), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_524), .A2(n_72), .B1(n_74), .B2(n_75), .Y(n_525) );
endmodule