module fake_jpeg_21250_n_270 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_270);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_18),
.B1(n_14),
.B2(n_16),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_42),
.B1(n_17),
.B2(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_34),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_14),
.B1(n_17),
.B2(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_14),
.B1(n_23),
.B2(n_17),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_46),
.B(n_50),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_39),
.B1(n_40),
.B2(n_45),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_42),
.B1(n_40),
.B2(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_52),
.B1(n_43),
.B2(n_49),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_35),
.B1(n_14),
.B2(n_37),
.Y(n_73)
);

OAI22x1_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_54),
.B1(n_56),
.B2(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_42),
.CI(n_39),
.CON(n_79),
.SN(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_87),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_71),
.C(n_65),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_86),
.B(n_90),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_98),
.B1(n_79),
.B2(n_36),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_68),
.B(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_55),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_78),
.B1(n_81),
.B2(n_62),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_57),
.B1(n_56),
.B2(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_63),
.B(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_67),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_92),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_64),
.A2(n_57),
.B1(n_61),
.B2(n_53),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_54),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_95),
.B(n_74),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_51),
.C(n_35),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_69),
.C(n_80),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_36),
.B1(n_54),
.B2(n_35),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_34),
.Y(n_99)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_70),
.B1(n_68),
.B2(n_79),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_106),
.B1(n_113),
.B2(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_109),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_105),
.A2(n_110),
.B1(n_33),
.B2(n_29),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_73),
.B1(n_36),
.B2(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_67),
.B1(n_54),
.B2(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_112),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_118),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_75),
.B1(n_80),
.B2(n_69),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_80),
.B1(n_69),
.B2(n_44),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_98),
.B1(n_99),
.B2(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_127),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_90),
.C(n_87),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_76),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_89),
.B(n_88),
.C(n_99),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_134),
.B(n_138),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_29),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_110),
.B1(n_105),
.B2(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_91),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_120),
.B(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_84),
.B(n_93),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_7),
.B(n_11),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_141),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_108),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_SL g164 ( 
.A(n_142),
.B(n_143),
.C(n_145),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_74),
.B(n_76),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_106),
.B1(n_111),
.B2(n_81),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_74),
.B1(n_76),
.B2(n_81),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_153),
.B1(n_167),
.B2(n_169),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_151),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_156),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_78),
.B1(n_33),
.B2(n_29),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_127),
.B(n_137),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_11),
.B(n_10),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_137),
.B(n_24),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_123),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_13),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_141),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_78),
.B1(n_28),
.B2(n_0),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_78),
.B1(n_28),
.B2(n_22),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_145),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_28),
.B1(n_1),
.B2(n_0),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_145),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_171),
.A2(n_175),
.B(n_126),
.Y(n_198)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_181),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_145),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_165),
.A2(n_130),
.B1(n_129),
.B2(n_143),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_22),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_143),
.B1(n_122),
.B2(n_124),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_143),
.B1(n_136),
.B2(n_131),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_125),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_134),
.C(n_132),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_158),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_136),
.C(n_131),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_156),
.C(n_162),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_147),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_173),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_184),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_150),
.B1(n_169),
.B2(n_153),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_197),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_13),
.B1(n_15),
.B2(n_2),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_126),
.C(n_167),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_201),
.C(n_202),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_8),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_22),
.C(n_21),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_22),
.C(n_21),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_177),
.C(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_203),
.B(n_207),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_175),
.B1(n_171),
.B2(n_188),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_221),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_210),
.A2(n_216),
.B1(n_193),
.B2(n_20),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_195),
.B(n_187),
.CI(n_179),
.CON(n_211),
.SN(n_211)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_214),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_191),
.A2(n_200),
.B1(n_196),
.B2(n_203),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_199),
.B1(n_192),
.B2(n_198),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_201),
.A2(n_183),
.B1(n_187),
.B2(n_21),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_208),
.B1(n_197),
.B2(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_8),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_15),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_204),
.A2(n_7),
.B(n_9),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_229),
.B1(n_210),
.B2(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_228),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_6),
.B1(n_10),
.B2(n_2),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_20),
.B1(n_19),
.B2(n_12),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_230),
.B(n_233),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_209),
.C(n_216),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_232),
.C(n_223),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_20),
.C(n_19),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_15),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_5),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_234),
.B1(n_227),
.B2(n_229),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_217),
.B(n_211),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_238),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_211),
.B(n_6),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_242),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_19),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_0),
.C(n_1),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_245),
.A2(n_3),
.B(n_4),
.Y(n_258)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_250),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_243),
.B(n_5),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_5),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_0),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_240),
.C(n_6),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_3),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_246),
.B(n_247),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_10),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_257),
.C(n_255),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_264),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_260),
.C(n_3),
.Y(n_266)
);

OAI221xp5_ASAP7_75t_L g267 ( 
.A1(n_266),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.C(n_1),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_267),
.A2(n_1),
.B(n_4),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_1),
.C(n_9),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);


endmodule