module fake_jpeg_13794_n_158 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_40),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_80),
.Y(n_83)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_77),
.B(n_79),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_49),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_50),
.Y(n_81)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_0),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_65),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_49),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_63),
.C(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_92),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_63),
.B1(n_57),
.B2(n_59),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_60),
.B1(n_52),
.B2(n_69),
.Y(n_104)
);

OR2x2_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_60),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_65),
.C(n_71),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_68),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_81),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_99),
.C(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_10),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_108),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_61),
.C(n_59),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_109),
.B1(n_112),
.B2(n_97),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_110),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_69),
.B1(n_75),
.B2(n_52),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_1),
.B(n_2),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_10),
.B(n_12),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_27),
.C(n_46),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_87),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_117),
.Y(n_135)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_89),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_28),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_3),
.B1(n_7),
.B2(n_9),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_124),
.B1(n_24),
.B2(n_29),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_9),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_122),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_130),
.B(n_13),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_34),
.B1(n_45),
.B2(n_15),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_125),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_47),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_22),
.Y(n_136)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_39),
.C(n_42),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_13),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_133),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_44),
.C(n_23),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_137),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

OA21x2_ASAP7_75t_SL g147 ( 
.A1(n_140),
.A2(n_142),
.B(n_143),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_43),
.B1(n_124),
.B2(n_121),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_114),
.B(n_123),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_148),
.A2(n_127),
.B(n_117),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_151),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_135),
.C(n_143),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_152),
.A2(n_148),
.B1(n_135),
.B2(n_149),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_153),
.B1(n_134),
.B2(n_147),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_154),
.Y(n_157)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_145),
.B1(n_138),
.B2(n_141),
.C(n_120),
.Y(n_158)
);


endmodule