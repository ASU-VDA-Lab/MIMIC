module fake_jpeg_19947_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx9p33_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_17),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g31 ( 
.A1(n_17),
.A2(n_0),
.B(n_2),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_35),
.Y(n_41)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_15),
.B1(n_19),
.B2(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_52),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_19),
.B1(n_27),
.B2(n_24),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_46),
.B1(n_56),
.B2(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_14),
.B1(n_23),
.B2(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_53),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_14),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_23),
.B1(n_18),
.B2(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_76),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_30),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_66),
.B(n_68),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_37),
.B(n_35),
.C(n_38),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_54),
.B1(n_45),
.B2(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_38),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_20),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_37),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_84),
.C(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_55),
.B1(n_67),
.B2(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_65),
.C(n_68),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_36),
.C(n_37),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_68),
.B(n_75),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_93),
.B(n_67),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_35),
.B(n_27),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_87),
.B1(n_88),
.B2(n_84),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_71),
.B1(n_72),
.B2(n_59),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_99),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_92),
.B(n_93),
.C(n_91),
.D(n_80),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_105),
.C(n_85),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_90),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_60),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_109),
.B(n_94),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_91),
.C(n_89),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_59),
.Y(n_119)
);

OAI321xp33_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_95),
.A3(n_100),
.B1(n_104),
.B2(n_102),
.C(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_117),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_106),
.B(n_110),
.C(n_101),
.D(n_113),
.Y(n_115)
);

AOI321xp33_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_118),
.A3(n_20),
.B1(n_36),
.B2(n_26),
.C(n_12),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_96),
.B1(n_94),
.B2(n_98),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_55),
.B1(n_77),
.B2(n_64),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_120),
.Y(n_121)
);

AOI221xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_57),
.B1(n_20),
.B2(n_26),
.C(n_99),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_78),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_2),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_124),
.A2(n_115),
.B(n_9),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_125),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_127),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_129),
.B1(n_121),
.B2(n_125),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_10),
.B1(n_11),
.B2(n_4),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_10),
.C(n_4),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_5),
.B1(n_127),
.B2(n_130),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_132),
.C(n_5),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);


endmodule