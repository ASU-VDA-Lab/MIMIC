module fake_netlist_5_1434_n_107 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_107);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_107;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVxp33_ASAP7_75t_SL g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_0),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_20),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_4),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_5),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2x1p5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NAND2x1p5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_46),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_53),
.B(n_55),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_60),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_56),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_44),
.B(n_32),
.C(n_35),
.Y(n_70)
);

AO21x2_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_44),
.B(n_54),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_67),
.B(n_68),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_63),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_21),
.B(n_22),
.C(n_63),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_74),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_65),
.C(n_70),
.Y(n_79)
);

AND2x4_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_51),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_81),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_71),
.Y(n_86)
);

OAI21x1_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_64),
.B(n_52),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_66),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_84),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_91),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_67),
.B(n_43),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_87),
.B(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_67),
.Y(n_101)
);

OAI221xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_96),
.B1(n_97),
.B2(n_68),
.C(n_64),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_101),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_100),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_102),
.B1(n_97),
.B2(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_39),
.B1(n_13),
.B2(n_11),
.C(n_64),
.Y(n_107)
);


endmodule