module fake_jpeg_2495_n_201 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_201);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_17),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_0),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_76),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_88),
.Y(n_93)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_63),
.B1(n_62),
.B2(n_65),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_66),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_73),
.Y(n_87)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_58),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_66),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_84),
.B1(n_88),
.B2(n_80),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_95),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_57),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_61),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_103),
.Y(n_127)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_82),
.B1(n_89),
.B2(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_82),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_53),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_113),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_62),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_49),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_53),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_125),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_50),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_124),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_48),
.B1(n_56),
.B2(n_55),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_51),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_150),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_127),
.A2(n_48),
.B1(n_92),
.B2(n_54),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_144),
.B1(n_67),
.B2(n_3),
.Y(n_157)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_136),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_67),
.B1(n_54),
.B2(n_20),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_139),
.B(n_141),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_111),
.B1(n_123),
.B2(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_1),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_145),
.B(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_149),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_1),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_67),
.C(n_54),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_158),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_21),
.C(n_45),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_156),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_146),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_161),
.B1(n_164),
.B2(n_167),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_169),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

NOR4xp25_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_22),
.C(n_43),
.D(n_41),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_18),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_129),
.C(n_130),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_175),
.C(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_174),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_153),
.B(n_44),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_39),
.B(n_37),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_175),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_36),
.C(n_35),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_179),
.A2(n_152),
.B1(n_154),
.B2(n_151),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_178),
.B1(n_159),
.B2(n_172),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_185),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_180),
.A2(n_157),
.B(n_155),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_29),
.B(n_28),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_152),
.C(n_33),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_190),
.B(n_186),
.Y(n_195)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_191),
.B(n_192),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_6),
.B(n_8),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_195),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_194),
.B(n_14),
.Y(n_197)
);

OAI221xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_196),
.B(n_12),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_10),
.B(n_13),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_13),
.Y(n_201)
);


endmodule