module fake_jpeg_14833_n_354 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_354);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_354;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_28),
.Y(n_74)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_29),
.B(n_27),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_23),
.Y(n_101)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_24),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_41),
.C(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_34),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_27),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_80),
.B(n_84),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_34),
.Y(n_81)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_37),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_91),
.Y(n_142)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_35),
.B1(n_45),
.B2(n_44),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_90),
.A2(n_30),
.B1(n_43),
.B2(n_53),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_28),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_31),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_102),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_37),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_103),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_35),
.B1(n_21),
.B2(n_30),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_98),
.B1(n_110),
.B2(n_66),
.Y(n_115)
);

BUFx2_ASAP7_75t_SL g97 ( 
.A(n_66),
.Y(n_97)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_70),
.Y(n_98)
);

BUFx4f_ASAP7_75t_SL g100 ( 
.A(n_71),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_100),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_51),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_21),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_64),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_109),
.Y(n_135)
);

CKINVDCx12_ASAP7_75t_R g109 ( 
.A(n_58),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_75),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_114),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_61),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_119),
.B1(n_140),
.B2(n_141),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_145),
.Y(n_154)
);

FAx1_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_68),
.CI(n_51),
.CON(n_118),
.SN(n_118)
);

XOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_118),
.B(n_146),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_68),
.B1(n_72),
.B2(n_67),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_41),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_96),
.Y(n_149)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_45),
.B1(n_44),
.B2(n_50),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

NAND2x1p5_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_49),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_158),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_152),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_117),
.B(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_49),
.C(n_100),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_89),
.B1(n_104),
.B2(n_83),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_155),
.B1(n_122),
.B2(n_140),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_119),
.A2(n_78),
.B1(n_83),
.B2(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_112),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_162),
.A2(n_169),
.B1(n_147),
.B2(n_144),
.Y(n_174)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

AOI22x1_ASAP7_75t_SL g165 ( 
.A1(n_146),
.A2(n_90),
.B1(n_38),
.B2(n_25),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_125),
.B(n_142),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_106),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_110),
.A3(n_22),
.B1(n_25),
.B2(n_38),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_141),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_174),
.A2(n_156),
.B1(n_98),
.B2(n_82),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_182),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_183),
.A2(n_185),
.B(n_187),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_117),
.B(n_118),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_133),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_192),
.B(n_171),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_201),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_135),
.B(n_133),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_26),
.B(n_32),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_196),
.A2(n_199),
.B1(n_85),
.B2(n_124),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_122),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_200),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_136),
.B1(n_144),
.B2(n_147),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_120),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

INVx4_ASAP7_75t_SL g208 ( 
.A(n_179),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_208),
.A2(n_179),
.B1(n_193),
.B2(n_182),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_157),
.Y(n_211)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_155),
.B1(n_168),
.B2(n_160),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_221),
.B1(n_228),
.B2(n_183),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_164),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_163),
.Y(n_216)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_218),
.B(n_226),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_SL g245 ( 
.A1(n_219),
.A2(n_222),
.B(n_224),
.Y(n_245)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_225),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_120),
.B1(n_156),
.B2(n_121),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_87),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_229),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_192),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_180),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_124),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_22),
.Y(n_251)
);

AND2x6_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_0),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_38),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_175),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_26),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_94),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_199),
.B(n_196),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_233),
.A2(n_240),
.B(n_232),
.Y(n_266)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_237),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_175),
.C(n_177),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_249),
.C(n_234),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_223),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_94),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_252),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_203),
.A2(n_207),
.B1(n_206),
.B2(n_214),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_256),
.B1(n_257),
.B2(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_26),
.C(n_32),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_25),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_254),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_20),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_22),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_206),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_257)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_212),
.B1(n_209),
.B2(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

HAxp5_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_229),
.CON(n_262),
.SN(n_262)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_267),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_204),
.B1(n_228),
.B2(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_225),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_266),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_R g267 ( 
.A1(n_245),
.A2(n_232),
.B1(n_222),
.B2(n_221),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_270),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_218),
.Y(n_271)
);

AOI21xp33_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_220),
.B(n_208),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_274),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_20),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_253),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_280),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_235),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_277),
.B1(n_256),
.B2(n_254),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_233),
.A2(n_20),
.B1(n_7),
.B2(n_8),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_255),
.C(n_249),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_238),
.A2(n_6),
.B(n_8),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_283),
.C(n_287),
.Y(n_310)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_248),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_242),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_291),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_244),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_244),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_259),
.Y(n_305)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_237),
.Y(n_300)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_269),
.C(n_243),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_282),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_261),
.B1(n_266),
.B2(n_265),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_303),
.A2(n_287),
.B1(n_291),
.B2(n_283),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_314),
.C(n_285),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_261),
.B(n_276),
.Y(n_307)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_277),
.B1(n_262),
.B2(n_280),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_6),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_286),
.B(n_14),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_296),
.B(n_8),
.Y(n_311)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_293),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_312),
.B(n_313),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_292),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_290),
.B(n_11),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_323),
.C(n_310),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_299),
.Y(n_317)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_317),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_303),
.B(n_15),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_319),
.B(n_302),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_326),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_281),
.C(n_285),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_329),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_321),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g337 ( 
.A1(n_330),
.A2(n_324),
.A3(n_318),
.B1(n_326),
.B2(n_323),
.C1(n_315),
.C2(n_40),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_320),
.A2(n_304),
.B1(n_306),
.B2(n_314),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_322),
.A2(n_306),
.B1(n_15),
.B2(n_16),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_333),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_40),
.Y(n_339)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_337),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_335),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_338),
.B(n_341),
.Y(n_346)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_339),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_11),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_17),
.Y(n_345)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_345),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_346),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_347),
.B(n_343),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_340),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_348),
.C(n_344),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_351),
.A2(n_336),
.B(n_342),
.Y(n_352)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_15),
.B(n_16),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_17),
.Y(n_354)
);


endmodule