module fake_jpeg_23025_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_42),
.Y(n_53)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_0),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_23),
.B(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_47),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_23),
.B1(n_34),
.B2(n_17),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_55),
.B1(n_23),
.B2(n_31),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_26),
.B1(n_21),
.B2(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_59),
.B(n_67),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_23),
.B1(n_26),
.B2(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_60),
.A2(n_68),
.B1(n_31),
.B2(n_24),
.Y(n_102)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_65),
.Y(n_88)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2x1_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_27),
.B1(n_26),
.B2(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_25),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_24),
.Y(n_89)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_74),
.Y(n_101)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_44),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_28),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_78),
.B(n_82),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_31),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_61),
.C(n_39),
.Y(n_142)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_64),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_83),
.A2(n_87),
.B1(n_100),
.B2(n_71),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_85),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_55),
.B1(n_21),
.B2(n_31),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_62),
.B1(n_66),
.B2(n_65),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_89),
.B(n_111),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_35),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_36),
.A3(n_44),
.B1(n_43),
.B2(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_94),
.Y(n_115)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_47),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_47),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_99),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_34),
.B(n_25),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_90),
.B(n_78),
.C(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_47),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_104),
.B(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_47),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_108),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_32),
.B1(n_24),
.B2(n_27),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_73),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_40),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_48),
.B(n_25),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_58),
.A2(n_32),
.B1(n_33),
.B2(n_30),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_123),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_0),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_119),
.B(n_125),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_54),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_79),
.A2(n_43),
.B(n_36),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_133),
.B1(n_82),
.B2(n_77),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_80),
.B(n_30),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_80),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_40),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_134),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_83),
.A2(n_33),
.B1(n_30),
.B2(n_39),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_19),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_0),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_142),
.C(n_81),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_19),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_86),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_61),
.B1(n_39),
.B2(n_16),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_112),
.B1(n_92),
.B2(n_77),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_105),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_145),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_147),
.B(n_150),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_131),
.Y(n_196)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_173),
.B(n_135),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_96),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_159),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_91),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_155),
.C(n_160),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_120),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_115),
.A2(n_86),
.B1(n_108),
.B2(n_103),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_167),
.B1(n_174),
.B2(n_139),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_100),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_88),
.B(n_107),
.C(n_101),
.D(n_85),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_175),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_105),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_112),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_168),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_128),
.B1(n_138),
.B2(n_137),
.Y(n_179)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_109),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_176),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_114),
.C(n_84),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_116),
.Y(n_192)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_124),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_131),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_95),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_172),
.B(n_118),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_114),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_115),
.A2(n_93),
.B1(n_33),
.B2(n_35),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_117),
.B(n_19),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_18),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_116),
.B(n_29),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_179),
.A2(n_182),
.B1(n_190),
.B2(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_138),
.B1(n_139),
.B2(n_123),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_183),
.A2(n_198),
.B1(n_20),
.B2(n_18),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_205),
.B(n_178),
.Y(n_223)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_200),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_173),
.A2(n_139),
.B1(n_135),
.B2(n_123),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_139),
.B1(n_124),
.B2(n_129),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_196),
.C(n_199),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_137),
.B1(n_121),
.B2(n_126),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_131),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_173),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_211),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_158),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_154),
.A2(n_121),
.B(n_35),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_118),
.B1(n_20),
.B2(n_127),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_208),
.B1(n_165),
.B2(n_168),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_149),
.B(n_127),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_177),
.C(n_176),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_167),
.A2(n_150),
.B1(n_161),
.B2(n_146),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_127),
.Y(n_209)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_145),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_183),
.A2(n_148),
.B1(n_146),
.B2(n_170),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_239),
.B1(n_210),
.B2(n_180),
.Y(n_242)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_225),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_218),
.B(n_219),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_187),
.B(n_160),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_230),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_211),
.B(n_147),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_222),
.B(n_228),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_SL g244 ( 
.A1(n_223),
.A2(n_234),
.B(n_197),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_184),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_157),
.B(n_154),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_226),
.A2(n_231),
.B(n_237),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_174),
.Y(n_228)
);

XOR2x2_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_153),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_229),
.B(n_199),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_236),
.C(n_7),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_18),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_1),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_20),
.C(n_18),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_189),
.Y(n_237)
);

BUFx12f_ASAP7_75t_SL g238 ( 
.A(n_190),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_238),
.A2(n_1),
.B(n_2),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_226),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_246),
.B1(n_259),
.B2(n_228),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_195),
.B1(n_202),
.B2(n_198),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_247),
.B1(n_249),
.B2(n_256),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_217),
.A2(n_195),
.B1(n_185),
.B2(n_201),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_205),
.B1(n_201),
.B2(n_192),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_251),
.C(n_254),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_207),
.B1(n_196),
.B2(n_3),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_1),
.C(n_2),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_227),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_255),
.B(n_221),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_7),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_260),
.C(n_262),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_217),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_233),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_212),
.B(n_3),
.C(n_4),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_280),
.B1(n_234),
.B2(n_249),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_243),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_271),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_237),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_274),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_220),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_219),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_276),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_213),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_250),
.B(n_215),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_279),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_282),
.B1(n_246),
.B2(n_254),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_259),
.B(n_235),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_263),
.A2(n_232),
.B1(n_243),
.B2(n_256),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_245),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_284),
.B(n_282),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_260),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_287),
.Y(n_298)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_248),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_258),
.C(n_242),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_292),
.C(n_296),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_247),
.C(n_251),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_267),
.A2(n_253),
.B1(n_223),
.B2(n_236),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_280),
.Y(n_301)
);

NOR2x1_ASAP7_75t_R g295 ( 
.A(n_274),
.B(n_11),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_295),
.A2(n_264),
.B(n_265),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_4),
.C(n_5),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_307),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_266),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_306),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_309),
.B1(n_310),
.B2(n_15),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_281),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_304),
.B(n_305),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_264),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_283),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_270),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_308),
.B(n_8),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_270),
.B1(n_5),
.B2(n_6),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_291),
.B1(n_292),
.B2(n_288),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_287),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_313),
.Y(n_321)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_295),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_8),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_320),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_306),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_4),
.C(n_6),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_325),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_302),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_316),
.A3(n_315),
.B1(n_320),
.B2(n_15),
.C1(n_12),
.C2(n_11),
.Y(n_328)
);

MAJx2_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_298),
.C(n_12),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_298),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_14),
.A3(n_15),
.B1(n_316),
.B2(n_321),
.C1(n_326),
.C2(n_324),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_328),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_332),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_330),
.B1(n_331),
.B2(n_14),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_14),
.Y(n_336)
);


endmodule