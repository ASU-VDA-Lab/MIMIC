module fake_jpeg_14472_n_199 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_199);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_5),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_4),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_19),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_91),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_1),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_89),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_61),
.B1(n_67),
.B2(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_88),
.B1(n_82),
.B2(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_104),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_61),
.B1(n_67),
.B2(n_63),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_60),
.B1(n_62),
.B2(n_78),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_58),
.B1(n_57),
.B2(n_68),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_76),
.B(n_79),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_85),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_69),
.B1(n_58),
.B2(n_70),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_109),
.B1(n_79),
.B2(n_3),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_69),
.B1(n_58),
.B2(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_126),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_116),
.Y(n_154)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_130),
.B(n_2),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_82),
.B1(n_81),
.B2(n_75),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_120),
.B1(n_124),
.B2(n_131),
.Y(n_149)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_108),
.B(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_125),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_72),
.B1(n_71),
.B2(n_65),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_84),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_1),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_9),
.Y(n_141)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_25),
.C(n_52),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_137),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_24),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_142),
.B1(n_29),
.B2(n_31),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_20),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_153),
.B1(n_21),
.B2(n_22),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_27),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_130),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_146),
.C(n_53),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_137),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_163),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_153),
.B1(n_144),
.B2(n_137),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_167),
.B1(n_168),
.B2(n_171),
.Y(n_180)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_147),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_146),
.B1(n_143),
.B2(n_43),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_40),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_45),
.B(n_51),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_136),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_179),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_41),
.C(n_44),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_181),
.B(n_172),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g184 ( 
.A(n_177),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_185),
.Y(n_189)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_178),
.A2(n_172),
.B1(n_160),
.B2(n_170),
.C(n_167),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_175),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_183),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_183),
.B(n_186),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_191),
.C(n_190),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_189),
.C(n_174),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_176),
.B(n_182),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_180),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_196),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_181),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_171),
.Y(n_199)
);


endmodule