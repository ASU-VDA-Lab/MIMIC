module fake_jpeg_24504_n_132 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_30),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_0),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_31),
.A2(n_28),
.B1(n_27),
.B2(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_38),
.Y(n_43)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_1),
.C(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_3),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_27),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_60),
.C(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_58),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_26),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_9),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_67),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_14),
.C(n_24),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_40),
.B1(n_35),
.B2(n_16),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_76),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_40),
.C(n_25),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_25),
.C(n_20),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_22),
.B1(n_6),
.B2(n_4),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_78),
.B1(n_50),
.B2(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_22),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_4),
.B1(n_6),
.B2(n_22),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_11),
.B(n_12),
.Y(n_88)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_59),
.B1(n_50),
.B2(n_52),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_78),
.B1(n_72),
.B2(n_46),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_77),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_80),
.B(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_95),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_52),
.B(n_43),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_73),
.B(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_63),
.B(n_46),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_82),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_72),
.B1(n_46),
.B2(n_53),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_85),
.B1(n_86),
.B2(n_44),
.Y(n_110)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_73),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_46),
.C(n_44),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_106),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_93),
.B1(n_83),
.B2(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_114),
.B(n_96),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_105),
.C(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_101),
.Y(n_118)
);

AOI321xp33_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_101),
.A3(n_106),
.B1(n_108),
.B2(n_103),
.C(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_103),
.B1(n_104),
.B2(n_87),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_107),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_107),
.C(n_108),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_116),
.B(n_84),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_115),
.C(n_105),
.Y(n_126)
);

OAI21x1_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_128),
.B(n_124),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_130),
.B1(n_44),
.B2(n_79),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_127),
.A2(n_102),
.B(n_85),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_79),
.Y(n_132)
);


endmodule