module fake_netlist_6_4094_n_334 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_98, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_77, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_104, n_95, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_103, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_334);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_77;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_104;
input n_95;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_103;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_334;

wire n_326;
wire n_256;
wire n_209;
wire n_223;
wire n_278;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_168;
wire n_125;
wire n_297;
wire n_106;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_142;
wire n_143;
wire n_180;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_280;
wire n_287;
wire n_230;
wire n_141;
wire n_200;
wire n_176;
wire n_114;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_111;
wire n_314;
wire n_183;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_129;
wire n_197;
wire n_137;
wire n_155;
wire n_109;
wire n_122;
wire n_218;
wire n_234;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_107;
wire n_272;
wire n_185;
wire n_293;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_265;
wire n_260;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_166;
wire n_184;
wire n_216;
wire n_323;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_204;
wire n_261;
wire n_312;
wire n_130;
wire n_164;
wire n_292;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_237;
wire n_244;
wire n_243;
wire n_124;
wire n_282;
wire n_116;
wire n_211;
wire n_175;
wire n_117;
wire n_322;
wire n_231;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_317;
wire n_149;
wire n_328;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_324;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_267;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_259;
wire n_177;
wire n_295;
wire n_190;
wire n_262;
wire n_187;
wire n_170;
wire n_332;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

INVxp33_ASAP7_75t_SL g107 ( 
.A(n_5),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_12),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_5),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_31),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_17),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_14),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_41),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_26),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_6),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_10),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_39),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_50),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_34),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_45),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_16),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_25),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_15),
.Y(n_144)
);

INVxp67_ASAP7_75t_SL g145 ( 
.A(n_78),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_49),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_10),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g149 ( 
.A(n_46),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_24),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_51),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_19),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_48),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_94),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_60),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_42),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_76),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_128),
.B(n_0),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_0),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_1),
.B(n_2),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_3),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_13),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_4),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_133),
.B(n_7),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g183 ( 
.A1(n_112),
.A2(n_8),
.B(n_9),
.Y(n_183)
);

AND3x2_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_9),
.C(n_11),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_164),
.B(n_107),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_123),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

AO22x2_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_119),
.B1(n_158),
.B2(n_136),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_187),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

OAI221xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_125),
.B1(n_147),
.B2(n_114),
.C(n_159),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_160),
.B1(n_126),
.B2(n_121),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_115),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_141),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_116),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_189),
.B(n_120),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_183),
.B1(n_170),
.B2(n_180),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_181),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_169),
.B1(n_172),
.B2(n_167),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_170),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_216),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_170),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_192),
.Y(n_230)
);

OR2x2_ASAP7_75t_SL g231 ( 
.A(n_210),
.B(n_183),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_117),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_145),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_149),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_155),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_206),
.B(n_214),
.C(n_215),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_237),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

BUFx8_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

OR2x6_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_196),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_224),
.A2(n_196),
.B1(n_190),
.B2(n_124),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_205),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_139),
.B(n_122),
.C(n_144),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_197),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_218),
.A2(n_130),
.B(n_134),
.C(n_137),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_152),
.B1(n_143),
.B2(n_146),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_231),
.A2(n_154),
.B1(n_153),
.B2(n_140),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_151),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_200),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_235),
.A2(n_195),
.B(n_201),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_156),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_238),
.A2(n_18),
.B(n_20),
.Y(n_268)
);

OAI22x1_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_184),
.B1(n_21),
.B2(n_23),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_271)
);

NAND2x1p5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_254),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_243),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_229),
.B(n_223),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_233),
.B(n_232),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_229),
.B(n_223),
.Y(n_281)
);

INVx5_ASAP7_75t_SL g282 ( 
.A(n_252),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g284 ( 
.A1(n_262),
.A2(n_246),
.B(n_268),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_259),
.A2(n_240),
.B1(n_33),
.B2(n_35),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_30),
.B(n_36),
.C(n_37),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_255),
.A2(n_38),
.B(n_40),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_43),
.B(n_44),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_252),
.A2(n_269),
.B1(n_263),
.B2(n_271),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_267),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

OAI221xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_248),
.B1(n_251),
.B2(n_56),
.C(n_57),
.Y(n_293)
);

AO21x2_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_54),
.B(n_55),
.Y(n_294)
);

OR2x6_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_58),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_61),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_66),
.B1(n_68),
.B2(n_71),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_275),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_80),
.B(n_81),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_L g301 ( 
.A1(n_274),
.A2(n_103),
.B1(n_84),
.B2(n_85),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_82),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_274),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_298),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_279),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_309),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_298),
.B1(n_299),
.B2(n_294),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_280),
.Y(n_315)
);

OAI211xp5_ASAP7_75t_SL g316 ( 
.A1(n_308),
.A2(n_297),
.B(n_301),
.C(n_281),
.Y(n_316)
);

NAND5xp2_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_272),
.C(n_288),
.D(n_300),
.E(n_289),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_R g318 ( 
.A(n_311),
.B(n_300),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_315),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_319),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_321),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_316),
.B(n_312),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_SL g328 ( 
.A(n_327),
.B(n_318),
.C(n_317),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_SL g329 ( 
.A(n_328),
.B(n_272),
.C(n_87),
.Y(n_329)
);

XNOR2x1_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_86),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_278),
.B1(n_90),
.B2(n_91),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

AOI221xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.C(n_102),
.Y(n_334)
);


endmodule