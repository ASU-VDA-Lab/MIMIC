module real_aes_2048_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_0), .B(n_140), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_1), .A2(n_149), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_2), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_3), .B(n_140), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_4), .B(n_156), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_5), .B(n_156), .Y(n_517) );
INVx1_ASAP7_75t_L g147 ( .A(n_6), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_7), .B(n_156), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_8), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g786 ( .A1(n_9), .A2(n_55), .B1(n_787), .B2(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_9), .Y(n_787) );
NAND2xp33_ASAP7_75t_L g538 ( .A(n_10), .B(n_158), .Y(n_538) );
AND2x2_ASAP7_75t_L g176 ( .A(n_11), .B(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g253 ( .A(n_12), .B(n_165), .Y(n_253) );
INVx2_ASAP7_75t_L g162 ( .A(n_13), .Y(n_162) );
AOI221x1_ASAP7_75t_L g562 ( .A1(n_14), .A2(n_26), .B1(n_140), .B2(n_149), .C(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_15), .B(n_156), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_16), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_17), .B(n_140), .Y(n_534) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_18), .A2(n_165), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_19), .B(n_160), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_20), .B(n_156), .Y(n_494) );
AO21x1_ASAP7_75t_L g512 ( .A1(n_21), .A2(n_140), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_22), .B(n_140), .Y(n_207) );
INVx1_ASAP7_75t_L g115 ( .A(n_23), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_24), .A2(n_91), .B1(n_140), .B2(n_182), .Y(n_181) );
AOI22xp5_ASAP7_75t_SL g124 ( .A1(n_25), .A2(n_48), .B1(n_125), .B2(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g126 ( .A(n_25), .Y(n_126) );
NAND2x1_ASAP7_75t_L g555 ( .A(n_27), .B(n_156), .Y(n_555) );
NAND2x1_ASAP7_75t_L g504 ( .A(n_28), .B(n_158), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_29), .A2(n_123), .B1(n_124), .B2(n_127), .Y(n_122) );
INVx1_ASAP7_75t_L g127 ( .A(n_29), .Y(n_127) );
OR2x2_ASAP7_75t_L g163 ( .A(n_30), .B(n_88), .Y(n_163) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_30), .A2(n_88), .B(n_162), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_31), .B(n_158), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_32), .B(n_156), .Y(n_537) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_33), .A2(n_177), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_34), .B(n_158), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_35), .A2(n_149), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_36), .B(n_156), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_37), .A2(n_149), .B(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g146 ( .A(n_38), .B(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g150 ( .A(n_38), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g190 ( .A(n_38), .Y(n_190) );
OR2x6_ASAP7_75t_L g113 ( .A(n_39), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_40), .B(n_140), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_41), .B(n_140), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_42), .B(n_156), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_43), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_44), .B(n_158), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_45), .B(n_140), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_46), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_47), .A2(n_149), .B(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g125 ( .A(n_48), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_49), .A2(n_149), .B(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_50), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_51), .B(n_158), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_52), .B(n_140), .Y(n_231) );
INVx1_ASAP7_75t_L g143 ( .A(n_53), .Y(n_143) );
INVx1_ASAP7_75t_L g153 ( .A(n_53), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_54), .B(n_156), .Y(n_174) );
INVx1_ASAP7_75t_L g788 ( .A(n_55), .Y(n_788) );
AND2x2_ASAP7_75t_L g197 ( .A(n_56), .B(n_160), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_57), .B(n_158), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_58), .B(n_156), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_59), .B(n_158), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_60), .A2(n_149), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_61), .B(n_140), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_62), .B(n_140), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_63), .A2(n_149), .B(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g213 ( .A(n_64), .B(n_161), .Y(n_213) );
AO21x1_ASAP7_75t_L g514 ( .A1(n_65), .A2(n_149), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_66), .B(n_140), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_67), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_68), .B(n_158), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_69), .B(n_140), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_70), .B(n_158), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_71), .A2(n_95), .B1(n_149), .B2(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_72), .B(n_156), .Y(n_210) );
AND2x2_ASAP7_75t_L g528 ( .A(n_73), .B(n_161), .Y(n_528) );
INVx1_ASAP7_75t_L g145 ( .A(n_74), .Y(n_145) );
INVx1_ASAP7_75t_L g151 ( .A(n_74), .Y(n_151) );
AND2x2_ASAP7_75t_L g507 ( .A(n_75), .B(n_177), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_76), .B(n_158), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_77), .A2(n_149), .B(n_201), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_78), .A2(n_149), .B(n_154), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_79), .A2(n_149), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g225 ( .A(n_80), .B(n_161), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_81), .B(n_160), .Y(n_179) );
INVx1_ASAP7_75t_L g116 ( .A(n_82), .Y(n_116) );
AND2x2_ASAP7_75t_L g480 ( .A(n_83), .B(n_177), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_84), .B(n_140), .Y(n_496) );
AND2x2_ASAP7_75t_L g164 ( .A(n_85), .B(n_165), .Y(n_164) );
OAI22x1_ASAP7_75t_L g781 ( .A1(n_86), .A2(n_782), .B1(n_789), .B2(n_790), .Y(n_781) );
INVx1_ASAP7_75t_L g789 ( .A(n_86), .Y(n_789) );
AND2x2_ASAP7_75t_L g513 ( .A(n_87), .B(n_204), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_89), .B(n_158), .Y(n_495) );
AND2x2_ASAP7_75t_L g558 ( .A(n_90), .B(n_177), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_92), .B(n_156), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_93), .A2(n_149), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_94), .B(n_158), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_96), .A2(n_149), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_97), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_98), .B(n_156), .Y(n_485) );
BUFx2_ASAP7_75t_L g212 ( .A(n_99), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_100), .Y(n_799) );
BUFx2_ASAP7_75t_L g780 ( .A(n_101), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_102), .A2(n_149), .B(n_536), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_120), .B(n_798), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g800 ( .A(n_107), .Y(n_800) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_117), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_SL g792 ( .A(n_110), .Y(n_792) );
BUFx3_ASAP7_75t_L g796 ( .A(n_110), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x6_ASAP7_75t_SL g471 ( .A(n_111), .B(n_113), .Y(n_471) );
OR2x6_ASAP7_75t_SL g771 ( .A(n_111), .B(n_112), .Y(n_771) );
OR2x2_ASAP7_75t_L g777 ( .A(n_111), .B(n_113), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AO221x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_778), .B1(n_781), .B2(n_791), .C(n_793), .Y(n_120) );
OAI222xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_128), .B1(n_772), .B2(n_773), .C1(n_774), .C2(n_775), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_122), .Y(n_772) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI22x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_471), .B1(n_472), .B2(n_770), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_130), .A2(n_471), .B1(n_473), .B2(n_770), .Y(n_773) );
OA22x2_ASAP7_75t_L g783 ( .A1(n_130), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_783) );
INVx2_ASAP7_75t_SL g784 ( .A(n_130), .Y(n_784) );
OA22x2_ASAP7_75t_L g790 ( .A1(n_130), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_790) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_396), .Y(n_130) );
NOR2xp67_ASAP7_75t_L g131 ( .A(n_132), .B(n_315), .Y(n_131) );
NAND5xp2_ASAP7_75t_L g132 ( .A(n_133), .B(n_259), .C(n_269), .D(n_286), .E(n_302), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_193), .B1(n_236), .B2(n_240), .Y(n_134) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_167), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g242 ( .A(n_137), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g261 ( .A(n_137), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g282 ( .A(n_137), .B(n_283), .Y(n_282) );
INVx4_ASAP7_75t_L g296 ( .A(n_137), .Y(n_296) );
AND2x2_ASAP7_75t_L g305 ( .A(n_137), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_SL g327 ( .A(n_137), .B(n_244), .Y(n_327) );
BUFx2_ASAP7_75t_L g370 ( .A(n_137), .Y(n_370) );
AND2x2_ASAP7_75t_L g385 ( .A(n_137), .B(n_168), .Y(n_385) );
OR2x2_ASAP7_75t_L g417 ( .A(n_137), .B(n_418), .Y(n_417) );
NOR4xp25_ASAP7_75t_L g466 ( .A(n_137), .B(n_467), .C(n_468), .D(n_469), .Y(n_466) );
OR2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_164), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_148), .B(n_160), .Y(n_138) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
AND2x6_ASAP7_75t_L g158 ( .A(n_142), .B(n_151), .Y(n_158) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g156 ( .A(n_144), .B(n_153), .Y(n_156) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx5_ASAP7_75t_L g159 ( .A(n_146), .Y(n_159) );
AND2x2_ASAP7_75t_L g152 ( .A(n_147), .B(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
BUFx3_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
INVx2_ASAP7_75t_L g192 ( .A(n_151), .Y(n_192) );
AND2x4_ASAP7_75t_L g188 ( .A(n_152), .B(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_158), .B(n_212), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_159), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_159), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_159), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_159), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_159), .A2(n_234), .B(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_159), .A2(n_250), .B(n_251), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_159), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_159), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_159), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_159), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_159), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_159), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_159), .A2(n_555), .B(n_556), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_159), .A2(n_564), .B(n_565), .Y(n_563) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_160), .A2(n_181), .B(n_187), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_160), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_160), .A2(n_482), .B(n_483), .Y(n_481) );
OA21x2_ASAP7_75t_L g561 ( .A1(n_160), .A2(n_562), .B(n_566), .Y(n_561) );
OA21x2_ASAP7_75t_L g606 ( .A1(n_160), .A2(n_562), .B(n_566), .Y(n_606) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_162), .B(n_163), .Y(n_161) );
AND2x4_ASAP7_75t_L g204 ( .A(n_162), .B(n_163), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_165), .A2(n_207), .B(n_208), .Y(n_206) );
BUFx4f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g169 ( .A(n_166), .Y(n_169) );
AOI31xp33_ASAP7_75t_L g334 ( .A1(n_167), .A2(n_335), .A3(n_337), .B(n_339), .Y(n_334) );
INVx2_ASAP7_75t_SL g451 ( .A(n_167), .Y(n_451) );
OR2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_178), .Y(n_167) );
INVx2_ASAP7_75t_L g258 ( .A(n_168), .Y(n_258) );
AND2x2_ASAP7_75t_L g262 ( .A(n_168), .B(n_245), .Y(n_262) );
INVx2_ASAP7_75t_L g285 ( .A(n_168), .Y(n_285) );
AND2x2_ASAP7_75t_L g304 ( .A(n_168), .B(n_244), .Y(n_304) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_176), .Y(n_168) );
INVx4_ASAP7_75t_L g177 ( .A(n_169), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_175), .Y(n_170) );
INVx3_ASAP7_75t_L g218 ( .A(n_177), .Y(n_218) );
AND2x2_ASAP7_75t_L g256 ( .A(n_178), .B(n_257), .Y(n_256) );
BUFx3_ASAP7_75t_L g263 ( .A(n_178), .Y(n_263) );
INVx2_ASAP7_75t_L g281 ( .A(n_178), .Y(n_281) );
AND2x2_ASAP7_75t_L g336 ( .A(n_178), .B(n_296), .Y(n_336) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
AND2x4_ASAP7_75t_L g307 ( .A(n_179), .B(n_180), .Y(n_307) );
AND2x4_ASAP7_75t_L g182 ( .A(n_183), .B(n_186), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
NOR2x1p5_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_226), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_214), .Y(n_194) );
OR2x2_ASAP7_75t_L g236 ( .A(n_195), .B(n_237), .Y(n_236) );
INVx3_ASAP7_75t_L g388 ( .A(n_195), .Y(n_388) );
OR2x2_ASAP7_75t_L g436 ( .A(n_195), .B(n_437), .Y(n_436) );
NAND2x1_ASAP7_75t_L g195 ( .A(n_196), .B(n_205), .Y(n_195) );
OR2x2_ASAP7_75t_SL g227 ( .A(n_196), .B(n_228), .Y(n_227) );
INVx4_ASAP7_75t_L g266 ( .A(n_196), .Y(n_266) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_196), .Y(n_310) );
INVx2_ASAP7_75t_L g318 ( .A(n_196), .Y(n_318) );
OR2x2_ASAP7_75t_L g353 ( .A(n_196), .B(n_216), .Y(n_353) );
AND2x2_ASAP7_75t_L g465 ( .A(n_196), .B(n_320), .Y(n_465) );
AND2x2_ASAP7_75t_L g470 ( .A(n_196), .B(n_229), .Y(n_470) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_204), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_204), .A2(n_231), .B(n_232), .Y(n_230) );
INVx1_ASAP7_75t_SL g490 ( .A(n_204), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_204), .B(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_204), .A2(n_534), .B(n_535), .Y(n_533) );
OR2x2_ASAP7_75t_L g228 ( .A(n_205), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g294 ( .A(n_205), .B(n_215), .Y(n_294) );
OR2x2_ASAP7_75t_L g301 ( .A(n_205), .B(n_266), .Y(n_301) );
NOR2x1_ASAP7_75t_SL g320 ( .A(n_205), .B(n_239), .Y(n_320) );
BUFx2_ASAP7_75t_L g352 ( .A(n_205), .Y(n_352) );
AND2x2_ASAP7_75t_L g361 ( .A(n_205), .B(n_266), .Y(n_361) );
AND2x2_ASAP7_75t_L g394 ( .A(n_205), .B(n_314), .Y(n_394) );
INVx2_ASAP7_75t_SL g403 ( .A(n_205), .Y(n_403) );
AND2x2_ASAP7_75t_L g406 ( .A(n_205), .B(n_216), .Y(n_406) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_213), .Y(n_205) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_214), .B(n_271), .C(n_356), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_214), .B(n_318), .Y(n_421) );
INVxp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_215), .B(n_403), .Y(n_424) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_216), .Y(n_268) );
AND2x2_ASAP7_75t_L g312 ( .A(n_216), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g377 ( .A(n_216), .B(n_378), .Y(n_377) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_225), .Y(n_217) );
AO21x1_ASAP7_75t_SL g239 ( .A1(n_218), .A2(n_219), .B(n_225), .Y(n_239) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_218), .A2(n_522), .B(n_528), .Y(n_521) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_218), .A2(n_522), .B(n_528), .Y(n_543) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_218), .A2(n_552), .B(n_558), .Y(n_551) );
AO21x2_ASAP7_75t_L g576 ( .A1(n_218), .A2(n_552), .B(n_558), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
AND2x4_ASAP7_75t_L g272 ( .A(n_226), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g408 ( .A(n_228), .B(n_353), .Y(n_408) );
AND2x2_ASAP7_75t_L g238 ( .A(n_229), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g276 ( .A(n_229), .Y(n_276) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_229), .Y(n_293) );
INVx2_ASAP7_75t_L g314 ( .A(n_229), .Y(n_314) );
INVx1_ASAP7_75t_L g378 ( .A(n_229), .Y(n_378) );
INVx2_ASAP7_75t_L g460 ( .A(n_236), .Y(n_460) );
OR2x2_ASAP7_75t_L g324 ( .A(n_237), .B(n_301), .Y(n_324) );
INVx2_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g464 ( .A(n_238), .B(n_361), .Y(n_464) );
AND2x2_ASAP7_75t_L g357 ( .A(n_239), .B(n_314), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_254), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_242), .A2(n_371), .B1(n_388), .B2(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g284 ( .A(n_244), .Y(n_284) );
AND2x2_ASAP7_75t_L g338 ( .A(n_244), .B(n_258), .Y(n_338) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_244), .Y(n_365) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_245), .Y(n_333) );
AOI21x1_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_253), .Y(n_245) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_246), .A2(n_501), .B(n_507), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_252), .Y(n_247) );
INVxp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_256), .B(n_370), .Y(n_369) );
OAI32xp33_ASAP7_75t_L g386 ( .A1(n_256), .A2(n_387), .A3(n_389), .B1(n_390), .B2(n_392), .Y(n_386) );
BUFx2_ASAP7_75t_L g271 ( .A(n_257), .Y(n_271) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g413 ( .A(n_258), .B(n_307), .Y(n_413) );
OR4x1_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .C(n_264), .D(n_267), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_260), .A2(n_351), .B1(n_445), .B2(n_446), .Y(n_444) );
INVx2_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_261), .Y(n_453) );
AND2x2_ASAP7_75t_L g295 ( .A(n_262), .B(n_296), .Y(n_295) );
BUFx2_ASAP7_75t_L g375 ( .A(n_262), .Y(n_375) );
INVx1_ASAP7_75t_L g391 ( .A(n_262), .Y(n_391) );
INVx1_ASAP7_75t_L g426 ( .A(n_262), .Y(n_426) );
OR2x2_ASAP7_75t_L g383 ( .A(n_263), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g427 ( .A(n_263), .B(n_428), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_264), .A2(n_301), .B1(n_345), .B2(n_364), .Y(n_366) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g410 ( .A(n_265), .B(n_319), .Y(n_410) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx2_ASAP7_75t_L g277 ( .A(n_266), .Y(n_277) );
NOR2xp67_ASAP7_75t_L g292 ( .A(n_266), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g273 ( .A(n_267), .Y(n_273) );
NAND4xp25_ASAP7_75t_L g400 ( .A(n_267), .B(n_271), .C(n_352), .D(n_364), .Y(n_400) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g437 ( .A(n_268), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_272), .B1(n_274), .B2(n_278), .Y(n_269) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_270), .A2(n_271), .B1(n_421), .B2(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVxp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx3_ASAP7_75t_L g299 ( .A(n_276), .Y(n_299) );
AOI32xp33_ASAP7_75t_L g415 ( .A1(n_276), .A2(n_416), .A3(n_420), .B1(n_425), .B2(n_429), .Y(n_415) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_282), .Y(n_278) );
NOR2xp67_ASAP7_75t_L g321 ( .A(n_279), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g374 ( .A(n_279), .B(n_375), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_279), .A2(n_287), .B1(n_399), .B2(n_404), .C(n_407), .Y(n_398) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g331 ( .A(n_280), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g446 ( .A(n_280), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_281), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g288 ( .A(n_283), .Y(n_288) );
AND2x2_ASAP7_75t_L g306 ( .A(n_283), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_SL g346 ( .A(n_284), .Y(n_346) );
INVx1_ASAP7_75t_L g330 ( .A(n_285), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_289), .B1(n_295), .B2(n_297), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g432 ( .A(n_288), .B(n_362), .Y(n_432) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g372 ( .A(n_291), .Y(n_372) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
AND2x2_ASAP7_75t_L g303 ( .A(n_296), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_296), .B(n_333), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_296), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_296), .B(n_338), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_297), .A2(n_457), .B1(n_458), .B2(n_460), .Y(n_456) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
OR2x2_ASAP7_75t_L g339 ( .A(n_299), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g349 ( .A(n_299), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_299), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_299), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_SL g404 ( .A(n_299), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g380 ( .A(n_301), .B(n_381), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .B(n_308), .Y(n_302) );
INVx1_ASAP7_75t_L g322 ( .A(n_304), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_305), .A2(n_342), .B1(n_349), .B2(n_354), .Y(n_341) );
INVx3_ASAP7_75t_L g344 ( .A(n_307), .Y(n_344) );
INVx2_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
OAI32xp33_ASAP7_75t_SL g399 ( .A1(n_310), .A2(n_370), .A3(n_400), .B1(n_401), .B2(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g319 ( .A(n_313), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND4xp25_ASAP7_75t_SL g315 ( .A(n_316), .B(n_341), .C(n_358), .D(n_373), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_321), .B1(n_323), .B2(n_325), .C(n_334), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g356 ( .A(n_318), .Y(n_356) );
AND2x2_ASAP7_75t_L g405 ( .A(n_318), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_318), .B(n_357), .Y(n_443) );
AND2x2_ASAP7_75t_L g454 ( .A(n_318), .B(n_377), .Y(n_454) );
INVx2_ASAP7_75t_L g340 ( .A(n_320), .Y(n_340) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B(n_331), .Y(n_325) );
AND2x2_ASAP7_75t_L g457 ( .A(n_326), .B(n_328), .Y(n_457) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_327), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g434 ( .A(n_332), .Y(n_434) );
INVx1_ASAP7_75t_L g419 ( .A(n_333), .Y(n_419) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_336), .B(n_391), .Y(n_390) );
NOR2x1_ASAP7_75t_L g348 ( .A(n_337), .B(n_344), .Y(n_348) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g447 ( .A(n_338), .Y(n_447) );
INVx1_ASAP7_75t_L g429 ( .A(n_340), .Y(n_429) );
OR2x2_ASAP7_75t_L g445 ( .A(n_340), .B(n_356), .Y(n_445) );
NAND2xp33_ASAP7_75t_SL g342 ( .A(n_343), .B(n_347), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx2_ASAP7_75t_L g362 ( .A(n_344), .Y(n_362) );
AND2x2_ASAP7_75t_L g367 ( .A(n_344), .B(n_357), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_344), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g441 ( .A(n_345), .Y(n_441) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_350), .A2(n_431), .B1(n_433), .B2(n_435), .Y(n_430) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g395 ( .A(n_353), .Y(n_395) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g381 ( .A(n_357), .Y(n_381) );
AOI322xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .A3(n_363), .B1(n_366), .B2(n_367), .C1(n_368), .C2(n_371), .Y(n_358) );
OAI21xp5_ASAP7_75t_SL g409 ( .A1(n_359), .A2(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g376 ( .A(n_361), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g433 ( .A(n_362), .B(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_369), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g389 ( .A(n_370), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_370), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B1(n_379), .B2(n_382), .C(n_386), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_375), .A2(n_462), .B1(n_464), .B2(n_465), .C(n_466), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_377), .B(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_L g428 ( .A(n_378), .Y(n_428) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_382), .A2(n_453), .B(n_454), .Y(n_452) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp33_ASAP7_75t_SL g462 ( .A(n_391), .B(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
NOR4xp75_ASAP7_75t_L g396 ( .A(n_397), .B(n_414), .C(n_438), .D(n_455), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_409), .Y(n_397) );
INVx1_ASAP7_75t_L g468 ( .A(n_406), .Y(n_468) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g440 ( .A(n_413), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g467 ( .A(n_413), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_415), .B(n_430), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_SL g463 ( .A(n_434), .Y(n_463) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND3x1_ASAP7_75t_L g438 ( .A(n_439), .B(n_448), .C(n_452), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_442), .B(n_444), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_461), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_655), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_610), .C(n_639), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_476), .B(n_583), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_508), .B1(n_529), .B2(n_540), .C(n_544), .Y(n_476) );
INVx3_ASAP7_75t_SL g700 ( .A(n_477), .Y(n_700) );
AND2x2_ASAP7_75t_SL g477 ( .A(n_478), .B(n_487), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g546 ( .A(n_478), .B(n_499), .Y(n_546) );
INVx4_ASAP7_75t_L g581 ( .A(n_478), .Y(n_581) );
AND2x2_ASAP7_75t_L g603 ( .A(n_478), .B(n_500), .Y(n_603) );
AND2x2_ASAP7_75t_L g609 ( .A(n_478), .B(n_548), .Y(n_609) );
INVx5_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g578 ( .A(n_479), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_479), .B(n_499), .Y(n_654) );
AND2x2_ASAP7_75t_L g659 ( .A(n_479), .B(n_500), .Y(n_659) );
AND2x2_ASAP7_75t_L g671 ( .A(n_479), .B(n_532), .Y(n_671) );
NOR2x1_ASAP7_75t_SL g710 ( .A(n_479), .B(n_548), .Y(n_710) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g539 ( .A(n_487), .Y(n_539) );
AND2x2_ASAP7_75t_L g643 ( .A(n_487), .B(n_592), .Y(n_643) );
AND2x2_ASAP7_75t_L g740 ( .A(n_487), .B(n_671), .Y(n_740) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_499), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g572 ( .A(n_489), .Y(n_572) );
INVx2_ASAP7_75t_L g594 ( .A(n_489), .Y(n_594) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B(n_497), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_490), .B(n_498), .Y(n_497) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_490), .A2(n_491), .B(n_497), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_496), .Y(n_491) );
AND2x2_ASAP7_75t_L g569 ( .A(n_499), .B(n_531), .Y(n_569) );
INVx2_ASAP7_75t_L g573 ( .A(n_499), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_499), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g672 ( .A(n_499), .B(n_637), .Y(n_672) );
OR2x2_ASAP7_75t_L g719 ( .A(n_499), .B(n_532), .Y(n_719) );
INVx4_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_500), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_506), .Y(n_501) );
AND2x2_ASAP7_75t_L g716 ( .A(n_508), .B(n_597), .Y(n_716) );
AND2x2_ASAP7_75t_L g766 ( .A(n_508), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g642 ( .A(n_509), .B(n_586), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
AND2x2_ASAP7_75t_L g575 ( .A(n_510), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g605 ( .A(n_510), .B(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g626 ( .A(n_510), .B(n_606), .Y(n_626) );
AND2x4_ASAP7_75t_L g661 ( .A(n_510), .B(n_649), .Y(n_661) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g542 ( .A(n_511), .Y(n_542) );
OAI21x1_ASAP7_75t_SL g511 ( .A1(n_512), .A2(n_514), .B(n_518), .Y(n_511) );
INVx1_ASAP7_75t_L g519 ( .A(n_513), .Y(n_519) );
AND2x2_ASAP7_75t_L g588 ( .A(n_520), .B(n_541), .Y(n_588) );
AND2x2_ASAP7_75t_L g674 ( .A(n_520), .B(n_606), .Y(n_674) );
AND2x2_ASAP7_75t_L g685 ( .A(n_520), .B(n_550), .Y(n_685) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g549 ( .A(n_521), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g616 ( .A(n_521), .B(n_551), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_523), .B(n_527), .Y(n_522) );
INVx2_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_539), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_531), .B(n_581), .Y(n_638) );
AND2x2_ASAP7_75t_L g682 ( .A(n_531), .B(n_548), .Y(n_682) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_532), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g592 ( .A(n_532), .Y(n_592) );
BUFx3_ASAP7_75t_L g601 ( .A(n_532), .Y(n_601) );
AND2x2_ASAP7_75t_L g624 ( .A(n_532), .B(n_594), .Y(n_624) );
OAI322xp33_ASAP7_75t_L g544 ( .A1(n_539), .A2(n_545), .A3(n_549), .B1(n_559), .B2(n_567), .C1(n_574), .C2(n_579), .Y(n_544) );
INVx1_ASAP7_75t_L g705 ( .A(n_539), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_540), .B(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g618 ( .A(n_540), .B(n_560), .Y(n_618) );
INVx2_ASAP7_75t_L g663 ( .A(n_540), .Y(n_663) );
AND2x2_ASAP7_75t_L g679 ( .A(n_540), .B(n_621), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_540), .B(n_697), .Y(n_727) );
AND2x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x2_ASAP7_75t_SL g630 ( .A(n_541), .B(n_606), .Y(n_630) );
OR2x2_ASAP7_75t_L g651 ( .A(n_541), .B(n_568), .Y(n_651) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g623 ( .A(n_542), .Y(n_623) );
INVx2_ASAP7_75t_L g568 ( .A(n_543), .Y(n_568) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_543), .Y(n_570) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g613 ( .A(n_546), .Y(n_613) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_547), .Y(n_633) );
INVx1_ASAP7_75t_L g731 ( .A(n_547), .Y(n_731) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_547), .Y(n_746) );
NAND2x1_ASAP7_75t_L g756 ( .A(n_549), .B(n_560), .Y(n_756) );
INVx1_ASAP7_75t_L g763 ( .A(n_549), .Y(n_763) );
BUFx2_ASAP7_75t_L g597 ( .A(n_550), .Y(n_597) );
AND2x2_ASAP7_75t_L g673 ( .A(n_550), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx3_ASAP7_75t_L g582 ( .A(n_551), .Y(n_582) );
INVxp67_ASAP7_75t_L g586 ( .A(n_551), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_559), .B(n_575), .C(n_577), .Y(n_574) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_SL g595 ( .A(n_560), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_560), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g747 ( .A(n_560), .B(n_696), .Y(n_747) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g649 ( .A(n_561), .Y(n_649) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_561), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_567) );
AND2x4_ASAP7_75t_SL g696 ( .A(n_568), .B(n_576), .Y(n_696) );
AND2x2_ASAP7_75t_L g709 ( .A(n_569), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_570), .Y(n_711) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx2_ASAP7_75t_L g668 ( .A(n_572), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_572), .B(n_581), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_573), .B(n_591), .Y(n_590) );
AND3x2_ASAP7_75t_L g608 ( .A(n_573), .B(n_601), .C(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g632 ( .A(n_573), .Y(n_632) );
AND2x2_ASAP7_75t_L g745 ( .A(n_573), .B(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g621 ( .A(n_576), .Y(n_621) );
INVx1_ASAP7_75t_L g699 ( .A(n_576), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_577), .B(n_600), .Y(n_738) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_578), .B(n_682), .Y(n_687) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g678 ( .A(n_581), .B(n_624), .Y(n_678) );
INVx1_ASAP7_75t_SL g629 ( .A(n_582), .Y(n_629) );
AND2x2_ASAP7_75t_L g737 ( .A(n_582), .B(n_649), .Y(n_737) );
AND2x2_ASAP7_75t_L g758 ( .A(n_582), .B(n_630), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_589), .B1(n_595), .B2(n_598), .C(n_604), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g750 ( .A(n_586), .Y(n_750) );
AOI21xp33_ASAP7_75t_SL g604 ( .A1(n_587), .A2(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g596 ( .A(n_588), .B(n_597), .Y(n_596) );
AOI222xp33_ASAP7_75t_L g619 ( .A1(n_588), .A2(n_620), .B1(n_622), .B2(n_627), .C1(n_631), .C2(n_634), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_588), .B(n_737), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_589), .A2(n_618), .B1(n_641), .B2(n_643), .Y(n_640) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g625 ( .A(n_592), .Y(n_625) );
AND2x2_ASAP7_75t_L g744 ( .A(n_592), .B(n_710), .Y(n_744) );
OAI32xp33_ASAP7_75t_L g748 ( .A1(n_592), .A2(n_617), .A3(n_669), .B1(n_677), .B2(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g753 ( .A(n_592), .B(n_603), .Y(n_753) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g637 ( .A(n_594), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g644 ( .A1(n_595), .A2(n_645), .B(n_652), .Y(n_644) );
INVx1_ASAP7_75t_L g708 ( .A(n_597), .Y(n_708) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
AND2x2_ASAP7_75t_L g612 ( .A(n_600), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g620 ( .A(n_603), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g693 ( .A(n_603), .B(n_624), .Y(n_693) );
INVx1_ASAP7_75t_SL g764 ( .A(n_605), .Y(n_764) );
AND2x2_ASAP7_75t_L g698 ( .A(n_606), .B(n_699), .Y(n_698) );
OAI222xp33_ASAP7_75t_L g751 ( .A1(n_607), .A2(n_660), .B1(n_739), .B2(n_752), .C1(n_754), .C2(n_756), .Y(n_751) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g724 ( .A(n_609), .B(n_725), .Y(n_724) );
OAI21xp33_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_614), .B(n_619), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_613), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g692 ( .A(n_615), .Y(n_692) );
INVx1_ASAP7_75t_L g660 ( .A(n_616), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_616), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g714 ( .A(n_621), .Y(n_714) );
AO22x1_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_625), .B2(n_626), .Y(n_622) );
OAI322xp33_ASAP7_75t_L g734 ( .A1(n_623), .A2(n_684), .A3(n_687), .B1(n_735), .B2(n_736), .C1(n_738), .C2(n_739), .Y(n_734) );
AND2x2_ASAP7_75t_SL g658 ( .A(n_624), .B(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g653 ( .A(n_625), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_626), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g755 ( .A(n_626), .B(n_685), .Y(n_755) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g735 ( .A(n_629), .Y(n_735) );
INVx1_ASAP7_75t_SL g664 ( .A(n_630), .Y(n_664) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
OR2x2_ASAP7_75t_L g666 ( .A(n_638), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g704 ( .A(n_638), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_644), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_650), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g677 ( .A(n_648), .B(n_663), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_648), .B(n_685), .Y(n_684) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g707 ( .A(n_651), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2x1_ASAP7_75t_L g655 ( .A(n_656), .B(n_720), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_657), .B(n_675), .C(n_688), .D(n_701), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .A3(n_661), .B1(n_662), .B2(n_665), .C1(n_670), .C2(n_673), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g757 ( .A1(n_658), .A2(n_758), .B(n_759), .C(n_762), .Y(n_757) );
AND2x2_ASAP7_75t_L g769 ( .A(n_659), .B(n_746), .Y(n_769) );
INVx1_ASAP7_75t_L g691 ( .A(n_661), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_661), .B(n_696), .Y(n_733) );
NAND2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_669), .B(n_682), .Y(n_749) );
AND2x4_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B1(n_679), .B2(n_680), .C1(n_683), .C2(n_686), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_678), .A2(n_689), .B1(n_692), .B2(n_693), .C(n_694), .Y(n_688) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI21xp33_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_697), .B(n_700), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_706), .B1(n_709), .B2(n_711), .C(n_712), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g761 ( .A(n_710), .Y(n_761) );
AOI21xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B(n_717), .Y(n_712) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx2_ASAP7_75t_L g725 ( .A(n_719), .Y(n_725) );
OR2x2_ASAP7_75t_L g760 ( .A(n_719), .B(n_761), .Y(n_760) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_741), .C(n_757), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_734), .Y(n_721) );
OAI21xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_726), .B(n_728), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_732), .Y(n_728) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_747), .B1(n_748), .B2(n_750), .C(n_751), .Y(n_741) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NOR2x1_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_756), .B(n_760), .Y(n_759) );
O2A1O1Ixp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B(n_765), .C(n_768), .Y(n_762) );
INVxp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
CKINVDCx11_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
INVx3_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
NOR2x1_ASAP7_75t_R g791 ( .A(n_780), .B(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_797), .Y(n_793) );
CKINVDCx11_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
endmodule