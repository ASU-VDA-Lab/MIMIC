module fake_jpeg_25209_n_169 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_38),
.Y(n_59)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_50),
.B1(n_27),
.B2(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_28),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_20),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_33),
.C(n_32),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_21),
.B1(n_20),
.B2(n_29),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_37),
.B1(n_32),
.B2(n_24),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_57),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_29),
.B1(n_27),
.B2(n_31),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_66),
.Y(n_90)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_68),
.Y(n_79)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_31),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_74),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_59),
.C(n_33),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_42),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_57),
.B1(n_15),
.B2(n_30),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_56),
.B1(n_49),
.B2(n_53),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_80),
.B1(n_87),
.B2(n_88),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_56),
.B1(n_37),
.B2(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_57),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_66),
.B1(n_73),
.B2(n_63),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_74),
.B1(n_72),
.B2(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_15),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_60),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_24),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_98),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_103),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_108),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_22),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_76),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_76),
.Y(n_124)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_114),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_79),
.B1(n_91),
.B2(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_119),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_83),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_86),
.Y(n_130)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_109),
.C(n_103),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_130),
.C(n_133),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_101),
.B(n_105),
.C(n_108),
.D(n_96),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_117),
.B(n_118),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_96),
.C(n_92),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_81),
.B1(n_62),
.B2(n_76),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_127),
.B1(n_38),
.B2(n_137),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_116),
.B(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_136),
.Y(n_145)
);

AO221x1_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_52),
.B1(n_54),
.B2(n_43),
.C(n_3),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_113),
.C(n_123),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_143),
.C(n_54),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_146),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_144),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_118),
.C(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_0),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_7),
.B(n_14),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_151),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_131),
.B1(n_135),
.B2(n_129),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_149),
.A2(n_150),
.B1(n_147),
.B2(n_152),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_13),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_12),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_157),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_138),
.B(n_13),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_1),
.B(n_2),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_151),
.B(n_8),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_8),
.C(n_7),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_161),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_4),
.B(n_5),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_6),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_164),
.B(n_6),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_166),
.Y(n_169)
);


endmodule