module real_jpeg_5151_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_188;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_1),
.A2(n_171),
.B1(n_172),
.B2(n_174),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_1),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_2),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_23),
.B1(n_51),
.B2(n_54),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_23),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_2),
.A2(n_23),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_2),
.A2(n_144),
.B(n_147),
.C(n_150),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_2),
.B(n_26),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_2),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_2),
.B(n_97),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_2),
.B(n_213),
.C(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_2),
.B(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_2),
.B(n_73),
.C(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_3),
.A2(n_24),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_3),
.A2(n_44),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_44),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_3),
.A2(n_44),
.B1(n_116),
.B2(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_6),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_6),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_7),
.Y(n_149)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_10),
.Y(n_213)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_190),
.B1(n_269),
.B2(n_270),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_13),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_188),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_160),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_15),
.B(n_160),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_118),
.C(n_151),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_16),
.B(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_46),
.B2(n_47),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_18),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_18),
.B(n_49),
.C(n_88),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_25),
.B1(n_41),
.B2(n_45),
.Y(n_18)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_19),
.A2(n_25),
.B1(n_41),
.B2(n_45),
.Y(n_163)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_23),
.A2(n_51),
.B(n_148),
.Y(n_147)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_24),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_26)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_88),
.B2(n_117),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_48),
.A2(n_49),
.B1(n_178),
.B2(n_179),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_48),
.B(n_178),
.C(n_235),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_57),
.B1(n_71),
.B2(n_82),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_50),
.A2(n_57),
.B1(n_71),
.B2(n_82),
.Y(n_153)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2x1_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_71),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_68),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_71),
.Y(n_224)
);

AOI22x1_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_75),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_87),
.Y(n_240)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_89),
.B(n_108),
.Y(n_180)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_89),
.Y(n_228)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_96),
.A2(n_107),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_97),
.B(n_182),
.Y(n_181)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_102),
.B2(n_105),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_110),
.B1(n_112),
.B2(n_115),
.Y(n_109)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_118),
.A2(n_119),
.B1(n_151),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_142),
.B2(n_143),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_143),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_120),
.A2(n_121),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_121),
.B(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_121),
.B(n_203),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_121),
.B(n_223),
.C(n_226),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_129),
.B1(n_135),
.B2(n_138),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_129),
.B1(n_138),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_128),
.Y(n_247)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_131),
.Y(n_216)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_138),
.B(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_151),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_158),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_153),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_152),
.A2(n_153),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_154),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_206),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_259)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_198),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_163),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_187),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_178),
.B1(n_179),
.B2(n_186),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B(n_175),
.Y(n_168)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_176),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_178),
.A2(n_179),
.B1(n_207),
.B2(n_217),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_217),
.Y(n_230)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_190),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_263),
.B(n_268),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_251),
.B(n_262),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_232),
.B(n_250),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_219),
.B(n_231),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_205),
.B(n_218),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_202),
.B(n_204),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_230),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_230),
.Y(n_231)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_229),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_225),
.A2(n_226),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_254),
.C(n_256),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_234),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_249),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_243),
.B2(n_248),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_248),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_261),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_261),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_256),
.B1(n_257),
.B2(n_260),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);


endmodule