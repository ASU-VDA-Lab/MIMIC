module fake_jpeg_31946_n_122 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_122);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_56),
.Y(n_67)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_20),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_2),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_61),
.B(n_62),
.C(n_48),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_44),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_59),
.B(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_5),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_72),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_51),
.B1(n_46),
.B2(n_41),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_46),
.B1(n_41),
.B2(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_4),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_62),
.B(n_52),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_83),
.B(n_90),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_86),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_58),
.B1(n_44),
.B2(n_23),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_21),
.B1(n_40),
.B2(n_39),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_19),
.B1(n_38),
.B2(n_36),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_16),
.B1(n_35),
.B2(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_88),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_58),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_11),
.C(n_12),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_5),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_15),
.B1(n_30),
.B2(n_29),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_65),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_13),
.B1(n_28),
.B2(n_27),
.Y(n_90)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_9),
.B1(n_10),
.B2(n_25),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_6),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_100),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_101),
.B1(n_10),
.B2(n_26),
.Y(n_112)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_18),
.CI(n_32),
.CON(n_100),
.SN(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_8),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_102),
.B(n_103),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_64),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_9),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_95),
.B1(n_98),
.B2(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_114),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_103),
.B(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_108),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_104),
.C(n_111),
.Y(n_118)
);

INVxp67_ASAP7_75t_SL g119 ( 
.A(n_118),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_117),
.A3(n_109),
.B1(n_114),
.B2(n_106),
.C1(n_94),
.C2(n_107),
.Y(n_121)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_93),
.C(n_92),
.Y(n_122)
);


endmodule