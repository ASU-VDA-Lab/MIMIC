module real_jpeg_23720_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_215;
wire n_300;
wire n_221;
wire n_249;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_1),
.B(n_43),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_1),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_1),
.B(n_31),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_1),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_2),
.B(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_2),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_2),
.B(n_31),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_2),
.B(n_137),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_2),
.B(n_36),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_3),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_3),
.B(n_51),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_3),
.B(n_45),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_3),
.B(n_43),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_3),
.B(n_31),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_3),
.B(n_36),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_3),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_3),
.B(n_25),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_4),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_4),
.B(n_43),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_4),
.B(n_25),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_45),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_4),
.B(n_17),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_4),
.B(n_36),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_4),
.B(n_31),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx8_ASAP7_75t_SL g53 ( 
.A(n_7),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_9),
.B(n_36),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_9),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_10),
.B(n_51),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_10),
.B(n_25),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_10),
.B(n_31),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_10),
.B(n_45),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_10),
.B(n_36),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_10),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_10),
.B(n_43),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_13),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_13),
.B(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_13),
.B(n_43),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_13),
.B(n_25),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_13),
.B(n_36),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_13),
.B(n_31),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_13),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_13),
.B(n_45),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_14),
.B(n_36),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_14),
.B(n_31),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_14),
.B(n_137),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_16),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_16),
.B(n_43),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_16),
.B(n_25),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_16),
.B(n_45),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_16),
.B(n_36),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_16),
.B(n_51),
.Y(n_247)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_17),
.Y(n_115)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_17),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_156),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_91),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_38),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_31),
.Y(n_219)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_38),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_33),
.B(n_57),
.C(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_35),
.B(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_47),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.C(n_44),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_42),
.CI(n_44),
.CON(n_69),
.SN(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_47),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.CI(n_50),
.CON(n_47),
.SN(n_47)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_70),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_63),
.C(n_69),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_56),
.B(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_61),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_64),
.C(n_65),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_69),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_66),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_69),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_84),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_82),
.C(n_83),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_73),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.C(n_79),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_79),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_82),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_83),
.B1(n_89),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_105),
.C(n_109),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.C(n_101),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_93),
.B(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_95),
.B(n_101),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.C(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_98),
.B(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_122),
.C(n_123),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.C(n_120),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_123),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_131),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_302)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_131),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_144),
.C(n_146),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_132),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.C(n_140),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_133),
.B(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_135),
.A2(n_136),
.B(n_139),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_135),
.B(n_140),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.C(n_143),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_141),
.B(n_142),
.CI(n_143),
.CON(n_261),
.SN(n_261)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_144),
.B(n_146),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.C(n_154),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_147),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_151),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_148),
.B(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_150),
.B(n_151),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_300),
.C(n_301),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_290),
.C(n_291),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_275),
.C(n_276),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_254),
.C(n_255),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_229),
.C(n_230),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_189),
.C(n_201),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_176),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_171),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_171),
.C(n_176),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_166),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_172),
.B(n_174),
.C(n_175),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_177),
.B(n_183),
.C(n_184),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_185),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_188),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_200),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_194),
.B1(n_200),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_225),
.C(n_226),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_210),
.C(n_216),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_208),
.C(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.C(n_220),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_244),
.C(n_253),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_238),
.C(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_234),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_237),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_239),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.CI(n_242),
.CON(n_239),
.SN(n_239)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_253),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_251),
.B2(n_252),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_247),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_250),
.C(n_252),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_267),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_259),
.C(n_267),
.Y(n_275)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_263),
.C(n_266),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_261),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_271),
.C(n_273),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_270),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_271),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_285),
.B2(n_289),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_286),
.C(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_281),
.C(n_283),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_298),
.B2(n_299),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_292),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_296),
.C(n_298),
.Y(n_300)
);


endmodule