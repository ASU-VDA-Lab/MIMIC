module fake_jpeg_20950_n_315 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_37),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_29),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_19),
.B1(n_34),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_72),
.B1(n_26),
.B2(n_33),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_22),
.B1(n_19),
.B2(n_33),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_58),
.B1(n_35),
.B2(n_30),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_19),
.B1(n_20),
.B2(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_20),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_65),
.B(n_66),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_28),
.C(n_18),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_74),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_31),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_29),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_19),
.B1(n_37),
.B2(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_38),
.A2(n_26),
.B1(n_33),
.B2(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_21),
.B1(n_27),
.B2(n_25),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_80),
.A2(n_84),
.B(n_92),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_23),
.B1(n_37),
.B2(n_18),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_81),
.A2(n_83),
.B1(n_85),
.B2(n_91),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_42),
.B(n_1),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_48),
.B1(n_21),
.B2(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_86),
.B(n_12),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_90),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_88),
.A2(n_102),
.B(n_95),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_48),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_115),
.C(n_50),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_26),
.B1(n_32),
.B2(n_21),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_0),
.B(n_1),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_25),
.B1(n_27),
.B2(n_32),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_107),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_25),
.B1(n_46),
.B2(n_30),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_35),
.B1(n_46),
.B2(n_28),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx5_ASAP7_75t_SL g141 ( 
.A(n_97),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_35),
.B1(n_36),
.B2(n_24),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_109),
.B1(n_62),
.B2(n_69),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_36),
.B(n_24),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_55),
.A2(n_36),
.B1(n_9),
.B2(n_15),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_54),
.A2(n_46),
.B1(n_7),
.B2(n_8),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_0),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

AO22x2_ASAP7_75t_SL g114 ( 
.A1(n_63),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_2),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_120),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_61),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_59),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_122),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_84),
.B1(n_102),
.B2(n_105),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_135),
.B1(n_139),
.B2(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_133),
.B(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_71),
.B1(n_60),
.B2(n_69),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_138),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_83),
.B(n_89),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_147),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_85),
.A2(n_52),
.B1(n_76),
.B2(n_50),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_114),
.B1(n_115),
.B2(n_103),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_76),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_149),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_8),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_150),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_100),
.C(n_89),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_164),
.C(n_169),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_94),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_171),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_129),
.B1(n_123),
.B2(n_119),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_153),
.A2(n_156),
.B1(n_173),
.B2(n_50),
.Y(n_204)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_166),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_52),
.B1(n_111),
.B2(n_114),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_114),
.B1(n_80),
.B2(n_91),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_177),
.B1(n_136),
.B2(n_138),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_143),
.B(n_130),
.C(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_137),
.Y(n_197)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_140),
.C(n_145),
.Y(n_164)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_111),
.C(n_92),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_116),
.B(n_78),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_115),
.C(n_96),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_146),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_141),
.A2(n_123),
.B1(n_119),
.B2(n_144),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_132),
.Y(n_174)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_93),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_175),
.B(n_180),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_93),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_186),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_142),
.B(n_125),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_185),
.A2(n_193),
.B(n_194),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_181),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_190),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_118),
.C(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_125),
.B(n_136),
.Y(n_193)
);

AND2x4_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_164),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_168),
.B1(n_159),
.B2(n_174),
.Y(n_224)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_207),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_200),
.B(n_208),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_124),
.B1(n_150),
.B2(n_127),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_198),
.A2(n_155),
.B1(n_170),
.B2(n_154),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_182),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_104),
.B(n_97),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_178),
.A2(n_127),
.B1(n_134),
.B2(n_79),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_203),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_167),
.A2(n_161),
.B1(n_151),
.B2(n_169),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_163),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_161),
.A2(n_93),
.B1(n_50),
.B2(n_4),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_211),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_182),
.B(n_7),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_176),
.A2(n_110),
.B(n_3),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_210),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_2),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_224),
.B1(n_236),
.B2(n_205),
.Y(n_243)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_225),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_218),
.B(n_212),
.Y(n_251)
);

XOR2x1_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_176),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_219),
.A2(n_231),
.B(n_200),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_221),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_170),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_154),
.C(n_168),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_203),
.C(n_208),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_191),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_210),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_212),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_159),
.B1(n_174),
.B2(n_166),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_198),
.B1(n_211),
.B2(n_209),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_163),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_222),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_195),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_185),
.B(n_197),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_241),
.B(n_235),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_226),
.B(n_231),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_242),
.A2(n_227),
.B(n_189),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_244),
.B1(n_250),
.B2(n_255),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_194),
.B1(n_187),
.B2(n_183),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_248),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_213),
.A2(n_219),
.B1(n_229),
.B2(n_194),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_213),
.C(n_221),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_184),
.B1(n_202),
.B2(n_192),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_220),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_215),
.A2(n_189),
.B1(n_206),
.B2(n_196),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_234),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_258),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_260),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_236),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_263),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_229),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_225),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_266),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_217),
.C(n_223),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g269 ( 
.A(n_239),
.B(n_241),
.CI(n_244),
.CON(n_269),
.SN(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_259),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_233),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_237),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_280),
.B(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_274),
.B(n_279),
.Y(n_286)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_243),
.B1(n_255),
.B2(n_245),
.Y(n_279)
);

XOR2x2_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_249),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_257),
.A2(n_245),
.B1(n_246),
.B2(n_238),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_283),
.Y(n_292)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

NAND4xp25_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_248),
.C(n_216),
.D(n_6),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_285),
.A2(n_276),
.B(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_284),
.Y(n_301)
);

A2O1A1O1Ixp25_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_261),
.B(n_264),
.C(n_266),
.D(n_260),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_289),
.A2(n_278),
.B(n_282),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_258),
.C(n_256),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_293),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_268),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_284),
.Y(n_300)
);

NAND3xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_289),
.C(n_293),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_281),
.Y(n_297)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_257),
.B1(n_272),
.B2(n_263),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_291),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_305),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_304),
.A2(n_296),
.B1(n_297),
.B2(n_301),
.Y(n_308)
);

OAI211xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_275),
.B(n_5),
.C(n_6),
.Y(n_305)
);

OAI21x1_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_309),
.B(n_5),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_306),
.A2(n_305),
.B1(n_303),
.B2(n_275),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_311),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_309),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_307),
.Y(n_313)
);

OAI221xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_4),
.B1(n_10),
.B2(n_13),
.C(n_311),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_13),
.Y(n_315)
);


endmodule