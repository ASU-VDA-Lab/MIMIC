module fake_jpeg_30893_n_517 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_61),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_46),
.Y(n_69)
);

INVx5_ASAP7_75t_SL g104 ( 
.A(n_69),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_24),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx5_ASAP7_75t_SL g134 ( 
.A(n_84),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_94),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_96),
.Y(n_116)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

BUFx24_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_95),
.B(n_97),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_18),
.B(n_31),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_98),
.B(n_99),
.Y(n_147)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_33),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_49),
.B1(n_36),
.B2(n_35),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_102),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_29),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_33),
.B1(n_50),
.B2(n_28),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_119),
.A2(n_135),
.B1(n_142),
.B2(n_78),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_31),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_123),
.B(n_144),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_54),
.A2(n_40),
.B1(n_38),
.B2(n_33),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_125),
.A2(n_127),
.B1(n_128),
.B2(n_137),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_56),
.A2(n_38),
.B1(n_20),
.B2(n_43),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_58),
.A2(n_38),
.B1(n_20),
.B2(n_43),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_82),
.A2(n_49),
.B1(n_36),
.B2(n_35),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_129),
.A2(n_64),
.B1(n_55),
.B2(n_60),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_68),
.A2(n_76),
.B1(n_38),
.B2(n_98),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_95),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_139),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_61),
.A2(n_21),
.B1(n_37),
.B2(n_25),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_94),
.A2(n_20),
.B1(n_44),
.B2(n_42),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_141),
.A2(n_145),
.B1(n_134),
.B2(n_107),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_87),
.A2(n_101),
.B1(n_96),
.B2(n_89),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_69),
.B(n_26),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_94),
.A2(n_47),
.B1(n_44),
.B2(n_42),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_92),
.B(n_30),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_70),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_47),
.C(n_32),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_37),
.C(n_92),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_161),
.B(n_163),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_32),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_172),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_106),
.B(n_30),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_166),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_167),
.B(n_175),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_154),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_181),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_170),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_171),
.B(n_174),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_29),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_91),
.B1(n_80),
.B2(n_73),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_111),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_176),
.B(n_186),
.Y(n_251)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_178),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_117),
.B(n_90),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_194),
.Y(n_218)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_112),
.B(n_70),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_121),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_182),
.B(n_184),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_183),
.A2(n_207),
.B1(n_128),
.B2(n_127),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_143),
.B(n_16),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_118),
.B(n_90),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_189),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_104),
.B(n_53),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_125),
.A2(n_72),
.B1(n_66),
.B2(n_53),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_107),
.B1(n_134),
.B2(n_126),
.Y(n_227)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_133),
.Y(n_192)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_0),
.Y(n_194)
);

INVx4_ASAP7_75t_SL g195 ( 
.A(n_104),
.Y(n_195)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_109),
.B(n_0),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_159),
.B(n_0),
.Y(n_197)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_105),
.Y(n_199)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_1),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_201),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_113),
.B(n_160),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_202),
.Y(n_231)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_120),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_204),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_1),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_206),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_155),
.B(n_1),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_150),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_113),
.B(n_2),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_208),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_115),
.B(n_124),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_213),
.Y(n_244)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_145),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_124),
.B(n_3),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_141),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_4),
.Y(n_256)
);

OR2x2_ASAP7_75t_SL g215 ( 
.A(n_130),
.B(n_137),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_215),
.A2(n_103),
.B1(n_131),
.B2(n_152),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_227),
.A2(n_174),
.B1(n_195),
.B2(n_198),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_228),
.B(n_248),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_110),
.B1(n_158),
.B2(n_136),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_233),
.A2(n_235),
.B1(n_245),
.B2(n_227),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_110),
.B1(n_158),
.B2(n_136),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_177),
.A2(n_131),
.B1(n_126),
.B2(n_132),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_237),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_187),
.A2(n_152),
.B1(n_130),
.B2(n_132),
.Y(n_245)
);

OAI32xp33_ASAP7_75t_L g254 ( 
.A1(n_164),
.A2(n_103),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_255),
.Y(n_272)
);

OAI32xp33_ASAP7_75t_L g255 ( 
.A1(n_161),
.A2(n_13),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_256),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_215),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

BUFx6f_ASAP7_75t_SL g259 ( 
.A(n_195),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_262),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_162),
.C(n_171),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_265),
.C(n_268),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_179),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_266),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_217),
.B(n_176),
.C(n_198),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_172),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_267),
.A2(n_270),
.B1(n_278),
.B2(n_228),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_194),
.C(n_182),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_269),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_261),
.A2(n_183),
.B1(n_184),
.B2(n_210),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_271),
.B(n_274),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_205),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_273),
.B(n_279),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_216),
.B(n_163),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_275),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_231),
.B(n_173),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_294),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_226),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_218),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_281),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_223),
.B(n_206),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_213),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_283),
.B(n_289),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_211),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_284),
.B(n_292),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_261),
.A2(n_191),
.B(n_207),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_286),
.A2(n_287),
.B(n_248),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_249),
.A2(n_170),
.B(n_178),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_288),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_180),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_259),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_290),
.Y(n_304)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_251),
.B(n_192),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_258),
.B(n_249),
.Y(n_293)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_293),
.B(n_263),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_256),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_230),
.Y(n_296)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_249),
.B(n_166),
.C(n_200),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_245),
.C(n_233),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_220),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_234),
.Y(n_319)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_299),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_225),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_300),
.Y(n_305)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_230),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_302),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_279),
.B(n_236),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_308),
.B(n_334),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_310),
.A2(n_313),
.B(n_322),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_312),
.A2(n_281),
.B1(n_273),
.B2(n_265),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_285),
.A2(n_241),
.B1(n_252),
.B2(n_246),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_318),
.B(n_337),
.C(n_338),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_319),
.B(n_327),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_293),
.A2(n_254),
.B(n_255),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_328),
.Y(n_350)
);

OAI32xp33_ASAP7_75t_L g326 ( 
.A1(n_272),
.A2(n_235),
.A3(n_221),
.B1(n_193),
.B2(n_190),
.Y(n_326)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_292),
.Y(n_327)
);

AO22x1_ASAP7_75t_SL g328 ( 
.A1(n_301),
.A2(n_219),
.B1(n_232),
.B2(n_240),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_272),
.A2(n_294),
.B1(n_283),
.B2(n_301),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_329),
.A2(n_331),
.B1(n_278),
.B2(n_267),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_284),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_271),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_286),
.A2(n_185),
.B1(n_229),
.B2(n_219),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_301),
.A2(n_260),
.B(n_234),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_332),
.A2(n_289),
.B(n_277),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_266),
.B(n_221),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_268),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_280),
.B(n_243),
.C(n_240),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_264),
.B(n_243),
.C(n_232),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_262),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_339),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_SL g390 ( 
.A(n_342),
.B(n_363),
.C(n_341),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_340),
.Y(n_344)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_344),
.Y(n_377)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_345),
.Y(n_381)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_312),
.A2(n_295),
.B1(n_270),
.B2(n_297),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_349),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_351),
.A2(n_357),
.B1(n_365),
.B2(n_367),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_288),
.Y(n_353)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

NAND3xp33_ASAP7_75t_L g354 ( 
.A(n_305),
.B(n_269),
.C(n_296),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_354),
.B(n_304),
.Y(n_393)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_315),
.Y(n_355)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_355),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_356),
.B(n_317),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_329),
.B1(n_324),
.B2(n_309),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_268),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_306),
.C(n_338),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_320),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_359),
.B(n_366),
.Y(n_376)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_316),
.Y(n_361)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_364),
.Y(n_398)
);

AOI21xp33_ASAP7_75t_L g363 ( 
.A1(n_314),
.A2(n_302),
.B(n_224),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_310),
.A2(n_299),
.B1(n_229),
.B2(n_290),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_322),
.A2(n_224),
.B1(n_253),
.B2(n_291),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_309),
.A2(n_275),
.B1(n_253),
.B2(n_260),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_321),
.B(n_282),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_368),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_305),
.B(n_222),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_369),
.B(n_372),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_323),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_308),
.B(n_282),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_373),
.B(n_303),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_342),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_306),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_389),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_337),
.C(n_336),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_395),
.C(n_399),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_382),
.B(n_395),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_350),
.B(n_332),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_383),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_351),
.A2(n_318),
.B1(n_336),
.B2(n_317),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_384),
.A2(n_392),
.B1(n_400),
.B2(n_311),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_359),
.A2(n_313),
.B1(n_330),
.B2(n_303),
.Y(n_387)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_387),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_352),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_390),
.A2(n_393),
.B1(n_371),
.B2(n_383),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_391),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_357),
.A2(n_326),
.B1(n_328),
.B2(n_307),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_334),
.C(n_307),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_348),
.B(n_328),
.C(n_340),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_343),
.A2(n_328),
.B1(n_304),
.B2(n_339),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_353),
.B(n_325),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_347),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_346),
.B(n_325),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_402),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_346),
.Y(n_406)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_406),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_398),
.A2(n_343),
.B1(n_350),
.B2(n_341),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_407),
.A2(n_375),
.B1(n_400),
.B2(n_401),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_373),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_412),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_417),
.C(n_421),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_368),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_410),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_370),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_376),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_414),
.Y(n_442)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_394),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_282),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_374),
.B(n_367),
.C(n_365),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_390),
.A2(n_370),
.B1(n_362),
.B2(n_366),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_9),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_378),
.B(n_389),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_420),
.B(n_422),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_379),
.B(n_364),
.C(n_355),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_382),
.B(n_361),
.C(n_360),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_377),
.C(n_397),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_384),
.B(n_372),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_424),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_422),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_388),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_427),
.B(n_9),
.Y(n_449)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_396),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_282),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_429),
.A2(n_399),
.B1(n_386),
.B2(n_375),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_411),
.A2(n_383),
.B(n_398),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_430),
.A2(n_406),
.B(n_417),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_432),
.Y(n_456)
);

AO21x1_ASAP7_75t_L g432 ( 
.A1(n_412),
.A2(n_386),
.B(n_392),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_447),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_423),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_403),
.C(n_323),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_439),
.C(n_441),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_311),
.C(n_222),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_415),
.C(n_421),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_443),
.B(n_449),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_199),
.C(n_203),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_169),
.C(n_204),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_448),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_9),
.Y(n_466)
);

AO22x1_ASAP7_75t_L g452 ( 
.A1(n_446),
.A2(n_407),
.B1(n_411),
.B2(n_410),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_453),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_405),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_425),
.Y(n_454)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_454),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_436),
.Y(n_455)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_455),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_439),
.Y(n_473)
);

NAND2x1_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_409),
.Y(n_458)
);

MAJx2_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_435),
.C(n_441),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_404),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_461),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_463),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_433),
.A2(n_414),
.B1(n_429),
.B2(n_426),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_444),
.C(n_447),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_466),
.B(n_9),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_456),
.A2(n_434),
.B1(n_450),
.B2(n_432),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_470),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_452),
.A2(n_431),
.B(n_438),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_471),
.A2(n_478),
.B(n_479),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_473),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_481),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_444),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_464),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_457),
.A2(n_451),
.B(n_462),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_458),
.A2(n_435),
.B(n_445),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_482),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g494 ( 
.A(n_481),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_169),
.Y(n_482)
);

AO21x1_ASAP7_75t_L g499 ( 
.A1(n_484),
.A2(n_486),
.B(n_492),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_473),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_478),
.A2(n_459),
.B(n_467),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_475),
.Y(n_487)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_487),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_472),
.B(n_461),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_491),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_468),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_459),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_468),
.A2(n_465),
.B(n_466),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_495),
.B(n_479),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_493),
.Y(n_496)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_496),
.Y(n_507)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_497),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_501),
.B(n_504),
.C(n_484),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_470),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_502),
.A2(n_503),
.B(n_474),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_490),
.B(n_469),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_492),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_505),
.B(n_506),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_497),
.A2(n_488),
.B(n_471),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_169),
.C(n_204),
.Y(n_512)
);

AOI331xp33_ASAP7_75t_L g511 ( 
.A1(n_509),
.A2(n_500),
.A3(n_499),
.B1(n_483),
.B2(n_498),
.B3(n_477),
.C1(n_204),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_511),
.B(n_512),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_510),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_514),
.A2(n_507),
.B(n_12),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_513),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_13),
.Y(n_517)
);


endmodule