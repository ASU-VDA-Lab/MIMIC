module fake_jpeg_8349_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_31),
.Y(n_35)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_20),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_36),
.B(n_26),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_21),
.B1(n_24),
.B2(n_15),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_15),
.B1(n_24),
.B2(n_13),
.Y(n_49)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_2),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_54),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_1),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_28),
.B1(n_17),
.B2(n_23),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_33),
.B1(n_23),
.B2(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_32),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_56),
.Y(n_73)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_40),
.B1(n_38),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_66),
.B1(n_19),
.B2(n_22),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_19),
.B1(n_22),
.B2(n_25),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_72),
.B1(n_46),
.B2(n_57),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_79),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_25),
.B1(n_32),
.B2(n_26),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_79),
.C(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_1),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_55),
.B1(n_56),
.B2(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_3),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_88),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_46),
.C(n_57),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_91),
.C(n_3),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_60),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_65),
.B1(n_45),
.B2(n_59),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

NAND2x1_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_45),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_75),
.B(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_104),
.B(n_86),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_67),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_90),
.C(n_5),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_81),
.B(n_67),
.C(n_78),
.D(n_69),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_109),
.B(n_95),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_81),
.A3(n_77),
.B1(n_69),
.B2(n_72),
.C1(n_71),
.C2(n_84),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_71),
.B(n_77),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_87),
.B(n_86),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_95),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_4),
.B(n_5),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_110),
.B(n_115),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_106),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_113),
.B1(n_99),
.B2(n_108),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_90),
.B1(n_94),
.B2(n_85),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_99),
.B1(n_105),
.B2(n_90),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_89),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_116),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_109),
.C(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_101),
.C(n_100),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_112),
.B1(n_103),
.B2(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_121),
.B(n_119),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_118),
.B1(n_5),
.B2(n_6),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_111),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_128),
.B(n_118),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_130),
.C(n_132),
.Y(n_135)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_125),
.B(n_7),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_4),
.Y(n_137)
);

OAI21x1_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_8),
.B(n_10),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_135),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_136),
.Y(n_140)
);


endmodule