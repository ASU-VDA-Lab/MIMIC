module fake_aes_41_n_19 (n_1, n_2, n_0, n_19);
input n_1;
input n_2;
input n_0;
output n_19;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_3;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_6;
wire n_4;
wire n_7;
INVxp67_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
BUFx6f_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
BUFx10_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
BUFx2_ASAP7_75t_L g7 ( .A(n_3), .Y(n_7) );
BUFx6f_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_7), .B(n_5), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_9), .B(n_7), .Y(n_12) );
OAI221xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_4), .B1(n_10), .B2(n_5), .C(n_8), .Y(n_13) );
AOI221xp5_ASAP7_75t_L g14 ( .A1(n_11), .A2(n_4), .B1(n_5), .B2(n_8), .C(n_0), .Y(n_14) );
AND2x2_ASAP7_75t_SL g15 ( .A(n_14), .B(n_11), .Y(n_15) );
OAI21xp33_ASAP7_75t_L g16 ( .A1(n_13), .A2(n_4), .B(n_1), .Y(n_16) );
AOI21xp33_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_2), .B(n_0), .Y(n_17) );
OAI22xp5_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_18) );
AOI22xp33_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_2), .B1(n_15), .B2(n_18), .Y(n_19) );
endmodule