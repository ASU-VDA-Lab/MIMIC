module fake_jpeg_5293_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_21),
.B1(n_24),
.B2(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_24),
.B1(n_21),
.B2(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_46),
.Y(n_65)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_52),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_31),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_68),
.C(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_23),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_73),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_64),
.B1(n_70),
.B2(n_13),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_37),
.B1(n_32),
.B2(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_71),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_35),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_74),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_29),
.B1(n_15),
.B2(n_13),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_16),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_23),
.B(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

XOR2x1_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_57),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_88),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_49),
.B1(n_56),
.B2(n_42),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_56),
.B1(n_42),
.B2(n_57),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_56),
.B1(n_41),
.B2(n_44),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_51),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_73),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_44),
.B1(n_41),
.B2(n_15),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_61),
.C(n_74),
.Y(n_100)
);

AO21x1_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_94),
.B(n_18),
.Y(n_112)
);

OAI22x1_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_68),
.B1(n_75),
.B2(n_41),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_75),
.B(n_63),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_98),
.B(n_101),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_100),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_82),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_72),
.C(n_61),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_89),
.C(n_72),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_68),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_82),
.B(n_79),
.C(n_81),
.D(n_74),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_109),
.Y(n_114)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_111),
.CI(n_95),
.CON(n_115),
.SN(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_78),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_76),
.B1(n_84),
.B2(n_86),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_66),
.B(n_51),
.Y(n_113)
);

OAI22x1_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_51),
.B1(n_67),
.B2(n_44),
.Y(n_119)
);

AOI321xp33_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_117),
.A3(n_121),
.B1(n_26),
.B2(n_19),
.C(n_17),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_92),
.B(n_97),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_120),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_59),
.B(n_19),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_92),
.B1(n_112),
.B2(n_103),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_109),
.C(n_106),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_115),
.C(n_59),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_26),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_59),
.Y(n_126)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_19),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_130),
.C(n_123),
.Y(n_134)
);

OAI31xp33_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_127),
.A3(n_122),
.B(n_17),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_0),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_134),
.B(n_135),
.Y(n_137)
);

AOI21x1_ASAP7_75t_L g135 ( 
.A1(n_128),
.A2(n_0),
.B(n_1),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_137),
.A2(n_5),
.B(n_6),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_138),
.B(n_7),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_7),
.Y(n_141)
);


endmodule