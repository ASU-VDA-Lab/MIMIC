module fake_jpeg_8053_n_70 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_70);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_70;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_67;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_17),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_13),
.B1(n_22),
.B2(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_47)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_50),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_24),
.B1(n_12),
.B2(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_15),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_53),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_62),
.B1(n_58),
.B2(n_44),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_46),
.C(n_42),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_57),
.B(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_67),
.B(n_56),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

XNOR2x2_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_16),
.Y(n_70)
);


endmodule