module fake_netlist_6_500_n_5374 (n_992, n_1, n_801, n_1234, n_1199, n_741, n_1027, n_625, n_1189, n_223, n_1212, n_226, n_208, n_68, n_726, n_212, n_700, n_50, n_1038, n_578, n_1003, n_365, n_168, n_1237, n_1061, n_77, n_783, n_798, n_188, n_509, n_245, n_1209, n_677, n_805, n_1151, n_396, n_350, n_78, n_442, n_480, n_142, n_1009, n_62, n_1160, n_883, n_1238, n_1032, n_1247, n_893, n_1099, n_1264, n_1192, n_471, n_424, n_369, n_287, n_415, n_830, n_65, n_230, n_461, n_873, n_141, n_383, n_1285, n_200, n_447, n_1172, n_852, n_71, n_229, n_1078, n_250, n_544, n_1140, n_35, n_1263, n_836, n_375, n_522, n_1261, n_945, n_1143, n_1232, n_616, n_658, n_1119, n_428, n_641, n_822, n_693, n_1056, n_758, n_516, n_1163, n_1180, n_943, n_491, n_42, n_772, n_666, n_371, n_940, n_770, n_567, n_405, n_213, n_538, n_1106, n_886, n_343, n_953, n_1094, n_494, n_539, n_493, n_155, n_45, n_454, n_638, n_1211, n_381, n_887, n_112, n_1280, n_713, n_126, n_58, n_976, n_224, n_48, n_734, n_1088, n_196, n_1231, n_917, n_574, n_9, n_907, n_6, n_14, n_659, n_407, n_913, n_808, n_867, n_1230, n_473, n_1193, n_1054, n_559, n_44, n_163, n_281, n_551, n_699, n_564, n_451, n_824, n_279, n_686, n_757, n_594, n_577, n_166, n_619, n_521, n_572, n_395, n_813, n_323, n_606, n_818, n_1123, n_92, n_513, n_645, n_331, n_916, n_483, n_102, n_608, n_261, n_630, n_32, n_541, n_512, n_121, n_433, n_792, n_476, n_2, n_219, n_264, n_263, n_1162, n_860, n_788, n_939, n_821, n_938, n_1068, n_329, n_982, n_549, n_1075, n_408, n_932, n_61, n_237, n_243, n_979, n_905, n_117, n_175, n_322, n_993, n_689, n_354, n_134, n_1278, n_547, n_558, n_1064, n_634, n_136, n_966, n_764, n_692, n_733, n_1233, n_487, n_241, n_30, n_1107, n_1014, n_882, n_586, n_423, n_318, n_1111, n_715, n_1251, n_1265, n_88, n_530, n_277, n_618, n_199, n_1167, n_674, n_871, n_922, n_268, n_210, n_1069, n_5, n_612, n_178, n_247, n_1165, n_355, n_702, n_347, n_1175, n_328, n_429, n_1012, n_195, n_780, n_675, n_903, n_286, n_254, n_242, n_835, n_1214, n_928, n_47, n_690, n_850, n_816, n_1157, n_1188, n_877, n_604, n_825, n_728, n_1063, n_26, n_55, n_267, n_1124, n_515, n_598, n_696, n_961, n_437, n_1082, n_593, n_514, n_687, n_697, n_890, n_637, n_295, n_701, n_950, n_388, n_190, n_484, n_170, n_891, n_949, n_678, n_283, n_91, n_507, n_968, n_909, n_881, n_1008, n_760, n_590, n_63, n_362, n_148, n_161, n_22, n_462, n_1033, n_1052, n_304, n_694, n_125, n_297, n_595, n_627, n_524, n_342, n_1044, n_449, n_131, n_1208, n_1164, n_1072, n_495, n_815, n_1100, n_585, n_840, n_874, n_1128, n_382, n_673, n_1071, n_1067, n_898, n_255, n_284, n_865, n_925, n_1101, n_15, n_1026, n_38, n_289, n_615, n_1249, n_59, n_1127, n_320, n_108, n_639, n_963, n_794, n_727, n_894, n_685, n_353, n_605, n_826, n_872, n_1139, n_86, n_104, n_718, n_1018, n_542, n_847, n_644, n_682, n_851, n_305, n_72, n_996, n_532, n_173, n_413, n_791, n_510, n_837, n_79, n_948, n_704, n_977, n_1005, n_536, n_622, n_147, n_581, n_765, n_432, n_987, n_631, n_720, n_153, n_842, n_156, n_145, n_843, n_656, n_989, n_1277, n_797, n_1246, n_899, n_189, n_738, n_1035, n_294, n_499, n_705, n_11, n_1004, n_1176, n_1022, n_614, n_529, n_425, n_684, n_1181, n_37, n_486, n_947, n_1117, n_1087, n_648, n_657, n_1049, n_803, n_290, n_118, n_926, n_927, n_919, n_478, n_929, n_107, n_1228, n_417, n_446, n_89, n_777, n_272, n_526, n_1183, n_69, n_293, n_53, n_458, n_1070, n_998, n_16, n_717, n_18, n_154, n_1178, n_98, n_1073, n_1000, n_796, n_252, n_1195, n_184, n_552, n_216, n_912, n_745, n_1284, n_1142, n_716, n_623, n_1048, n_1201, n_884, n_731, n_755, n_931, n_1021, n_474, n_527, n_683, n_811, n_1207, n_312, n_66, n_958, n_292, n_1250, n_100, n_1137, n_880, n_889, n_150, n_589, n_819, n_767, n_600, n_964, n_831, n_477, n_954, n_864, n_1110, n_399, n_124, n_211, n_231, n_40, n_505, n_319, n_537, n_311, n_10, n_403, n_1080, n_723, n_596, n_123, n_546, n_562, n_1141, n_1268, n_386, n_1220, n_556, n_162, n_1136, n_128, n_1125, n_970, n_642, n_995, n_276, n_1159, n_1092, n_441, n_221, n_1060, n_444, n_146, n_1252, n_1223, n_303, n_511, n_193, n_1286, n_1053, n_416, n_520, n_418, n_1093, n_113, n_4, n_266, n_296, n_775, n_651, n_1153, n_439, n_217, n_518, n_1185, n_453, n_215, n_914, n_759, n_426, n_317, n_90, n_54, n_488, n_497, n_773, n_920, n_99, n_13, n_1224, n_1135, n_1169, n_1179, n_401, n_324, n_335, n_463, n_1243, n_848, n_120, n_301, n_274, n_1096, n_1091, n_36, n_1267, n_1281, n_983, n_427, n_496, n_906, n_688, n_1077, n_351, n_259, n_177, n_385, n_858, n_613, n_736, n_501, n_956, n_960, n_663, n_856, n_379, n_778, n_1134, n_410, n_1129, n_554, n_602, n_664, n_171, n_169, n_435, n_793, n_326, n_587, n_580, n_762, n_1030, n_1202, n_465, n_1079, n_341, n_828, n_607, n_316, n_419, n_28, n_1103, n_144, n_1203, n_820, n_951, n_106, n_725, n_952, n_999, n_358, n_1254, n_160, n_186, n_0, n_368, n_575, n_994, n_732, n_974, n_392, n_724, n_1020, n_1042, n_628, n_1273, n_557, n_349, n_617, n_845, n_807, n_1036, n_140, n_1138, n_1275, n_485, n_67, n_443, n_892, n_768, n_421, n_238, n_1095, n_202, n_597, n_280, n_1270, n_1187, n_610, n_1024, n_198, n_179, n_248, n_517, n_667, n_1206, n_621, n_1037, n_1279, n_1115, n_750, n_901, n_468, n_923, n_504, n_183, n_1015, n_466, n_1057, n_603, n_991, n_235, n_1126, n_340, n_710, n_1108, n_1182, n_39, n_73, n_785, n_746, n_609, n_101, n_167, n_127, n_1168, n_1216, n_133, n_96, n_1287, n_302, n_380, n_137, n_20, n_1190, n_397, n_122, n_34, n_1262, n_218, n_1213, n_70, n_172, n_1272, n_239, n_97, n_782, n_490, n_220, n_809, n_1043, n_986, n_80, n_1081, n_402, n_352, n_800, n_1084, n_1171, n_460, n_662, n_374, n_1152, n_450, n_921, n_711, n_579, n_937, n_370, n_650, n_1046, n_1145, n_330, n_1121, n_1102, n_972, n_258, n_456, n_260, n_313, n_624, n_962, n_1041, n_565, n_356, n_936, n_1288, n_1186, n_1062, n_885, n_896, n_83, n_654, n_411, n_152, n_1222, n_599, n_776, n_321, n_105, n_227, n_204, n_482, n_934, n_420, n_394, n_164, n_23, n_942, n_543, n_1271, n_1225, n_325, n_804, n_464, n_533, n_806, n_879, n_959, n_584, n_244, n_76, n_548, n_94, n_282, n_833, n_523, n_707, n_345, n_799, n_1155, n_139, n_41, n_273, n_787, n_1146, n_159, n_1086, n_1066, n_157, n_1282, n_550, n_275, n_652, n_560, n_1241, n_569, n_737, n_1235, n_1229, n_306, n_21, n_346, n_3, n_1029, n_790, n_138, n_1210, n_49, n_299, n_1248, n_902, n_333, n_1047, n_431, n_24, n_459, n_1269, n_502, n_672, n_1257, n_285, n_85, n_655, n_706, n_1045, n_786, n_1236, n_834, n_19, n_29, n_75, n_743, n_766, n_430, n_1002, n_545, n_489, n_251, n_1019, n_636, n_729, n_110, n_151, n_876, n_774, n_660, n_438, n_1200, n_479, n_869, n_1154, n_1113, n_646, n_528, n_391, n_1098, n_817, n_262, n_187, n_897, n_846, n_841, n_1001, n_508, n_1050, n_1177, n_332, n_1150, n_398, n_1191, n_566, n_1023, n_1076, n_1118, n_194, n_57, n_1007, n_855, n_52, n_591, n_256, n_853, n_440, n_695, n_875, n_209, n_367, n_680, n_661, n_278, n_1256, n_671, n_7, n_933, n_740, n_703, n_978, n_384, n_1217, n_751, n_749, n_310, n_969, n_988, n_1065, n_84, n_1255, n_568, n_143, n_180, n_1204, n_823, n_1132, n_643, n_233, n_698, n_1074, n_739, n_400, n_955, n_337, n_214, n_246, n_1097, n_935, n_781, n_789, n_1130, n_181, n_182, n_573, n_769, n_676, n_327, n_1120, n_832, n_555, n_389, n_814, n_669, n_176, n_114, n_300, n_222, n_747, n_74, n_1105, n_721, n_742, n_535, n_691, n_372, n_111, n_314, n_378, n_1196, n_377, n_863, n_601, n_338, n_1283, n_918, n_748, n_506, n_1114, n_56, n_763, n_1147, n_360, n_119, n_957, n_895, n_866, n_1227, n_191, n_387, n_452, n_744, n_971, n_946, n_344, n_761, n_1205, n_1258, n_174, n_1173, n_525, n_1116, n_611, n_1219, n_8, n_1174, n_1016, n_795, n_1221, n_1245, n_838, n_129, n_647, n_197, n_844, n_17, n_448, n_1017, n_1083, n_109, n_445, n_930, n_888, n_1112, n_234, n_910, n_911, n_82, n_27, n_236, n_653, n_752, n_908, n_944, n_576, n_1028, n_472, n_270, n_414, n_563, n_1011, n_1215, n_25, n_93, n_839, n_708, n_668, n_626, n_990, n_779, n_1104, n_854, n_1058, n_498, n_1122, n_870, n_904, n_1253, n_709, n_1266, n_366, n_103, n_1109, n_185, n_712, n_348, n_1276, n_376, n_390, n_1148, n_31, n_334, n_1161, n_1085, n_232, n_46, n_1239, n_771, n_470, n_475, n_924, n_298, n_492, n_1149, n_265, n_1184, n_228, n_719, n_455, n_363, n_1090, n_592, n_829, n_1156, n_393, n_984, n_503, n_132, n_868, n_570, n_859, n_406, n_735, n_878, n_620, n_130, n_519, n_307, n_469, n_1218, n_500, n_981, n_714, n_291, n_1144, n_357, n_985, n_481, n_997, n_802, n_561, n_33, n_980, n_1198, n_436, n_116, n_409, n_1244, n_240, n_756, n_810, n_1133, n_635, n_95, n_1194, n_1051, n_253, n_583, n_249, n_201, n_1039, n_1034, n_1158, n_754, n_941, n_975, n_1031, n_115, n_553, n_43, n_849, n_753, n_467, n_269, n_359, n_973, n_1055, n_582, n_861, n_857, n_967, n_571, n_271, n_404, n_158, n_206, n_679, n_633, n_1170, n_665, n_588, n_225, n_1260, n_308, n_309, n_1010, n_149, n_1040, n_915, n_632, n_1166, n_812, n_1131, n_534, n_1006, n_373, n_87, n_257, n_730, n_670, n_203, n_207, n_1089, n_205, n_1242, n_681, n_1226, n_1274, n_412, n_640, n_81, n_965, n_339, n_784, n_315, n_434, n_64, n_288, n_1059, n_1197, n_422, n_722, n_862, n_135, n_165, n_540, n_457, n_364, n_629, n_900, n_531, n_827, n_60, n_361, n_1025, n_336, n_12, n_1013, n_1259, n_192, n_51, n_649, n_1240, n_5374);

input n_992;
input n_1;
input n_801;
input n_1234;
input n_1199;
input n_741;
input n_1027;
input n_625;
input n_1189;
input n_223;
input n_1212;
input n_226;
input n_208;
input n_68;
input n_726;
input n_212;
input n_700;
input n_50;
input n_1038;
input n_578;
input n_1003;
input n_365;
input n_168;
input n_1237;
input n_1061;
input n_77;
input n_783;
input n_798;
input n_188;
input n_509;
input n_245;
input n_1209;
input n_677;
input n_805;
input n_1151;
input n_396;
input n_350;
input n_78;
input n_442;
input n_480;
input n_142;
input n_1009;
input n_62;
input n_1160;
input n_883;
input n_1238;
input n_1032;
input n_1247;
input n_893;
input n_1099;
input n_1264;
input n_1192;
input n_471;
input n_424;
input n_369;
input n_287;
input n_415;
input n_830;
input n_65;
input n_230;
input n_461;
input n_873;
input n_141;
input n_383;
input n_1285;
input n_200;
input n_447;
input n_1172;
input n_852;
input n_71;
input n_229;
input n_1078;
input n_250;
input n_544;
input n_1140;
input n_35;
input n_1263;
input n_836;
input n_375;
input n_522;
input n_1261;
input n_945;
input n_1143;
input n_1232;
input n_616;
input n_658;
input n_1119;
input n_428;
input n_641;
input n_822;
input n_693;
input n_1056;
input n_758;
input n_516;
input n_1163;
input n_1180;
input n_943;
input n_491;
input n_42;
input n_772;
input n_666;
input n_371;
input n_940;
input n_770;
input n_567;
input n_405;
input n_213;
input n_538;
input n_1106;
input n_886;
input n_343;
input n_953;
input n_1094;
input n_494;
input n_539;
input n_493;
input n_155;
input n_45;
input n_454;
input n_638;
input n_1211;
input n_381;
input n_887;
input n_112;
input n_1280;
input n_713;
input n_126;
input n_58;
input n_976;
input n_224;
input n_48;
input n_734;
input n_1088;
input n_196;
input n_1231;
input n_917;
input n_574;
input n_9;
input n_907;
input n_6;
input n_14;
input n_659;
input n_407;
input n_913;
input n_808;
input n_867;
input n_1230;
input n_473;
input n_1193;
input n_1054;
input n_559;
input n_44;
input n_163;
input n_281;
input n_551;
input n_699;
input n_564;
input n_451;
input n_824;
input n_279;
input n_686;
input n_757;
input n_594;
input n_577;
input n_166;
input n_619;
input n_521;
input n_572;
input n_395;
input n_813;
input n_323;
input n_606;
input n_818;
input n_1123;
input n_92;
input n_513;
input n_645;
input n_331;
input n_916;
input n_483;
input n_102;
input n_608;
input n_261;
input n_630;
input n_32;
input n_541;
input n_512;
input n_121;
input n_433;
input n_792;
input n_476;
input n_2;
input n_219;
input n_264;
input n_263;
input n_1162;
input n_860;
input n_788;
input n_939;
input n_821;
input n_938;
input n_1068;
input n_329;
input n_982;
input n_549;
input n_1075;
input n_408;
input n_932;
input n_61;
input n_237;
input n_243;
input n_979;
input n_905;
input n_117;
input n_175;
input n_322;
input n_993;
input n_689;
input n_354;
input n_134;
input n_1278;
input n_547;
input n_558;
input n_1064;
input n_634;
input n_136;
input n_966;
input n_764;
input n_692;
input n_733;
input n_1233;
input n_487;
input n_241;
input n_30;
input n_1107;
input n_1014;
input n_882;
input n_586;
input n_423;
input n_318;
input n_1111;
input n_715;
input n_1251;
input n_1265;
input n_88;
input n_530;
input n_277;
input n_618;
input n_199;
input n_1167;
input n_674;
input n_871;
input n_922;
input n_268;
input n_210;
input n_1069;
input n_5;
input n_612;
input n_178;
input n_247;
input n_1165;
input n_355;
input n_702;
input n_347;
input n_1175;
input n_328;
input n_429;
input n_1012;
input n_195;
input n_780;
input n_675;
input n_903;
input n_286;
input n_254;
input n_242;
input n_835;
input n_1214;
input n_928;
input n_47;
input n_690;
input n_850;
input n_816;
input n_1157;
input n_1188;
input n_877;
input n_604;
input n_825;
input n_728;
input n_1063;
input n_26;
input n_55;
input n_267;
input n_1124;
input n_515;
input n_598;
input n_696;
input n_961;
input n_437;
input n_1082;
input n_593;
input n_514;
input n_687;
input n_697;
input n_890;
input n_637;
input n_295;
input n_701;
input n_950;
input n_388;
input n_190;
input n_484;
input n_170;
input n_891;
input n_949;
input n_678;
input n_283;
input n_91;
input n_507;
input n_968;
input n_909;
input n_881;
input n_1008;
input n_760;
input n_590;
input n_63;
input n_362;
input n_148;
input n_161;
input n_22;
input n_462;
input n_1033;
input n_1052;
input n_304;
input n_694;
input n_125;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_1044;
input n_449;
input n_131;
input n_1208;
input n_1164;
input n_1072;
input n_495;
input n_815;
input n_1100;
input n_585;
input n_840;
input n_874;
input n_1128;
input n_382;
input n_673;
input n_1071;
input n_1067;
input n_898;
input n_255;
input n_284;
input n_865;
input n_925;
input n_1101;
input n_15;
input n_1026;
input n_38;
input n_289;
input n_615;
input n_1249;
input n_59;
input n_1127;
input n_320;
input n_108;
input n_639;
input n_963;
input n_794;
input n_727;
input n_894;
input n_685;
input n_353;
input n_605;
input n_826;
input n_872;
input n_1139;
input n_86;
input n_104;
input n_718;
input n_1018;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_305;
input n_72;
input n_996;
input n_532;
input n_173;
input n_413;
input n_791;
input n_510;
input n_837;
input n_79;
input n_948;
input n_704;
input n_977;
input n_1005;
input n_536;
input n_622;
input n_147;
input n_581;
input n_765;
input n_432;
input n_987;
input n_631;
input n_720;
input n_153;
input n_842;
input n_156;
input n_145;
input n_843;
input n_656;
input n_989;
input n_1277;
input n_797;
input n_1246;
input n_899;
input n_189;
input n_738;
input n_1035;
input n_294;
input n_499;
input n_705;
input n_11;
input n_1004;
input n_1176;
input n_1022;
input n_614;
input n_529;
input n_425;
input n_684;
input n_1181;
input n_37;
input n_486;
input n_947;
input n_1117;
input n_1087;
input n_648;
input n_657;
input n_1049;
input n_803;
input n_290;
input n_118;
input n_926;
input n_927;
input n_919;
input n_478;
input n_929;
input n_107;
input n_1228;
input n_417;
input n_446;
input n_89;
input n_777;
input n_272;
input n_526;
input n_1183;
input n_69;
input n_293;
input n_53;
input n_458;
input n_1070;
input n_998;
input n_16;
input n_717;
input n_18;
input n_154;
input n_1178;
input n_98;
input n_1073;
input n_1000;
input n_796;
input n_252;
input n_1195;
input n_184;
input n_552;
input n_216;
input n_912;
input n_745;
input n_1284;
input n_1142;
input n_716;
input n_623;
input n_1048;
input n_1201;
input n_884;
input n_731;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_683;
input n_811;
input n_1207;
input n_312;
input n_66;
input n_958;
input n_292;
input n_1250;
input n_100;
input n_1137;
input n_880;
input n_889;
input n_150;
input n_589;
input n_819;
input n_767;
input n_600;
input n_964;
input n_831;
input n_477;
input n_954;
input n_864;
input n_1110;
input n_399;
input n_124;
input n_211;
input n_231;
input n_40;
input n_505;
input n_319;
input n_537;
input n_311;
input n_10;
input n_403;
input n_1080;
input n_723;
input n_596;
input n_123;
input n_546;
input n_562;
input n_1141;
input n_1268;
input n_386;
input n_1220;
input n_556;
input n_162;
input n_1136;
input n_128;
input n_1125;
input n_970;
input n_642;
input n_995;
input n_276;
input n_1159;
input n_1092;
input n_441;
input n_221;
input n_1060;
input n_444;
input n_146;
input n_1252;
input n_1223;
input n_303;
input n_511;
input n_193;
input n_1286;
input n_1053;
input n_416;
input n_520;
input n_418;
input n_1093;
input n_113;
input n_4;
input n_266;
input n_296;
input n_775;
input n_651;
input n_1153;
input n_439;
input n_217;
input n_518;
input n_1185;
input n_453;
input n_215;
input n_914;
input n_759;
input n_426;
input n_317;
input n_90;
input n_54;
input n_488;
input n_497;
input n_773;
input n_920;
input n_99;
input n_13;
input n_1224;
input n_1135;
input n_1169;
input n_1179;
input n_401;
input n_324;
input n_335;
input n_463;
input n_1243;
input n_848;
input n_120;
input n_301;
input n_274;
input n_1096;
input n_1091;
input n_36;
input n_1267;
input n_1281;
input n_983;
input n_427;
input n_496;
input n_906;
input n_688;
input n_1077;
input n_351;
input n_259;
input n_177;
input n_385;
input n_858;
input n_613;
input n_736;
input n_501;
input n_956;
input n_960;
input n_663;
input n_856;
input n_379;
input n_778;
input n_1134;
input n_410;
input n_1129;
input n_554;
input n_602;
input n_664;
input n_171;
input n_169;
input n_435;
input n_793;
input n_326;
input n_587;
input n_580;
input n_762;
input n_1030;
input n_1202;
input n_465;
input n_1079;
input n_341;
input n_828;
input n_607;
input n_316;
input n_419;
input n_28;
input n_1103;
input n_144;
input n_1203;
input n_820;
input n_951;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_1254;
input n_160;
input n_186;
input n_0;
input n_368;
input n_575;
input n_994;
input n_732;
input n_974;
input n_392;
input n_724;
input n_1020;
input n_1042;
input n_628;
input n_1273;
input n_557;
input n_349;
input n_617;
input n_845;
input n_807;
input n_1036;
input n_140;
input n_1138;
input n_1275;
input n_485;
input n_67;
input n_443;
input n_892;
input n_768;
input n_421;
input n_238;
input n_1095;
input n_202;
input n_597;
input n_280;
input n_1270;
input n_1187;
input n_610;
input n_1024;
input n_198;
input n_179;
input n_248;
input n_517;
input n_667;
input n_1206;
input n_621;
input n_1037;
input n_1279;
input n_1115;
input n_750;
input n_901;
input n_468;
input n_923;
input n_504;
input n_183;
input n_1015;
input n_466;
input n_1057;
input n_603;
input n_991;
input n_235;
input n_1126;
input n_340;
input n_710;
input n_1108;
input n_1182;
input n_39;
input n_73;
input n_785;
input n_746;
input n_609;
input n_101;
input n_167;
input n_127;
input n_1168;
input n_1216;
input n_133;
input n_96;
input n_1287;
input n_302;
input n_380;
input n_137;
input n_20;
input n_1190;
input n_397;
input n_122;
input n_34;
input n_1262;
input n_218;
input n_1213;
input n_70;
input n_172;
input n_1272;
input n_239;
input n_97;
input n_782;
input n_490;
input n_220;
input n_809;
input n_1043;
input n_986;
input n_80;
input n_1081;
input n_402;
input n_352;
input n_800;
input n_1084;
input n_1171;
input n_460;
input n_662;
input n_374;
input n_1152;
input n_450;
input n_921;
input n_711;
input n_579;
input n_937;
input n_370;
input n_650;
input n_1046;
input n_1145;
input n_330;
input n_1121;
input n_1102;
input n_972;
input n_258;
input n_456;
input n_260;
input n_313;
input n_624;
input n_962;
input n_1041;
input n_565;
input n_356;
input n_936;
input n_1288;
input n_1186;
input n_1062;
input n_885;
input n_896;
input n_83;
input n_654;
input n_411;
input n_152;
input n_1222;
input n_599;
input n_776;
input n_321;
input n_105;
input n_227;
input n_204;
input n_482;
input n_934;
input n_420;
input n_394;
input n_164;
input n_23;
input n_942;
input n_543;
input n_1271;
input n_1225;
input n_325;
input n_804;
input n_464;
input n_533;
input n_806;
input n_879;
input n_959;
input n_584;
input n_244;
input n_76;
input n_548;
input n_94;
input n_282;
input n_833;
input n_523;
input n_707;
input n_345;
input n_799;
input n_1155;
input n_139;
input n_41;
input n_273;
input n_787;
input n_1146;
input n_159;
input n_1086;
input n_1066;
input n_157;
input n_1282;
input n_550;
input n_275;
input n_652;
input n_560;
input n_1241;
input n_569;
input n_737;
input n_1235;
input n_1229;
input n_306;
input n_21;
input n_346;
input n_3;
input n_1029;
input n_790;
input n_138;
input n_1210;
input n_49;
input n_299;
input n_1248;
input n_902;
input n_333;
input n_1047;
input n_431;
input n_24;
input n_459;
input n_1269;
input n_502;
input n_672;
input n_1257;
input n_285;
input n_85;
input n_655;
input n_706;
input n_1045;
input n_786;
input n_1236;
input n_834;
input n_19;
input n_29;
input n_75;
input n_743;
input n_766;
input n_430;
input n_1002;
input n_545;
input n_489;
input n_251;
input n_1019;
input n_636;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_660;
input n_438;
input n_1200;
input n_479;
input n_869;
input n_1154;
input n_1113;
input n_646;
input n_528;
input n_391;
input n_1098;
input n_817;
input n_262;
input n_187;
input n_897;
input n_846;
input n_841;
input n_1001;
input n_508;
input n_1050;
input n_1177;
input n_332;
input n_1150;
input n_398;
input n_1191;
input n_566;
input n_1023;
input n_1076;
input n_1118;
input n_194;
input n_57;
input n_1007;
input n_855;
input n_52;
input n_591;
input n_256;
input n_853;
input n_440;
input n_695;
input n_875;
input n_209;
input n_367;
input n_680;
input n_661;
input n_278;
input n_1256;
input n_671;
input n_7;
input n_933;
input n_740;
input n_703;
input n_978;
input n_384;
input n_1217;
input n_751;
input n_749;
input n_310;
input n_969;
input n_988;
input n_1065;
input n_84;
input n_1255;
input n_568;
input n_143;
input n_180;
input n_1204;
input n_823;
input n_1132;
input n_643;
input n_233;
input n_698;
input n_1074;
input n_739;
input n_400;
input n_955;
input n_337;
input n_214;
input n_246;
input n_1097;
input n_935;
input n_781;
input n_789;
input n_1130;
input n_181;
input n_182;
input n_573;
input n_769;
input n_676;
input n_327;
input n_1120;
input n_832;
input n_555;
input n_389;
input n_814;
input n_669;
input n_176;
input n_114;
input n_300;
input n_222;
input n_747;
input n_74;
input n_1105;
input n_721;
input n_742;
input n_535;
input n_691;
input n_372;
input n_111;
input n_314;
input n_378;
input n_1196;
input n_377;
input n_863;
input n_601;
input n_338;
input n_1283;
input n_918;
input n_748;
input n_506;
input n_1114;
input n_56;
input n_763;
input n_1147;
input n_360;
input n_119;
input n_957;
input n_895;
input n_866;
input n_1227;
input n_191;
input n_387;
input n_452;
input n_744;
input n_971;
input n_946;
input n_344;
input n_761;
input n_1205;
input n_1258;
input n_174;
input n_1173;
input n_525;
input n_1116;
input n_611;
input n_1219;
input n_8;
input n_1174;
input n_1016;
input n_795;
input n_1221;
input n_1245;
input n_838;
input n_129;
input n_647;
input n_197;
input n_844;
input n_17;
input n_448;
input n_1017;
input n_1083;
input n_109;
input n_445;
input n_930;
input n_888;
input n_1112;
input n_234;
input n_910;
input n_911;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_908;
input n_944;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_414;
input n_563;
input n_1011;
input n_1215;
input n_25;
input n_93;
input n_839;
input n_708;
input n_668;
input n_626;
input n_990;
input n_779;
input n_1104;
input n_854;
input n_1058;
input n_498;
input n_1122;
input n_870;
input n_904;
input n_1253;
input n_709;
input n_1266;
input n_366;
input n_103;
input n_1109;
input n_185;
input n_712;
input n_348;
input n_1276;
input n_376;
input n_390;
input n_1148;
input n_31;
input n_334;
input n_1161;
input n_1085;
input n_232;
input n_46;
input n_1239;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_492;
input n_1149;
input n_265;
input n_1184;
input n_228;
input n_719;
input n_455;
input n_363;
input n_1090;
input n_592;
input n_829;
input n_1156;
input n_393;
input n_984;
input n_503;
input n_132;
input n_868;
input n_570;
input n_859;
input n_406;
input n_735;
input n_878;
input n_620;
input n_130;
input n_519;
input n_307;
input n_469;
input n_1218;
input n_500;
input n_981;
input n_714;
input n_291;
input n_1144;
input n_357;
input n_985;
input n_481;
input n_997;
input n_802;
input n_561;
input n_33;
input n_980;
input n_1198;
input n_436;
input n_116;
input n_409;
input n_1244;
input n_240;
input n_756;
input n_810;
input n_1133;
input n_635;
input n_95;
input n_1194;
input n_1051;
input n_253;
input n_583;
input n_249;
input n_201;
input n_1039;
input n_1034;
input n_1158;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_553;
input n_43;
input n_849;
input n_753;
input n_467;
input n_269;
input n_359;
input n_973;
input n_1055;
input n_582;
input n_861;
input n_857;
input n_967;
input n_571;
input n_271;
input n_404;
input n_158;
input n_206;
input n_679;
input n_633;
input n_1170;
input n_665;
input n_588;
input n_225;
input n_1260;
input n_308;
input n_309;
input n_1010;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_1166;
input n_812;
input n_1131;
input n_534;
input n_1006;
input n_373;
input n_87;
input n_257;
input n_730;
input n_670;
input n_203;
input n_207;
input n_1089;
input n_205;
input n_1242;
input n_681;
input n_1226;
input n_1274;
input n_412;
input n_640;
input n_81;
input n_965;
input n_339;
input n_784;
input n_315;
input n_434;
input n_64;
input n_288;
input n_1059;
input n_1197;
input n_422;
input n_722;
input n_862;
input n_135;
input n_165;
input n_540;
input n_457;
input n_364;
input n_629;
input n_900;
input n_531;
input n_827;
input n_60;
input n_361;
input n_1025;
input n_336;
input n_12;
input n_1013;
input n_1259;
input n_192;
input n_51;
input n_649;
input n_1240;

output n_5374;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_1351;
wire n_5254;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_3089;
wire n_4978;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_4686;
wire n_2317;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_5279;
wire n_2786;
wire n_5239;
wire n_1971;
wire n_1781;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_4814;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_2625;
wire n_1400;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_2764;
wire n_2895;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5226;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_4697;
wire n_4289;
wire n_4288;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_5183;
wire n_2145;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_1932;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1512;
wire n_1451;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_3179;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_4345;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_4528;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_1529;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_5035;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1398;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_5359;
wire n_1955;
wire n_1791;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_3299;
wire n_1419;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_5180;
wire n_2049;
wire n_5182;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_4761;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_4189;
wire n_3817;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_1642;
wire n_3210;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_3292;
wire n_1496;
wire n_2007;
wire n_2039;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_4512;
wire n_1378;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_5124;
wire n_3951;
wire n_3569;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_1338;
wire n_3027;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1461;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_4027;
wire n_3154;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1570;
wire n_1702;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_3552;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_5335;
wire n_3444;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_1890;
wire n_3017;
wire n_2477;
wire n_1805;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_5274;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_3266;
wire n_3574;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_4504;
wire n_3844;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_5248;
wire n_1708;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_2356;
wire n_1511;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_2739;
wire n_1620;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_4047;
wire n_3413;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_4320;
wire n_3884;
wire n_5139;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_3798;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_4277;
wire n_4526;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_3725;
wire n_3933;
wire n_2311;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_1987;
wire n_2271;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_2954;
wire n_2728;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_3405;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_3442;
wire n_1880;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_4991;
wire n_2554;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_5087;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_3133;
wire n_1959;
wire n_5257;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_2604;
wire n_2407;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_3654;
wire n_2848;
wire n_1849;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5015;
wire n_4339;
wire n_2338;
wire n_3324;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_5282;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1951;
wire n_4362;
wire n_3311;
wire n_3913;
wire n_5121;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_4404;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_3869;
wire n_1901;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_2315;
wire n_4132;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_3234;
wire n_2276;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_3250;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_2598;
wire n_1683;
wire n_1916;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_4016;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2808;
wire n_2037;
wire n_4567;
wire n_5150;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_5348;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_3045;
wire n_3821;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_2390;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_4170;
wire n_4143;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_3515;
wire n_2951;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_4543;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_4910;
wire n_3083;
wire n_3049;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5203;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_4521;
wire n_1566;
wire n_3204;
wire n_4920;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_5266;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_4730;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_2256;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_2806;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_2378;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_2593;
wire n_4255;
wire n_4071;
wire n_3568;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_4297;
wire n_2907;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_1309;
wire n_2961;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_1530;
wire n_4745;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_3599;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_4800;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_3785;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_3519;
wire n_2082;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_3805;
wire n_1990;
wire n_2943;
wire n_5205;
wire n_3252;
wire n_1634;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_5372;
wire n_2691;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_3053;
wire n_1808;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_1809;
wire n_4280;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_4097;
wire n_1666;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_3505;
wire n_3540;
wire n_3577;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_5271;
wire n_2323;
wire n_2784;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_3407;
wire n_5313;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_2289;
wire n_1390;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_5278;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_3016;
wire n_2993;
wire n_4754;
wire n_4647;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_4983;
wire n_1778;
wire n_5287;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_3636;
wire n_2327;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_2755;
wire n_3141;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_5153;
wire n_4611;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1692;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_2699;
wire n_1828;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_2376;
wire n_1405;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_2458;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_2141;
wire n_5316;
wire n_3930;
wire n_4943;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_2021;
wire n_4942;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_3157;
wire n_4841;
wire n_3221;
wire n_1758;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_1498;
wire n_2417;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_2045;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_1994;
wire n_2566;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_4106;
wire n_3604;
wire n_1501;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_1721;
wire n_3494;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_4913;
wire n_2312;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_2042;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_4845;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_1770;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_4089;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_4865;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_5368;
wire n_4263;
wire n_1819;
wire n_3555;
wire n_3155;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_2405;
wire n_4050;
wire n_2647;
wire n_2336;
wire n_2521;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1985;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_3626;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_5022;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_3822;
wire n_4163;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_4372;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_5108;
wire n_4032;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_3921;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_4673;
wire n_2519;
wire n_3415;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_4019;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_1475;
wire n_1774;
wire n_3103;
wire n_2354;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_3144;
wire n_3244;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2357;
wire n_2025;
wire n_4654;
wire n_3640;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_2278;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_3595;
wire n_1661;
wire n_5360;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_2560;
wire n_2704;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_2901;
wire n_2611;
wire n_4358;
wire n_2653;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_1794;
wire n_4493;
wire n_4924;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_2066;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5236;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1327;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_2380;
wire n_4786;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_3493;
wire n_3774;
wire n_2910;
wire n_3268;
wire n_1785;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_2287;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_3334;
wire n_5097;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_2600;
wire n_3508;
wire n_4353;
wire n_4787;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_2440;
wire n_3521;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_2909;
wire n_5369;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_4210;
wire n_4981;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_2280;
wire n_1557;
wire n_3945;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_5065;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_966),
.Y(n_1289)
);

CKINVDCx14_ASAP7_75t_R g1290 ( 
.A(n_119),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_829),
.Y(n_1291)
);

BUFx10_ASAP7_75t_L g1292 ( 
.A(n_987),
.Y(n_1292)
);

BUFx5_ASAP7_75t_L g1293 ( 
.A(n_1172),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1034),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_588),
.Y(n_1295)
);

BUFx5_ASAP7_75t_L g1296 ( 
.A(n_258),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1125),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1234),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_202),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_730),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1283),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_452),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_945),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_391),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_620),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1009),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1161),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1018),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_289),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_715),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_176),
.Y(n_1311)
);

BUFx10_ASAP7_75t_L g1312 ( 
.A(n_974),
.Y(n_1312)
);

INVx4_ASAP7_75t_R g1313 ( 
.A(n_1150),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_609),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1028),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1255),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_708),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1210),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1211),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1199),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1223),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_675),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_877),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_548),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_993),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_614),
.Y(n_1326)
);

INVxp67_ASAP7_75t_L g1327 ( 
.A(n_740),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1214),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_256),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1195),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1209),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1239),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_307),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1259),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_87),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_999),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_948),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_407),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_453),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_337),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_452),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_839),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_838),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_881),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_574),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_957),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_78),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1019),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1080),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_480),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1136),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1025),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1037),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1267),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_920),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_320),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_206),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_855),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_227),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1055),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1031),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1038),
.Y(n_1362)
);

BUFx10_ASAP7_75t_L g1363 ( 
.A(n_142),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1010),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1184),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_582),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1227),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1279),
.Y(n_1368)
);

BUFx8_ASAP7_75t_SL g1369 ( 
.A(n_978),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_880),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1014),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_205),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1171),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_347),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_31),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_550),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_811),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1266),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_652),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_189),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1158),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_101),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_489),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_534),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1166),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_71),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_953),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_700),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_223),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_647),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_21),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1257),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_708),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1107),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_342),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_596),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_487),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1026),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1144),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_373),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_538),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_484),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1242),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1212),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_779),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_737),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1047),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1188),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1032),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_183),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_996),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1201),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_815),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_568),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_775),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_664),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_440),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_720),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_790),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1272),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_36),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1024),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1217),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_46),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_793),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_781),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1197),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_321),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1046),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_551),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_960),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_221),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_591),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_702),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1216),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_760),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_680),
.Y(n_1437)
);

BUFx10_ASAP7_75t_L g1438 ( 
.A(n_73),
.Y(n_1438)
);

BUFx10_ASAP7_75t_L g1439 ( 
.A(n_784),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1002),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_440),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_643),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_33),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1202),
.Y(n_1444)
);

CKINVDCx16_ASAP7_75t_R g1445 ( 
.A(n_1260),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_234),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1208),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_289),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_62),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_58),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1205),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_441),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_443),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_67),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_184),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_850),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_148),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_339),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1282),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_344),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1162),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1149),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_99),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_682),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1157),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_292),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_532),
.Y(n_1467)
);

INVxp67_ASAP7_75t_L g1468 ( 
.A(n_946),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_82),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1001),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_899),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_995),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_328),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1010),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_243),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1132),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_1192),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1253),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_308),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_186),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_926),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_788),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1041),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1281),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_899),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_294),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_572),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_943),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_317),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1035),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_282),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_62),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_95),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_395),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_879),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_661),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_15),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1176),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1167),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_982),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_490),
.Y(n_1501)
);

CKINVDCx16_ASAP7_75t_R g1502 ( 
.A(n_1179),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1215),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_484),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1018),
.Y(n_1505)
);

BUFx10_ASAP7_75t_L g1506 ( 
.A(n_485),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_685),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1155),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1043),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_990),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_700),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_985),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1269),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_659),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_509),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_335),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_946),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_941),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_574),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_344),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_833),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1222),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_23),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_222),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1088),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_140),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1140),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_989),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_349),
.Y(n_1529)
);

CKINVDCx16_ASAP7_75t_R g1530 ( 
.A(n_1173),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1207),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_926),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_203),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_516),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_406),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1262),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1037),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_891),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_827),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_52),
.Y(n_1540)
);

BUFx10_ASAP7_75t_L g1541 ( 
.A(n_1247),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_988),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_924),
.Y(n_1543)
);

CKINVDCx16_ASAP7_75t_R g1544 ( 
.A(n_796),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_326),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_436),
.Y(n_1546)
);

CKINVDCx14_ASAP7_75t_R g1547 ( 
.A(n_713),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1041),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_956),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1005),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_131),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_758),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_375),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1134),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1268),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1163),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_408),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1142),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1187),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_247),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_569),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_816),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_996),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_522),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_282),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_249),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_495),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_582),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1170),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_321),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_20),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1091),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_793),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1277),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_310),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_266),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1177),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_492),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_787),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1011),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1113),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_998),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_760),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1225),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1034),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_807),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1095),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_430),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_74),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_481),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_688),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_193),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_348),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1263),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_29),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_776),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_757),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1165),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_775),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1021),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1241),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_850),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_105),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1060),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_497),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_185),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_396),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_837),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_999),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_182),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_920),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1050),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1250),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1273),
.Y(n_1614)
);

BUFx10_ASAP7_75t_L g1615 ( 
.A(n_780),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_497),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_158),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1084),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1160),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_969),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_211),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_962),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_162),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_979),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_982),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_409),
.Y(n_1626)
);

CKINVDCx16_ASAP7_75t_R g1627 ( 
.A(n_1249),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_735),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_255),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1146),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_955),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1246),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_483),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1022),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1186),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1032),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_383),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_222),
.Y(n_1638)
);

CKINVDCx20_ASAP7_75t_R g1639 ( 
.A(n_121),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_59),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_190),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_508),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1000),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1228),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1220),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_486),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_342),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_204),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1015),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_238),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1013),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1048),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1196),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_707),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1139),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_811),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_515),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_462),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_103),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_561),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_593),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_549),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1198),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1178),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1203),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_618),
.Y(n_1666)
);

CKINVDCx20_ASAP7_75t_R g1667 ( 
.A(n_745),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_994),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_806),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_715),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_626),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1248),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1036),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_959),
.Y(n_1674)
);

BUFx10_ASAP7_75t_L g1675 ( 
.A(n_980),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_213),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_370),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_9),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_83),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_149),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_514),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1154),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_385),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1236),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_594),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_950),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_15),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_299),
.Y(n_1688)
);

CKINVDCx20_ASAP7_75t_R g1689 ( 
.A(n_90),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1183),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_225),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_447),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_633),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_137),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_959),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_740),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1033),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_111),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_970),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1169),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_872),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_88),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1286),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1256),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_465),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1194),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_972),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_401),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_353),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_437),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_707),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_395),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1245),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_161),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_59),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_906),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1270),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1152),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_374),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1278),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_995),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_949),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1252),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1126),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_983),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1022),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_261),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_586),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1175),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_736),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_986),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_947),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1174),
.Y(n_1733)
);

INVxp67_ASAP7_75t_SL g1734 ( 
.A(n_883),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_565),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_456),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_595),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_3),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_810),
.Y(n_1739)
);

CKINVDCx14_ASAP7_75t_R g1740 ( 
.A(n_595),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_317),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1185),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1016),
.Y(n_1743)
);

CKINVDCx20_ASAP7_75t_R g1744 ( 
.A(n_81),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_240),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_322),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_962),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1131),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1229),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_997),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1124),
.Y(n_1751)
);

CKINVDCx20_ASAP7_75t_R g1752 ( 
.A(n_827),
.Y(n_1752)
);

CKINVDCx16_ASAP7_75t_R g1753 ( 
.A(n_1012),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_891),
.Y(n_1754)
);

BUFx10_ASAP7_75t_L g1755 ( 
.A(n_1193),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_656),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1092),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_785),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_52),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_256),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_502),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_284),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_268),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_578),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1151),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_875),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1137),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_965),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1280),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_895),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_223),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1226),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_917),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1020),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_26),
.Y(n_1775)
);

CKINVDCx16_ASAP7_75t_R g1776 ( 
.A(n_677),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_667),
.Y(n_1777)
);

BUFx3_ASAP7_75t_L g1778 ( 
.A(n_463),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1067),
.Y(n_1779)
);

CKINVDCx20_ASAP7_75t_R g1780 ( 
.A(n_541),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_292),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1168),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_855),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_339),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_314),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_268),
.Y(n_1786)
);

CKINVDCx16_ASAP7_75t_R g1787 ( 
.A(n_984),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_614),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_332),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1264),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_630),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1156),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_408),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_466),
.Y(n_1794)
);

BUFx10_ASAP7_75t_L g1795 ( 
.A(n_1129),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_751),
.Y(n_1796)
);

CKINVDCx20_ASAP7_75t_R g1797 ( 
.A(n_261),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_470),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_1244),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1147),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_714),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1122),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1030),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_947),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_666),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1121),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1089),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_56),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_153),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_583),
.Y(n_1810)
);

CKINVDCx20_ASAP7_75t_R g1811 ( 
.A(n_963),
.Y(n_1811)
);

BUFx3_ASAP7_75t_L g1812 ( 
.A(n_1189),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_217),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_968),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1153),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1276),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_306),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_389),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_463),
.Y(n_1819)
);

CKINVDCx20_ASAP7_75t_R g1820 ( 
.A(n_991),
.Y(n_1820)
);

CKINVDCx20_ASAP7_75t_R g1821 ( 
.A(n_1218),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_546),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1231),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1027),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_628),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1054),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_887),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_865),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_885),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1180),
.Y(n_1830)
);

CKINVDCx20_ASAP7_75t_R g1831 ( 
.A(n_863),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1240),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_943),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_126),
.Y(n_1834)
);

CKINVDCx20_ASAP7_75t_R g1835 ( 
.A(n_432),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_255),
.Y(n_1836)
);

CKINVDCx20_ASAP7_75t_R g1837 ( 
.A(n_68),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_390),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_674),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1004),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_977),
.Y(n_1841)
);

BUFx10_ASAP7_75t_L g1842 ( 
.A(n_576),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_531),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_868),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_917),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_985),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_7),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_419),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_424),
.Y(n_1849)
);

BUFx3_ASAP7_75t_L g1850 ( 
.A(n_314),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_801),
.Y(n_1851)
);

BUFx3_ASAP7_75t_L g1852 ( 
.A(n_4),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1101),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_756),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_60),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1021),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_415),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_838),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1221),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_634),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_60),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1254),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_961),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_679),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1023),
.Y(n_1865)
);

CKINVDCx20_ASAP7_75t_R g1866 ( 
.A(n_605),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1053),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1191),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_611),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1029),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_245),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_686),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_286),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_964),
.Y(n_1874)
);

BUFx3_ASAP7_75t_L g1875 ( 
.A(n_1001),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_172),
.Y(n_1876)
);

BUFx6f_ASAP7_75t_L g1877 ( 
.A(n_1051),
.Y(n_1877)
);

BUFx10_ASAP7_75t_L g1878 ( 
.A(n_902),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_841),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_259),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1258),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1078),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_620),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_910),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_180),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_690),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_969),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_613),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_524),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_1284),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_28),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_208),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1143),
.Y(n_1893)
);

CKINVDCx20_ASAP7_75t_R g1894 ( 
.A(n_1148),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1288),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_486),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_457),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_28),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_35),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_575),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_263),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_630),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1052),
.Y(n_1903)
);

BUFx10_ASAP7_75t_L g1904 ( 
.A(n_1096),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1213),
.Y(n_1905)
);

CKINVDCx20_ASAP7_75t_R g1906 ( 
.A(n_1042),
.Y(n_1906)
);

BUFx3_ASAP7_75t_L g1907 ( 
.A(n_832),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1076),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1261),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_41),
.Y(n_1910)
);

CKINVDCx14_ASAP7_75t_R g1911 ( 
.A(n_391),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1200),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_973),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1232),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_896),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_421),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_950),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1206),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_682),
.Y(n_1919)
);

CKINVDCx20_ASAP7_75t_R g1920 ( 
.A(n_1049),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_930),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_971),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_210),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1045),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_107),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_951),
.Y(n_1926)
);

CKINVDCx20_ASAP7_75t_R g1927 ( 
.A(n_963),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_173),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1003),
.Y(n_1929)
);

CKINVDCx20_ASAP7_75t_R g1930 ( 
.A(n_695),
.Y(n_1930)
);

BUFx2_ASAP7_75t_L g1931 ( 
.A(n_535),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_480),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_365),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_L g1934 ( 
.A(n_585),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_758),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_333),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_967),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_88),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_885),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1238),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_297),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1038),
.Y(n_1942)
);

CKINVDCx16_ASAP7_75t_R g1943 ( 
.A(n_20),
.Y(n_1943)
);

BUFx6f_ASAP7_75t_L g1944 ( 
.A(n_209),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1128),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_273),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_713),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_35),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1275),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1138),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1127),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1233),
.Y(n_1952)
);

INVxp67_ASAP7_75t_SL g1953 ( 
.A(n_625),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_636),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_967),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_590),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1069),
.Y(n_1957)
);

CKINVDCx20_ASAP7_75t_R g1958 ( 
.A(n_1224),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_403),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_733),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_984),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_1028),
.Y(n_1962)
);

CKINVDCx5p33_ASAP7_75t_R g1963 ( 
.A(n_184),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_753),
.Y(n_1964)
);

BUFx3_ASAP7_75t_L g1965 ( 
.A(n_1271),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_638),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1049),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1130),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1285),
.Y(n_1969)
);

BUFx10_ASAP7_75t_L g1970 ( 
.A(n_784),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_302),
.Y(n_1971)
);

CKINVDCx20_ASAP7_75t_R g1972 ( 
.A(n_881),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_876),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1164),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1017),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1190),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_636),
.Y(n_1977)
);

INVx1_ASAP7_75t_SL g1978 ( 
.A(n_1287),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_472),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_70),
.Y(n_1980)
);

CKINVDCx20_ASAP7_75t_R g1981 ( 
.A(n_122),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_1243),
.Y(n_1982)
);

CKINVDCx20_ASAP7_75t_R g1983 ( 
.A(n_165),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_485),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1230),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1039),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_942),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_1181),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_229),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_124),
.Y(n_1990)
);

BUFx5_ASAP7_75t_L g1991 ( 
.A(n_857),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_424),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_875),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_847),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_24),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1274),
.Y(n_1996)
);

CKINVDCx20_ASAP7_75t_R g1997 ( 
.A(n_955),
.Y(n_1997)
);

BUFx10_ASAP7_75t_L g1998 ( 
.A(n_249),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_992),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1052),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_1237),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1123),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_92),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_493),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_650),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_193),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_481),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_981),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_448),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_102),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_24),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_861),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_5),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_688),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_554),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_402),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1007),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_623),
.Y(n_2018)
);

CKINVDCx14_ASAP7_75t_R g2019 ( 
.A(n_1204),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_669),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_711),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_865),
.Y(n_2022)
);

BUFx3_ASAP7_75t_L g2023 ( 
.A(n_294),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1135),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_175),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1141),
.Y(n_2026)
);

INVxp67_ASAP7_75t_L g2027 ( 
.A(n_954),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_575),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_558),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_810),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_907),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_581),
.Y(n_2032)
);

INVx1_ASAP7_75t_SL g2033 ( 
.A(n_1182),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_73),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1159),
.Y(n_2035)
);

BUFx3_ASAP7_75t_L g2036 ( 
.A(n_1235),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_161),
.Y(n_2037)
);

BUFx5_ASAP7_75t_L g2038 ( 
.A(n_976),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_555),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_115),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_695),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_654),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_163),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_975),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_951),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_351),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_492),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_131),
.Y(n_2048)
);

BUFx3_ASAP7_75t_L g2049 ( 
.A(n_446),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1040),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1044),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_645),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_563),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_70),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_470),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_422),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_515),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_443),
.Y(n_2058)
);

BUFx10_ASAP7_75t_L g2059 ( 
.A(n_952),
.Y(n_2059)
);

BUFx3_ASAP7_75t_L g2060 ( 
.A(n_958),
.Y(n_2060)
);

INVxp67_ASAP7_75t_L g2061 ( 
.A(n_114),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1265),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_578),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_1145),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1133),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_340),
.Y(n_2066)
);

CKINVDCx20_ASAP7_75t_R g2067 ( 
.A(n_1008),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1251),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_94),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_773),
.Y(n_2070)
);

BUFx6f_ASAP7_75t_L g2071 ( 
.A(n_26),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_800),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1112),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_180),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_221),
.Y(n_2075)
);

CKINVDCx20_ASAP7_75t_R g2076 ( 
.A(n_676),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_944),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_41),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_465),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_248),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1006),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_120),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_656),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_464),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_129),
.Y(n_2085)
);

CKINVDCx14_ASAP7_75t_R g2086 ( 
.A(n_767),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_725),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_819),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_1219),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_162),
.Y(n_2090)
);

CKINVDCx20_ASAP7_75t_R g2091 ( 
.A(n_1064),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1296),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1296),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1296),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1394),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1296),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1296),
.Y(n_2097)
);

CKINVDCx5p33_ASAP7_75t_R g2098 ( 
.A(n_1369),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1991),
.Y(n_2099)
);

INVxp67_ASAP7_75t_SL g2100 ( 
.A(n_1524),
.Y(n_2100)
);

INVxp33_ASAP7_75t_L g2101 ( 
.A(n_1311),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1991),
.Y(n_2102)
);

CKINVDCx20_ASAP7_75t_R g2103 ( 
.A(n_1331),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1991),
.Y(n_2104)
);

BUFx3_ASAP7_75t_L g2105 ( 
.A(n_1541),
.Y(n_2105)
);

INVxp33_ASAP7_75t_L g2106 ( 
.A(n_1338),
.Y(n_2106)
);

INVxp67_ASAP7_75t_L g2107 ( 
.A(n_1585),
.Y(n_2107)
);

CKINVDCx14_ASAP7_75t_R g2108 ( 
.A(n_1290),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1991),
.Y(n_2109)
);

INVxp33_ASAP7_75t_SL g2110 ( 
.A(n_1605),
.Y(n_2110)
);

BUFx3_ASAP7_75t_L g2111 ( 
.A(n_1541),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1991),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_1341),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2038),
.Y(n_2114)
);

INVxp67_ASAP7_75t_L g2115 ( 
.A(n_1697),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_1544),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2038),
.Y(n_2117)
);

CKINVDCx20_ASAP7_75t_R g2118 ( 
.A(n_2091),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2038),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2038),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2038),
.Y(n_2121)
);

INVxp33_ASAP7_75t_SL g2122 ( 
.A(n_1699),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1524),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1341),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1341),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_1298),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1421),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1421),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1421),
.Y(n_2129)
);

BUFx2_ASAP7_75t_L g2130 ( 
.A(n_1756),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1485),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1485),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1485),
.Y(n_2133)
);

INVxp67_ASAP7_75t_SL g2134 ( 
.A(n_1316),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1505),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1505),
.Y(n_2136)
);

INVxp67_ASAP7_75t_L g2137 ( 
.A(n_1931),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1307),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1505),
.Y(n_2139)
);

INVxp67_ASAP7_75t_SL g2140 ( 
.A(n_1321),
.Y(n_2140)
);

CKINVDCx16_ASAP7_75t_R g2141 ( 
.A(n_1753),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1532),
.Y(n_2142)
);

INVxp67_ASAP7_75t_SL g2143 ( 
.A(n_1508),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1532),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1532),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1580),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1580),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1318),
.Y(n_2148)
);

INVxp33_ASAP7_75t_L g2149 ( 
.A(n_1962),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1580),
.Y(n_2150)
);

CKINVDCx20_ASAP7_75t_R g2151 ( 
.A(n_1461),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1588),
.Y(n_2152)
);

INVxp33_ASAP7_75t_SL g2153 ( 
.A(n_1289),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1588),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1588),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_1547),
.B(n_1),
.Y(n_2156)
);

INVxp33_ASAP7_75t_L g2157 ( 
.A(n_1294),
.Y(n_2157)
);

INVxp67_ASAP7_75t_L g2158 ( 
.A(n_1292),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1636),
.Y(n_2159)
);

BUFx3_ASAP7_75t_L g2160 ( 
.A(n_1755),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_1636),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1636),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1711),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1711),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1711),
.Y(n_2165)
);

INVxp67_ASAP7_75t_SL g2166 ( 
.A(n_1802),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1745),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1745),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1745),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1813),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1813),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1813),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1825),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1825),
.Y(n_2174)
);

INVxp67_ASAP7_75t_L g2175 ( 
.A(n_1292),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1825),
.Y(n_2176)
);

CKINVDCx16_ASAP7_75t_R g2177 ( 
.A(n_1776),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1877),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1877),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1877),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1926),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_1319),
.Y(n_2182)
);

INVxp67_ASAP7_75t_L g2183 ( 
.A(n_1312),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1926),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1926),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1934),
.Y(n_2186)
);

BUFx3_ASAP7_75t_L g2187 ( 
.A(n_1755),
.Y(n_2187)
);

INVxp67_ASAP7_75t_SL g2188 ( 
.A(n_1812),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1934),
.Y(n_2189)
);

BUFx2_ASAP7_75t_L g2190 ( 
.A(n_1740),
.Y(n_2190)
);

INVx2_ASAP7_75t_SL g2191 ( 
.A(n_1312),
.Y(n_2191)
);

INVxp67_ASAP7_75t_SL g2192 ( 
.A(n_1895),
.Y(n_2192)
);

INVxp33_ASAP7_75t_SL g2193 ( 
.A(n_1295),
.Y(n_2193)
);

INVxp67_ASAP7_75t_SL g2194 ( 
.A(n_1965),
.Y(n_2194)
);

CKINVDCx16_ASAP7_75t_R g2195 ( 
.A(n_1787),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1934),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1320),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_1328),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1944),
.Y(n_2199)
);

INVxp67_ASAP7_75t_L g2200 ( 
.A(n_1363),
.Y(n_2200)
);

INVxp67_ASAP7_75t_L g2201 ( 
.A(n_1363),
.Y(n_2201)
);

INVxp33_ASAP7_75t_SL g2202 ( 
.A(n_1304),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1944),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_1332),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1944),
.Y(n_2205)
);

INVx1_ASAP7_75t_SL g2206 ( 
.A(n_1291),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1987),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1987),
.Y(n_2208)
);

CKINVDCx20_ASAP7_75t_R g2209 ( 
.A(n_1477),
.Y(n_2209)
);

XOR2xp5_ASAP7_75t_L g2210 ( 
.A(n_1911),
.B(n_0),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1987),
.Y(n_2211)
);

CKINVDCx20_ASAP7_75t_R g2212 ( 
.A(n_1587),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2003),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2003),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2003),
.Y(n_2215)
);

CKINVDCx20_ASAP7_75t_R g2216 ( 
.A(n_1635),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2071),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2071),
.Y(n_2218)
);

INVxp67_ASAP7_75t_SL g2219 ( 
.A(n_2036),
.Y(n_2219)
);

INVx1_ASAP7_75t_SL g2220 ( 
.A(n_1667),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2071),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1382),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1387),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1450),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1543),
.Y(n_2225)
);

NOR2xp67_ASAP7_75t_L g2226 ( 
.A(n_1327),
.B(n_0),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1293),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1646),
.Y(n_2228)
);

INVxp67_ASAP7_75t_SL g2229 ( 
.A(n_1451),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1739),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1746),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1778),
.Y(n_2232)
);

CKINVDCx5p33_ASAP7_75t_R g2233 ( 
.A(n_1334),
.Y(n_2233)
);

BUFx2_ASAP7_75t_L g2234 ( 
.A(n_2086),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1850),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1293),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1852),
.Y(n_2237)
);

INVxp67_ASAP7_75t_SL g2238 ( 
.A(n_1862),
.Y(n_2238)
);

BUFx2_ASAP7_75t_L g2239 ( 
.A(n_1874),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1875),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_1394),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1907),
.Y(n_2242)
);

INVxp33_ASAP7_75t_SL g2243 ( 
.A(n_1308),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2023),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_1349),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2049),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2060),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1293),
.Y(n_2248)
);

INVxp67_ASAP7_75t_SL g2249 ( 
.A(n_1945),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2090),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1299),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1300),
.Y(n_2252)
);

INVxp67_ASAP7_75t_L g2253 ( 
.A(n_1438),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2074),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2075),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2081),
.Y(n_2256)
);

INVxp67_ASAP7_75t_SL g2257 ( 
.A(n_1330),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2135),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2159),
.Y(n_2259)
);

INVx4_ASAP7_75t_L g2260 ( 
.A(n_2126),
.Y(n_2260)
);

BUFx3_ASAP7_75t_L g2261 ( 
.A(n_2239),
.Y(n_2261)
);

OA22x2_ASAP7_75t_SL g2262 ( 
.A1(n_2210),
.A2(n_1953),
.B1(n_1734),
.B2(n_1305),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2138),
.B(n_2019),
.Y(n_2263)
);

BUFx3_ASAP7_75t_L g2264 ( 
.A(n_2222),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2168),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2185),
.Y(n_2266)
);

BUFx6f_ASAP7_75t_L g2267 ( 
.A(n_2199),
.Y(n_2267)
);

CKINVDCx8_ASAP7_75t_R g2268 ( 
.A(n_2141),
.Y(n_2268)
);

OA21x2_ASAP7_75t_L g2269 ( 
.A1(n_2092),
.A2(n_1392),
.B(n_1367),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_2190),
.B(n_1385),
.Y(n_2270)
);

BUFx8_ASAP7_75t_SL g2271 ( 
.A(n_2098),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2217),
.Y(n_2272)
);

OAI22x1_ASAP7_75t_SL g2273 ( 
.A1(n_2110),
.A2(n_1370),
.B1(n_1411),
.B2(n_1362),
.Y(n_2273)
);

OAI22x1_ASAP7_75t_R g2274 ( 
.A1(n_2103),
.A2(n_1516),
.B1(n_1538),
.B2(n_1432),
.Y(n_2274)
);

OAI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2122),
.A2(n_1943),
.B1(n_1502),
.B2(n_1530),
.Y(n_2275)
);

INVx3_ASAP7_75t_L g2276 ( 
.A(n_2113),
.Y(n_2276)
);

INVx5_ASAP7_75t_L g2277 ( 
.A(n_2191),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2124),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2125),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2148),
.B(n_1351),
.Y(n_2280)
);

AOI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2156),
.A2(n_1627),
.B1(n_1445),
.B2(n_1821),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2095),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2127),
.Y(n_2283)
);

OA21x2_ASAP7_75t_L g2284 ( 
.A1(n_2093),
.A2(n_1403),
.B(n_1399),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_2095),
.Y(n_2285)
);

BUFx6f_ASAP7_75t_L g2286 ( 
.A(n_2095),
.Y(n_2286)
);

INVx5_ASAP7_75t_L g2287 ( 
.A(n_2113),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2128),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_L g2289 ( 
.A(n_2153),
.B(n_1408),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2241),
.Y(n_2290)
);

INVx5_ASAP7_75t_L g2291 ( 
.A(n_2241),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2129),
.Y(n_2292)
);

INVx5_ASAP7_75t_L g2293 ( 
.A(n_2161),
.Y(n_2293)
);

BUFx8_ASAP7_75t_L g2294 ( 
.A(n_2234),
.Y(n_2294)
);

INVx3_ASAP7_75t_L g2295 ( 
.A(n_2161),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2182),
.B(n_1381),
.Y(n_2296)
);

BUFx3_ASAP7_75t_L g2297 ( 
.A(n_2223),
.Y(n_2297)
);

AOI22xp5_ASAP7_75t_L g2298 ( 
.A1(n_2177),
.A2(n_1918),
.B1(n_1958),
.B2(n_1894),
.Y(n_2298)
);

BUFx6f_ASAP7_75t_L g2299 ( 
.A(n_2241),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_2131),
.Y(n_2300)
);

AND2x4_ASAP7_75t_L g2301 ( 
.A(n_2105),
.B(n_1830),
.Y(n_2301)
);

BUFx12f_ASAP7_75t_L g2302 ( 
.A(n_2197),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2195),
.A2(n_2115),
.B1(n_2137),
.B2(n_2107),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2132),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2133),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2198),
.B(n_1427),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2204),
.B(n_1598),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2108),
.B(n_1795),
.Y(n_2308)
);

CKINVDCx16_ASAP7_75t_R g2309 ( 
.A(n_2118),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2136),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_2116),
.B(n_1303),
.Y(n_2311)
);

BUFx3_ASAP7_75t_L g2312 ( 
.A(n_2224),
.Y(n_2312)
);

OAI22x1_ASAP7_75t_R g2313 ( 
.A1(n_2151),
.A2(n_1597),
.B1(n_1629),
.B2(n_1576),
.Y(n_2313)
);

OA21x2_ASAP7_75t_L g2314 ( 
.A1(n_2094),
.A2(n_1498),
.B(n_1484),
.Y(n_2314)
);

BUFx6f_ASAP7_75t_L g2315 ( 
.A(n_2139),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2142),
.Y(n_2316)
);

BUFx6f_ASAP7_75t_L g2317 ( 
.A(n_2144),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2233),
.B(n_1614),
.Y(n_2318)
);

BUFx3_ASAP7_75t_L g2319 ( 
.A(n_2225),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2193),
.B(n_1968),
.Y(n_2320)
);

AND2x2_ASAP7_75t_SL g2321 ( 
.A(n_2130),
.B(n_1302),
.Y(n_2321)
);

HB1xp67_ASAP7_75t_L g2322 ( 
.A(n_2111),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2245),
.B(n_1723),
.Y(n_2323)
);

BUFx3_ASAP7_75t_L g2324 ( 
.A(n_2228),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2145),
.Y(n_2325)
);

OAI22xp5_ASAP7_75t_L g2326 ( 
.A1(n_2149),
.A2(n_1519),
.B1(n_2027),
.B2(n_1468),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2146),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2147),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_2202),
.B(n_1978),
.Y(n_2329)
);

BUFx6f_ASAP7_75t_L g2330 ( 
.A(n_2150),
.Y(n_2330)
);

OAI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2101),
.A2(n_2061),
.B1(n_1314),
.B2(n_1315),
.Y(n_2331)
);

BUFx12f_ASAP7_75t_L g2332 ( 
.A(n_2160),
.Y(n_2332)
);

BUFx8_ASAP7_75t_SL g2333 ( 
.A(n_2209),
.Y(n_2333)
);

AND2x6_ASAP7_75t_L g2334 ( 
.A(n_2187),
.B(n_1352),
.Y(n_2334)
);

HB1xp67_ASAP7_75t_L g2335 ( 
.A(n_2206),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2152),
.Y(n_2336)
);

OAI21x1_ASAP7_75t_L g2337 ( 
.A1(n_2096),
.A2(n_1301),
.B(n_1297),
.Y(n_2337)
);

BUFx6f_ASAP7_75t_L g2338 ( 
.A(n_2154),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2155),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2162),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_2134),
.B(n_1795),
.Y(n_2341)
);

INVx4_ASAP7_75t_L g2342 ( 
.A(n_2097),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2163),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2164),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_2165),
.Y(n_2345)
);

BUFx2_ASAP7_75t_L g2346 ( 
.A(n_2158),
.Y(n_2346)
);

OAI22x1_ASAP7_75t_SL g2347 ( 
.A1(n_2220),
.A2(n_1676),
.B1(n_1677),
.B2(n_1639),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2167),
.Y(n_2348)
);

HB1xp67_ASAP7_75t_L g2349 ( 
.A(n_2175),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_2183),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2169),
.Y(n_2351)
);

HB1xp67_ASAP7_75t_L g2352 ( 
.A(n_2200),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2170),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2171),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2172),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2173),
.Y(n_2356)
);

BUFx6f_ASAP7_75t_L g2357 ( 
.A(n_2174),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2176),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2178),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2179),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2180),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2181),
.Y(n_2362)
);

OA21x2_ASAP7_75t_L g2363 ( 
.A1(n_2099),
.A2(n_1536),
.B(n_1503),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2184),
.Y(n_2364)
);

BUFx6f_ASAP7_75t_L g2365 ( 
.A(n_2186),
.Y(n_2365)
);

AND2x4_ASAP7_75t_L g2366 ( 
.A(n_2140),
.B(n_2033),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2143),
.B(n_2166),
.Y(n_2367)
);

CKINVDCx5p33_ASAP7_75t_R g2368 ( 
.A(n_2212),
.Y(n_2368)
);

OAI22xp33_ASAP7_75t_SL g2369 ( 
.A1(n_2100),
.A2(n_1418),
.B1(n_1456),
.B2(n_1374),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2189),
.Y(n_2370)
);

HB1xp67_ASAP7_75t_L g2371 ( 
.A(n_2201),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2196),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2188),
.B(n_1951),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2203),
.Y(n_2374)
);

BUFx6f_ASAP7_75t_L g2375 ( 
.A(n_2205),
.Y(n_2375)
);

BUFx6f_ASAP7_75t_L g2376 ( 
.A(n_2207),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2208),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2211),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2213),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2214),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_2215),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2218),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_2253),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_L g2384 ( 
.A(n_2243),
.B(n_1952),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2221),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2192),
.B(n_1904),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_2106),
.B(n_1904),
.Y(n_2387)
);

BUFx3_ASAP7_75t_L g2388 ( 
.A(n_2230),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2102),
.Y(n_2389)
);

CKINVDCx6p67_ASAP7_75t_R g2390 ( 
.A(n_2216),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2104),
.Y(n_2391)
);

CKINVDCx16_ASAP7_75t_R g2392 ( 
.A(n_2231),
.Y(n_2392)
);

AND2x4_ASAP7_75t_L g2393 ( 
.A(n_2194),
.B(n_1555),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_2219),
.B(n_1556),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2109),
.Y(n_2395)
);

BUFx6f_ASAP7_75t_L g2396 ( 
.A(n_2250),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_2251),
.Y(n_2397)
);

INVx5_ASAP7_75t_L g2398 ( 
.A(n_2227),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2112),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2114),
.Y(n_2400)
);

OR2x2_ASAP7_75t_L g2401 ( 
.A(n_2232),
.B(n_1398),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2117),
.Y(n_2402)
);

AND2x4_ASAP7_75t_L g2403 ( 
.A(n_2229),
.B(n_1584),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_2238),
.B(n_1594),
.Y(n_2404)
);

BUFx6f_ASAP7_75t_L g2405 ( 
.A(n_2252),
.Y(n_2405)
);

OAI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2249),
.A2(n_1325),
.B1(n_1326),
.B2(n_1310),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_2257),
.Y(n_2407)
);

BUFx6f_ASAP7_75t_L g2408 ( 
.A(n_2254),
.Y(n_2408)
);

AND2x6_ASAP7_75t_L g2409 ( 
.A(n_2235),
.B(n_1553),
.Y(n_2409)
);

AOI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2226),
.A2(n_1333),
.B1(n_1335),
.B2(n_1329),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2237),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2119),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2157),
.B(n_1460),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2240),
.B(n_2242),
.Y(n_2414)
);

OAI21x1_ASAP7_75t_L g2415 ( 
.A1(n_2236),
.A2(n_1462),
.B(n_1378),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2120),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2121),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2255),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2123),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2256),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2248),
.Y(n_2421)
);

BUFx6f_ASAP7_75t_L g2422 ( 
.A(n_2244),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2246),
.B(n_1604),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2247),
.Y(n_2424)
);

OAI22x1_ASAP7_75t_R g2425 ( 
.A1(n_2103),
.A2(n_1744),
.B1(n_1752),
.B2(n_1689),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2108),
.B(n_1471),
.Y(n_2426)
);

CKINVDCx16_ASAP7_75t_R g2427 ( 
.A(n_2141),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2135),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2135),
.Y(n_2429)
);

BUFx8_ASAP7_75t_SL g2430 ( 
.A(n_2098),
.Y(n_2430)
);

OA21x2_ASAP7_75t_L g2431 ( 
.A1(n_2092),
.A2(n_1619),
.B(n_1618),
.Y(n_2431)
);

BUFx6f_ASAP7_75t_L g2432 ( 
.A(n_2135),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_2190),
.B(n_1644),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2126),
.B(n_1782),
.Y(n_2434)
);

BUFx3_ASAP7_75t_L g2435 ( 
.A(n_2239),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_2153),
.B(n_1655),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_2153),
.B(n_1665),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2116),
.Y(n_2438)
);

BUFx6f_ASAP7_75t_L g2439 ( 
.A(n_2135),
.Y(n_2439)
);

OAI21x1_ASAP7_75t_L g2440 ( 
.A1(n_2096),
.A2(n_1682),
.B(n_1672),
.Y(n_2440)
);

OA21x2_ASAP7_75t_L g2441 ( 
.A1(n_2092),
.A2(n_1704),
.B(n_1703),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2135),
.Y(n_2442)
);

BUFx6f_ASAP7_75t_L g2443 ( 
.A(n_2135),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2108),
.B(n_1533),
.Y(n_2444)
);

BUFx6f_ASAP7_75t_L g2445 ( 
.A(n_2135),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2135),
.Y(n_2446)
);

INVx5_ASAP7_75t_L g2447 ( 
.A(n_2191),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2126),
.B(n_1706),
.Y(n_2448)
);

BUFx8_ASAP7_75t_L g2449 ( 
.A(n_2190),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2135),
.Y(n_2450)
);

BUFx6f_ASAP7_75t_L g2451 ( 
.A(n_2135),
.Y(n_2451)
);

BUFx6f_ASAP7_75t_L g2452 ( 
.A(n_2135),
.Y(n_2452)
);

BUFx8_ASAP7_75t_SL g2453 ( 
.A(n_2098),
.Y(n_2453)
);

INVx2_ASAP7_75t_SL g2454 ( 
.A(n_2105),
.Y(n_2454)
);

BUFx6f_ASAP7_75t_L g2455 ( 
.A(n_2135),
.Y(n_2455)
);

AND2x6_ASAP7_75t_L g2456 ( 
.A(n_2156),
.B(n_1571),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_2135),
.Y(n_2457)
);

HB1xp67_ASAP7_75t_L g2458 ( 
.A(n_2116),
.Y(n_2458)
);

BUFx6f_ASAP7_75t_L g2459 ( 
.A(n_2135),
.Y(n_2459)
);

BUFx6f_ASAP7_75t_L g2460 ( 
.A(n_2135),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2135),
.Y(n_2461)
);

AND2x4_ASAP7_75t_L g2462 ( 
.A(n_2190),
.B(n_1718),
.Y(n_2462)
);

INVx4_ASAP7_75t_L g2463 ( 
.A(n_2126),
.Y(n_2463)
);

AOI22x1_ASAP7_75t_SL g2464 ( 
.A1(n_2103),
.A2(n_1780),
.B1(n_1797),
.B2(n_1771),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2135),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_SL g2466 ( 
.A(n_2190),
.B(n_1438),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2135),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2135),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2135),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2135),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2190),
.B(n_1765),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_L g2472 ( 
.A(n_2135),
.Y(n_2472)
);

BUFx6f_ASAP7_75t_L g2473 ( 
.A(n_2135),
.Y(n_2473)
);

BUFx6f_ASAP7_75t_L g2474 ( 
.A(n_2135),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2135),
.Y(n_2475)
);

OAI22xp5_ASAP7_75t_L g2476 ( 
.A1(n_2110),
.A2(n_1339),
.B1(n_1340),
.B2(n_1337),
.Y(n_2476)
);

CKINVDCx11_ASAP7_75t_R g2477 ( 
.A(n_2103),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2135),
.Y(n_2478)
);

HB1xp67_ASAP7_75t_L g2479 ( 
.A(n_2116),
.Y(n_2479)
);

BUFx2_ASAP7_75t_L g2480 ( 
.A(n_2108),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2135),
.Y(n_2481)
);

NOR2x1_ASAP7_75t_L g2482 ( 
.A(n_2105),
.B(n_1767),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2135),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2135),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_2126),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2135),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2135),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2135),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2135),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2126),
.B(n_1823),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2135),
.Y(n_2491)
);

BUFx3_ASAP7_75t_L g2492 ( 
.A(n_2239),
.Y(n_2492)
);

BUFx2_ASAP7_75t_L g2493 ( 
.A(n_2108),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2135),
.Y(n_2494)
);

BUFx3_ASAP7_75t_L g2495 ( 
.A(n_2239),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2135),
.Y(n_2496)
);

BUFx6f_ASAP7_75t_L g2497 ( 
.A(n_2135),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2135),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2135),
.Y(n_2499)
);

BUFx6f_ASAP7_75t_L g2500 ( 
.A(n_2135),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2135),
.Y(n_2501)
);

BUFx6f_ASAP7_75t_L g2502 ( 
.A(n_2135),
.Y(n_2502)
);

INVx5_ASAP7_75t_L g2503 ( 
.A(n_2191),
.Y(n_2503)
);

BUFx3_ASAP7_75t_L g2504 ( 
.A(n_2239),
.Y(n_2504)
);

BUFx2_ASAP7_75t_L g2505 ( 
.A(n_2108),
.Y(n_2505)
);

BUFx12f_ASAP7_75t_L g2506 ( 
.A(n_2098),
.Y(n_2506)
);

HB1xp67_ASAP7_75t_L g2507 ( 
.A(n_2116),
.Y(n_2507)
);

INVx5_ASAP7_75t_L g2508 ( 
.A(n_2191),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2135),
.Y(n_2509)
);

OAI22xp5_ASAP7_75t_R g2510 ( 
.A1(n_2110),
.A2(n_1343),
.B1(n_1344),
.B2(n_1342),
.Y(n_2510)
);

BUFx3_ASAP7_75t_L g2511 ( 
.A(n_2239),
.Y(n_2511)
);

BUFx6f_ASAP7_75t_L g2512 ( 
.A(n_2135),
.Y(n_2512)
);

OAI22x1_ASAP7_75t_L g2513 ( 
.A1(n_2210),
.A2(n_1595),
.B1(n_1649),
.B2(n_1607),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2135),
.Y(n_2514)
);

AND2x4_ASAP7_75t_L g2515 ( 
.A(n_2190),
.B(n_1832),
.Y(n_2515)
);

BUFx6f_ASAP7_75t_L g2516 ( 
.A(n_2135),
.Y(n_2516)
);

INVx6_ASAP7_75t_L g2517 ( 
.A(n_2105),
.Y(n_2517)
);

CKINVDCx16_ASAP7_75t_R g2518 ( 
.A(n_2141),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2135),
.Y(n_2519)
);

BUFx6f_ASAP7_75t_L g2520 ( 
.A(n_2135),
.Y(n_2520)
);

CKINVDCx6p67_ASAP7_75t_R g2521 ( 
.A(n_2141),
.Y(n_2521)
);

AND2x4_ASAP7_75t_L g2522 ( 
.A(n_2190),
.B(n_1908),
.Y(n_2522)
);

INVx5_ASAP7_75t_L g2523 ( 
.A(n_2191),
.Y(n_2523)
);

BUFx6f_ASAP7_75t_L g2524 ( 
.A(n_2135),
.Y(n_2524)
);

AND2x2_ASAP7_75t_SL g2525 ( 
.A(n_2141),
.B(n_1360),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_L g2526 ( 
.A(n_2153),
.B(n_1909),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2135),
.Y(n_2527)
);

OAI22xp5_ASAP7_75t_L g2528 ( 
.A1(n_2110),
.A2(n_1346),
.B1(n_1347),
.B2(n_1345),
.Y(n_2528)
);

OAI21x1_ASAP7_75t_L g2529 ( 
.A1(n_2096),
.A2(n_1940),
.B(n_1914),
.Y(n_2529)
);

INVxp33_ASAP7_75t_SL g2530 ( 
.A(n_2210),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2135),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2135),
.Y(n_2532)
);

AND2x4_ASAP7_75t_L g2533 ( 
.A(n_2190),
.B(n_1949),
.Y(n_2533)
);

INVx5_ASAP7_75t_L g2534 ( 
.A(n_2191),
.Y(n_2534)
);

INVx5_ASAP7_75t_L g2535 ( 
.A(n_2191),
.Y(n_2535)
);

BUFx6f_ASAP7_75t_L g2536 ( 
.A(n_2135),
.Y(n_2536)
);

BUFx12f_ASAP7_75t_L g2537 ( 
.A(n_2098),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2135),
.Y(n_2538)
);

BUFx6f_ASAP7_75t_L g2539 ( 
.A(n_2135),
.Y(n_2539)
);

AOI22xp5_ASAP7_75t_L g2540 ( 
.A1(n_2110),
.A2(n_1350),
.B1(n_1353),
.B2(n_1348),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2108),
.B(n_1564),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2108),
.B(n_1637),
.Y(n_2542)
);

BUFx12f_ASAP7_75t_L g2543 ( 
.A(n_2098),
.Y(n_2543)
);

INVx3_ASAP7_75t_L g2544 ( 
.A(n_2113),
.Y(n_2544)
);

OAI21x1_ASAP7_75t_L g2545 ( 
.A1(n_2096),
.A2(n_2026),
.B(n_1976),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2126),
.B(n_2062),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2135),
.Y(n_2547)
);

OAI22x1_ASAP7_75t_SL g2548 ( 
.A1(n_2110),
.A2(n_1818),
.B1(n_1820),
.B2(n_1811),
.Y(n_2548)
);

INVx3_ASAP7_75t_L g2549 ( 
.A(n_2113),
.Y(n_2549)
);

OAI22xp5_ASAP7_75t_SL g2550 ( 
.A1(n_2210),
.A2(n_1835),
.B1(n_1837),
.B2(n_1831),
.Y(n_2550)
);

BUFx12f_ASAP7_75t_L g2551 ( 
.A(n_2098),
.Y(n_2551)
);

BUFx8_ASAP7_75t_SL g2552 ( 
.A(n_2098),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2126),
.B(n_1354),
.Y(n_2553)
);

INVx3_ASAP7_75t_L g2554 ( 
.A(n_2113),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2135),
.Y(n_2555)
);

BUFx2_ASAP7_75t_L g2556 ( 
.A(n_2108),
.Y(n_2556)
);

INVxp67_ASAP7_75t_L g2557 ( 
.A(n_2116),
.Y(n_2557)
);

AND2x2_ASAP7_75t_SL g2558 ( 
.A(n_2141),
.B(n_1388),
.Y(n_2558)
);

INVx2_ASAP7_75t_SL g2559 ( 
.A(n_2105),
.Y(n_2559)
);

CKINVDCx20_ASAP7_75t_R g2560 ( 
.A(n_2103),
.Y(n_2560)
);

BUFx6f_ASAP7_75t_L g2561 ( 
.A(n_2135),
.Y(n_2561)
);

CKINVDCx5p33_ASAP7_75t_R g2562 ( 
.A(n_2126),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2153),
.B(n_1365),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2135),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2135),
.Y(n_2565)
);

AND2x4_ASAP7_75t_L g2566 ( 
.A(n_2190),
.B(n_1650),
.Y(n_2566)
);

BUFx12f_ASAP7_75t_L g2567 ( 
.A(n_2098),
.Y(n_2567)
);

BUFx6f_ASAP7_75t_L g2568 ( 
.A(n_2135),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_2126),
.Y(n_2569)
);

INVx4_ASAP7_75t_L g2570 ( 
.A(n_2126),
.Y(n_2570)
);

AND2x2_ASAP7_75t_L g2571 ( 
.A(n_2108),
.B(n_1654),
.Y(n_2571)
);

BUFx12f_ASAP7_75t_L g2572 ( 
.A(n_2098),
.Y(n_2572)
);

OAI22x1_ASAP7_75t_R g2573 ( 
.A1(n_2103),
.A2(n_1906),
.B1(n_1920),
.B2(n_1866),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2126),
.B(n_1368),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2135),
.Y(n_2575)
);

BUFx6f_ASAP7_75t_L g2576 ( 
.A(n_2135),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2135),
.Y(n_2577)
);

BUFx2_ASAP7_75t_L g2578 ( 
.A(n_2108),
.Y(n_2578)
);

AOI22x1_ASAP7_75t_SL g2579 ( 
.A1(n_2103),
.A2(n_1930),
.B1(n_1966),
.B2(n_1927),
.Y(n_2579)
);

BUFx6f_ASAP7_75t_L g2580 ( 
.A(n_2135),
.Y(n_2580)
);

CKINVDCx5p33_ASAP7_75t_R g2581 ( 
.A(n_2126),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2126),
.B(n_1373),
.Y(n_2582)
);

BUFx8_ASAP7_75t_SL g2583 ( 
.A(n_2098),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2135),
.Y(n_2584)
);

INVx2_ASAP7_75t_SL g2585 ( 
.A(n_2105),
.Y(n_2585)
);

INVx5_ASAP7_75t_L g2586 ( 
.A(n_2191),
.Y(n_2586)
);

BUFx6f_ASAP7_75t_L g2587 ( 
.A(n_2135),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_2333),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2396),
.Y(n_2589)
);

BUFx3_ASAP7_75t_L g2590 ( 
.A(n_2517),
.Y(n_2590)
);

AND3x1_ASAP7_75t_L g2591 ( 
.A(n_2281),
.B(n_1863),
.C(n_1763),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2397),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2485),
.Y(n_2593)
);

INVx3_ASAP7_75t_L g2594 ( 
.A(n_2285),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2405),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2562),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2282),
.Y(n_2597)
);

INVx4_ASAP7_75t_L g2598 ( 
.A(n_2302),
.Y(n_2598)
);

BUFx2_ASAP7_75t_L g2599 ( 
.A(n_2335),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2290),
.Y(n_2600)
);

NAND2x1p5_ASAP7_75t_L g2601 ( 
.A(n_2480),
.B(n_1394),
.Y(n_2601)
);

CKINVDCx5p33_ASAP7_75t_R g2602 ( 
.A(n_2569),
.Y(n_2602)
);

BUFx8_ASAP7_75t_L g2603 ( 
.A(n_2506),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2408),
.Y(n_2604)
);

NAND2xp33_ASAP7_75t_L g2605 ( 
.A(n_2456),
.B(n_1581),
.Y(n_2605)
);

AND2x4_ASAP7_75t_L g2606 ( 
.A(n_2261),
.B(n_2043),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2267),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2391),
.Y(n_2608)
);

OA21x2_ASAP7_75t_L g2609 ( 
.A1(n_2337),
.A2(n_1412),
.B(n_1404),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2432),
.Y(n_2610)
);

INVx3_ASAP7_75t_L g2611 ( 
.A(n_2286),
.Y(n_2611)
);

INVx4_ASAP7_75t_L g2612 ( 
.A(n_2581),
.Y(n_2612)
);

INVx4_ASAP7_75t_L g2613 ( 
.A(n_2411),
.Y(n_2613)
);

HB1xp67_ASAP7_75t_L g2614 ( 
.A(n_2435),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2407),
.B(n_1420),
.Y(n_2615)
);

BUFx6f_ASAP7_75t_L g2616 ( 
.A(n_2299),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2439),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2395),
.Y(n_2618)
);

INVx4_ASAP7_75t_L g2619 ( 
.A(n_2260),
.Y(n_2619)
);

CKINVDCx20_ASAP7_75t_R g2620 ( 
.A(n_2560),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2413),
.B(n_2366),
.Y(n_2621)
);

CKINVDCx20_ASAP7_75t_R g2622 ( 
.A(n_2309),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2341),
.B(n_2386),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_SL g2624 ( 
.A(n_2301),
.B(n_1423),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_2477),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2402),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2443),
.Y(n_2627)
);

INVx3_ASAP7_75t_L g2628 ( 
.A(n_2422),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2368),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2416),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2367),
.B(n_1435),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2424),
.Y(n_2632)
);

INVx3_ASAP7_75t_L g2633 ( 
.A(n_2445),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2389),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2399),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2400),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2451),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2412),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2271),
.Y(n_2639)
);

BUFx6f_ASAP7_75t_L g2640 ( 
.A(n_2452),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2417),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2455),
.Y(n_2642)
);

CKINVDCx5p33_ASAP7_75t_R g2643 ( 
.A(n_2430),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2421),
.Y(n_2644)
);

INVx3_ASAP7_75t_L g2645 ( 
.A(n_2457),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_2453),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_2552),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_L g2648 ( 
.A(n_2459),
.Y(n_2648)
);

BUFx6f_ASAP7_75t_L g2649 ( 
.A(n_2460),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2472),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2583),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_2390),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2264),
.Y(n_2653)
);

CKINVDCx20_ASAP7_75t_R g2654 ( 
.A(n_2427),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2473),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_2537),
.Y(n_2656)
);

BUFx2_ASAP7_75t_L g2657 ( 
.A(n_2492),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_2543),
.Y(n_2658)
);

CKINVDCx20_ASAP7_75t_R g2659 ( 
.A(n_2518),
.Y(n_2659)
);

CKINVDCx20_ASAP7_75t_R g2660 ( 
.A(n_2521),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2297),
.Y(n_2661)
);

CKINVDCx5p33_ASAP7_75t_R g2662 ( 
.A(n_2551),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2312),
.Y(n_2663)
);

AND2x6_ASAP7_75t_L g2664 ( 
.A(n_2308),
.B(n_1581),
.Y(n_2664)
);

BUFx6f_ASAP7_75t_L g2665 ( 
.A(n_2474),
.Y(n_2665)
);

CKINVDCx5p33_ASAP7_75t_R g2666 ( 
.A(n_2567),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2434),
.B(n_1444),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2497),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2319),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2324),
.Y(n_2670)
);

CKINVDCx5p33_ASAP7_75t_R g2671 ( 
.A(n_2572),
.Y(n_2671)
);

CKINVDCx5p33_ASAP7_75t_R g2672 ( 
.A(n_2463),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2498),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2388),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2500),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2501),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2419),
.Y(n_2677)
);

CKINVDCx20_ASAP7_75t_R g2678 ( 
.A(n_2268),
.Y(n_2678)
);

CKINVDCx16_ASAP7_75t_R g2679 ( 
.A(n_2274),
.Y(n_2679)
);

AND2x4_ASAP7_75t_L g2680 ( 
.A(n_2495),
.B(n_1306),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2418),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2289),
.B(n_2320),
.Y(n_2682)
);

CKINVDCx5p33_ASAP7_75t_R g2683 ( 
.A(n_2570),
.Y(n_2683)
);

CKINVDCx5p33_ASAP7_75t_R g2684 ( 
.A(n_2493),
.Y(n_2684)
);

CKINVDCx5p33_ASAP7_75t_R g2685 ( 
.A(n_2505),
.Y(n_2685)
);

CKINVDCx20_ASAP7_75t_R g2686 ( 
.A(n_2294),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2420),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2502),
.Y(n_2688)
);

CKINVDCx5p33_ASAP7_75t_R g2689 ( 
.A(n_2556),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2276),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2270),
.B(n_1439),
.Y(n_2691)
);

BUFx6f_ASAP7_75t_L g2692 ( 
.A(n_2512),
.Y(n_2692)
);

AND2x4_ASAP7_75t_L g2693 ( 
.A(n_2504),
.B(n_1309),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2295),
.Y(n_2694)
);

NOR2x1_ASAP7_75t_L g2695 ( 
.A(n_2263),
.B(n_1317),
.Y(n_2695)
);

HB1xp67_ASAP7_75t_L g2696 ( 
.A(n_2511),
.Y(n_2696)
);

BUFx6f_ASAP7_75t_L g2697 ( 
.A(n_2516),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2544),
.Y(n_2698)
);

INVx3_ASAP7_75t_L g2699 ( 
.A(n_2520),
.Y(n_2699)
);

CKINVDCx20_ASAP7_75t_R g2700 ( 
.A(n_2449),
.Y(n_2700)
);

INVx3_ASAP7_75t_L g2701 ( 
.A(n_2524),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2549),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2527),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2448),
.B(n_1447),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2554),
.Y(n_2705)
);

AND2x4_ASAP7_75t_L g2706 ( 
.A(n_2454),
.B(n_1322),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2414),
.Y(n_2707)
);

CKINVDCx5p33_ASAP7_75t_R g2708 ( 
.A(n_2578),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2342),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2490),
.B(n_1459),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_2563),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2546),
.B(n_1465),
.Y(n_2712)
);

OAI21x1_ASAP7_75t_L g2713 ( 
.A1(n_2415),
.A2(n_1429),
.B(n_1428),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_2332),
.Y(n_2714)
);

BUFx6f_ASAP7_75t_L g2715 ( 
.A(n_2536),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_2530),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2278),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_2329),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2279),
.Y(n_2719)
);

CKINVDCx5p33_ASAP7_75t_R g2720 ( 
.A(n_2392),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2283),
.Y(n_2721)
);

HB1xp67_ASAP7_75t_L g2722 ( 
.A(n_2438),
.Y(n_2722)
);

INVxp67_ASAP7_75t_L g2723 ( 
.A(n_2349),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2288),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2292),
.Y(n_2725)
);

BUFx3_ASAP7_75t_L g2726 ( 
.A(n_2539),
.Y(n_2726)
);

INVxp67_ASAP7_75t_L g2727 ( 
.A(n_2350),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2304),
.Y(n_2728)
);

INVx3_ASAP7_75t_L g2729 ( 
.A(n_2561),
.Y(n_2729)
);

CKINVDCx20_ASAP7_75t_R g2730 ( 
.A(n_2298),
.Y(n_2730)
);

CKINVDCx20_ASAP7_75t_R g2731 ( 
.A(n_2458),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2568),
.Y(n_2732)
);

AND2x6_ASAP7_75t_L g2733 ( 
.A(n_2426),
.B(n_1581),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2305),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2325),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2436),
.B(n_1476),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2576),
.Y(n_2737)
);

OA21x2_ASAP7_75t_L g2738 ( 
.A1(n_2440),
.A2(n_1499),
.B(n_1478),
.Y(n_2738)
);

INVx3_ASAP7_75t_L g2739 ( 
.A(n_2580),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2553),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2327),
.Y(n_2741)
);

HB1xp67_ASAP7_75t_L g2742 ( 
.A(n_2479),
.Y(n_2742)
);

CKINVDCx20_ASAP7_75t_R g2743 ( 
.A(n_2507),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_2574),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2587),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2336),
.Y(n_2746)
);

BUFx6f_ASAP7_75t_L g2747 ( 
.A(n_2300),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2429),
.Y(n_2748)
);

BUFx6f_ASAP7_75t_L g2749 ( 
.A(n_2315),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2437),
.B(n_2526),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2317),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2442),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_2582),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2280),
.B(n_1513),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2296),
.B(n_1522),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2340),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_SL g2757 ( 
.A(n_2525),
.B(n_1525),
.Y(n_2757)
);

AND2x4_ASAP7_75t_L g2758 ( 
.A(n_2559),
.B(n_1323),
.Y(n_2758)
);

INVxp67_ASAP7_75t_SL g2759 ( 
.A(n_2330),
.Y(n_2759)
);

INVx3_ASAP7_75t_L g2760 ( 
.A(n_2338),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2343),
.Y(n_2761)
);

CKINVDCx5p33_ASAP7_75t_R g2762 ( 
.A(n_2322),
.Y(n_2762)
);

CKINVDCx20_ASAP7_75t_R g2763 ( 
.A(n_2313),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2348),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2351),
.Y(n_2765)
);

NOR2xp33_ASAP7_75t_R g2766 ( 
.A(n_2585),
.B(n_1527),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2356),
.Y(n_2767)
);

INVx3_ASAP7_75t_L g2768 ( 
.A(n_2345),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_2346),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2450),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2461),
.Y(n_2771)
);

CKINVDCx20_ASAP7_75t_R g2772 ( 
.A(n_2425),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2444),
.B(n_1439),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2359),
.Y(n_2774)
);

INVxp33_ASAP7_75t_L g2775 ( 
.A(n_2573),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_2306),
.Y(n_2776)
);

CKINVDCx5p33_ASAP7_75t_R g2777 ( 
.A(n_2307),
.Y(n_2777)
);

BUFx2_ASAP7_75t_L g2778 ( 
.A(n_2334),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2361),
.Y(n_2779)
);

HB1xp67_ASAP7_75t_L g2780 ( 
.A(n_2311),
.Y(n_2780)
);

HB1xp67_ASAP7_75t_L g2781 ( 
.A(n_2541),
.Y(n_2781)
);

INVx3_ASAP7_75t_L g2782 ( 
.A(n_2357),
.Y(n_2782)
);

NOR2xp33_ASAP7_75t_R g2783 ( 
.A(n_2384),
.B(n_1531),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2481),
.Y(n_2784)
);

INVx2_ASAP7_75t_SL g2785 ( 
.A(n_2542),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2362),
.Y(n_2786)
);

CKINVDCx5p33_ASAP7_75t_R g2787 ( 
.A(n_2318),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2374),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2484),
.Y(n_2789)
);

NOR2xp33_ASAP7_75t_L g2790 ( 
.A(n_2323),
.B(n_1356),
.Y(n_2790)
);

INVx3_ASAP7_75t_L g2791 ( 
.A(n_2365),
.Y(n_2791)
);

CKINVDCx5p33_ASAP7_75t_R g2792 ( 
.A(n_2510),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2486),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2571),
.B(n_1506),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_SL g2795 ( 
.A(n_2558),
.B(n_1554),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2378),
.Y(n_2796)
);

BUFx6f_ASAP7_75t_L g2797 ( 
.A(n_2375),
.Y(n_2797)
);

INVx5_ASAP7_75t_L g2798 ( 
.A(n_2334),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2379),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_L g2800 ( 
.A(n_2376),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2275),
.B(n_1357),
.Y(n_2801)
);

HB1xp67_ASAP7_75t_L g2802 ( 
.A(n_2557),
.Y(n_2802)
);

CKINVDCx5p33_ASAP7_75t_R g2803 ( 
.A(n_2347),
.Y(n_2803)
);

CKINVDCx20_ASAP7_75t_R g2804 ( 
.A(n_2550),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_2464),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2385),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2352),
.Y(n_2807)
);

INVx4_ASAP7_75t_L g2808 ( 
.A(n_2393),
.Y(n_2808)
);

BUFx6f_ASAP7_75t_L g2809 ( 
.A(n_2381),
.Y(n_2809)
);

HB1xp67_ASAP7_75t_L g2810 ( 
.A(n_2371),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2488),
.Y(n_2811)
);

CKINVDCx5p33_ASAP7_75t_R g2812 ( 
.A(n_2579),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2509),
.Y(n_2813)
);

CKINVDCx5p33_ASAP7_75t_R g2814 ( 
.A(n_2456),
.Y(n_2814)
);

BUFx2_ASAP7_75t_L g2815 ( 
.A(n_2409),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2321),
.B(n_1506),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2514),
.Y(n_2817)
);

CKINVDCx5p33_ASAP7_75t_R g2818 ( 
.A(n_2383),
.Y(n_2818)
);

INVx3_ASAP7_75t_L g2819 ( 
.A(n_2291),
.Y(n_2819)
);

CKINVDCx5p33_ASAP7_75t_R g2820 ( 
.A(n_2476),
.Y(n_2820)
);

BUFx3_ASAP7_75t_L g2821 ( 
.A(n_2398),
.Y(n_2821)
);

CKINVDCx5p33_ASAP7_75t_R g2822 ( 
.A(n_2528),
.Y(n_2822)
);

CKINVDCx20_ASAP7_75t_R g2823 ( 
.A(n_2303),
.Y(n_2823)
);

BUFx2_ASAP7_75t_L g2824 ( 
.A(n_2409),
.Y(n_2824)
);

XOR2xp5_ASAP7_75t_L g2825 ( 
.A(n_2273),
.B(n_1558),
.Y(n_2825)
);

INVx3_ASAP7_75t_L g2826 ( 
.A(n_2291),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2531),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2532),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2538),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2555),
.Y(n_2830)
);

INVx4_ASAP7_75t_L g2831 ( 
.A(n_2394),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2565),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2586),
.B(n_1615),
.Y(n_2833)
);

CKINVDCx5p33_ASAP7_75t_R g2834 ( 
.A(n_2406),
.Y(n_2834)
);

CKINVDCx5p33_ASAP7_75t_R g2835 ( 
.A(n_2277),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2447),
.B(n_1615),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2575),
.Y(n_2837)
);

HB1xp67_ASAP7_75t_L g2838 ( 
.A(n_2401),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2577),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2529),
.Y(n_2840)
);

CKINVDCx5p33_ASAP7_75t_R g2841 ( 
.A(n_2503),
.Y(n_2841)
);

CKINVDCx5p33_ASAP7_75t_R g2842 ( 
.A(n_2508),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2545),
.Y(n_2843)
);

OAI21x1_ASAP7_75t_L g2844 ( 
.A1(n_2269),
.A2(n_2314),
.B(n_2284),
.Y(n_2844)
);

CKINVDCx20_ASAP7_75t_R g2845 ( 
.A(n_2466),
.Y(n_2845)
);

CKINVDCx5p33_ASAP7_75t_R g2846 ( 
.A(n_2523),
.Y(n_2846)
);

AND2x4_ASAP7_75t_L g2847 ( 
.A(n_2433),
.B(n_1324),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2310),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2316),
.Y(n_2849)
);

CKINVDCx5p33_ASAP7_75t_R g2850 ( 
.A(n_2534),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2328),
.Y(n_2851)
);

HB1xp67_ASAP7_75t_L g2852 ( 
.A(n_2566),
.Y(n_2852)
);

CKINVDCx5p33_ASAP7_75t_R g2853 ( 
.A(n_2535),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_2540),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2339),
.Y(n_2855)
);

CKINVDCx5p33_ASAP7_75t_R g2856 ( 
.A(n_2410),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2344),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2353),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2354),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2355),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_R g2861 ( 
.A(n_2373),
.B(n_1559),
.Y(n_2861)
);

AND2x2_ASAP7_75t_L g2862 ( 
.A(n_2404),
.B(n_1675),
.Y(n_2862)
);

CKINVDCx5p33_ASAP7_75t_R g2863 ( 
.A(n_2548),
.Y(n_2863)
);

CKINVDCx5p33_ASAP7_75t_R g2864 ( 
.A(n_2403),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2387),
.B(n_1359),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2358),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2360),
.Y(n_2867)
);

BUFx2_ASAP7_75t_L g2868 ( 
.A(n_2462),
.Y(n_2868)
);

CKINVDCx5p33_ASAP7_75t_R g2869 ( 
.A(n_2331),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2364),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2471),
.B(n_1569),
.Y(n_2871)
);

BUFx6f_ASAP7_75t_L g2872 ( 
.A(n_2370),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2515),
.B(n_1572),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2372),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2377),
.Y(n_2875)
);

CKINVDCx5p33_ASAP7_75t_R g2876 ( 
.A(n_2522),
.Y(n_2876)
);

CKINVDCx5p33_ASAP7_75t_R g2877 ( 
.A(n_2533),
.Y(n_2877)
);

NAND2xp33_ASAP7_75t_L g2878 ( 
.A(n_2482),
.B(n_1868),
.Y(n_2878)
);

CKINVDCx20_ASAP7_75t_R g2879 ( 
.A(n_2326),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2380),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2382),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2258),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2259),
.Y(n_2883)
);

CKINVDCx5p33_ASAP7_75t_R g2884 ( 
.A(n_2513),
.Y(n_2884)
);

AND2x2_ASAP7_75t_L g2885 ( 
.A(n_2265),
.B(n_1675),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2423),
.B(n_2363),
.Y(n_2886)
);

CKINVDCx5p33_ASAP7_75t_R g2887 ( 
.A(n_2369),
.Y(n_2887)
);

HB1xp67_ASAP7_75t_L g2888 ( 
.A(n_2287),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2266),
.Y(n_2889)
);

INVxp67_ASAP7_75t_L g2890 ( 
.A(n_2272),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2428),
.Y(n_2891)
);

CKINVDCx5p33_ASAP7_75t_R g2892 ( 
.A(n_2293),
.Y(n_2892)
);

CKINVDCx5p33_ASAP7_75t_R g2893 ( 
.A(n_2446),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2465),
.Y(n_2894)
);

BUFx6f_ASAP7_75t_L g2895 ( 
.A(n_2431),
.Y(n_2895)
);

CKINVDCx5p33_ASAP7_75t_R g2896 ( 
.A(n_2467),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2468),
.Y(n_2897)
);

CKINVDCx5p33_ASAP7_75t_R g2898 ( 
.A(n_2469),
.Y(n_2898)
);

NAND2xp33_ASAP7_75t_SL g2899 ( 
.A(n_2262),
.B(n_1972),
.Y(n_2899)
);

HB1xp67_ASAP7_75t_L g2900 ( 
.A(n_2470),
.Y(n_2900)
);

INVx2_ASAP7_75t_SL g2901 ( 
.A(n_2475),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2748),
.Y(n_2902)
);

INVx2_ASAP7_75t_SL g2903 ( 
.A(n_2599),
.Y(n_2903)
);

INVx1_ASAP7_75t_SL g2904 ( 
.A(n_2838),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2752),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2682),
.B(n_2750),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2900),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2718),
.B(n_2711),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_SL g2909 ( 
.A(n_2776),
.B(n_2777),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2740),
.B(n_2744),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2770),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2771),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_SL g2913 ( 
.A(n_2787),
.B(n_1574),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2784),
.Y(n_2914)
);

INVx2_ASAP7_75t_SL g2915 ( 
.A(n_2621),
.Y(n_2915)
);

BUFx3_ASAP7_75t_L g2916 ( 
.A(n_2590),
.Y(n_2916)
);

BUFx3_ASAP7_75t_L g2917 ( 
.A(n_2620),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_SL g2918 ( 
.A(n_2623),
.B(n_1577),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2789),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2753),
.B(n_2441),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_2798),
.B(n_1601),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2677),
.Y(n_2922)
);

CKINVDCx20_ASAP7_75t_R g2923 ( 
.A(n_2622),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2790),
.B(n_1613),
.Y(n_2924)
);

INVx5_ASAP7_75t_L g2925 ( 
.A(n_2747),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_SL g2926 ( 
.A(n_2798),
.B(n_1630),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2717),
.Y(n_2927)
);

INVx3_ASAP7_75t_L g2928 ( 
.A(n_2616),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2719),
.Y(n_2929)
);

AOI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2869),
.A2(n_1632),
.B1(n_1653),
.B2(n_1645),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2721),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2793),
.Y(n_2932)
);

INVx3_ASAP7_75t_L g2933 ( 
.A(n_2616),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2785),
.B(n_1663),
.Y(n_2934)
);

NAND2xp33_ASAP7_75t_SL g2935 ( 
.A(n_2778),
.B(n_1981),
.Y(n_2935)
);

INVxp67_ASAP7_75t_SL g2936 ( 
.A(n_2895),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2724),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_L g2938 ( 
.A(n_2615),
.B(n_1679),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2827),
.Y(n_2939)
);

BUFx4f_ASAP7_75t_L g2940 ( 
.A(n_2601),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2725),
.Y(n_2941)
);

OR2x2_ASAP7_75t_L g2942 ( 
.A(n_2780),
.B(n_1693),
.Y(n_2942)
);

OAI22xp5_ASAP7_75t_L g2943 ( 
.A1(n_2736),
.A2(n_1684),
.B1(n_1690),
.B2(n_1664),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2728),
.Y(n_2944)
);

AOI22xp33_ASAP7_75t_L g2945 ( 
.A1(n_2895),
.A2(n_2886),
.B1(n_2801),
.B2(n_2862),
.Y(n_2945)
);

INVxp67_ASAP7_75t_SL g2946 ( 
.A(n_2872),
.Y(n_2946)
);

INVx2_ASAP7_75t_SL g2947 ( 
.A(n_2885),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2734),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2735),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2741),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_SL g2951 ( 
.A(n_2613),
.B(n_1700),
.Y(n_2951)
);

INVxp67_ASAP7_75t_SL g2952 ( 
.A(n_2872),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2672),
.B(n_1713),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2829),
.Y(n_2954)
);

INVx3_ASAP7_75t_L g2955 ( 
.A(n_2640),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2631),
.B(n_1717),
.Y(n_2956)
);

AND2x2_ASAP7_75t_SL g2957 ( 
.A(n_2679),
.B(n_1481),
.Y(n_2957)
);

AND2x2_ASAP7_75t_SL g2958 ( 
.A(n_2815),
.B(n_1489),
.Y(n_2958)
);

NAND2xp33_ASAP7_75t_L g2959 ( 
.A(n_2695),
.B(n_1720),
.Y(n_2959)
);

BUFx6f_ASAP7_75t_L g2960 ( 
.A(n_2640),
.Y(n_2960)
);

NAND2xp33_ASAP7_75t_L g2961 ( 
.A(n_2664),
.B(n_2783),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2832),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2644),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2851),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_SL g2965 ( 
.A(n_2683),
.B(n_1724),
.Y(n_2965)
);

INVx1_ASAP7_75t_SL g2966 ( 
.A(n_2731),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2859),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2746),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2870),
.Y(n_2969)
);

OR2x6_ASAP7_75t_L g2970 ( 
.A(n_2598),
.B(n_1336),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2894),
.Y(n_2971)
);

INVx3_ASAP7_75t_L g2972 ( 
.A(n_2648),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2756),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2761),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_SL g2975 ( 
.A(n_2861),
.B(n_2864),
.Y(n_2975)
);

HB1xp67_ASAP7_75t_L g2976 ( 
.A(n_2722),
.Y(n_2976)
);

INVx3_ASAP7_75t_L g2977 ( 
.A(n_2648),
.Y(n_2977)
);

NAND3xp33_ASAP7_75t_L g2978 ( 
.A(n_2605),
.B(n_1364),
.C(n_1361),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2764),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_SL g2980 ( 
.A(n_2816),
.B(n_1729),
.Y(n_2980)
);

AND2x2_ASAP7_75t_SL g2981 ( 
.A(n_2824),
.B(n_2591),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_L g2982 ( 
.A(n_2723),
.B(n_1766),
.Y(n_2982)
);

AOI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2856),
.A2(n_2834),
.B1(n_2854),
.B2(n_2822),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_SL g2984 ( 
.A(n_2781),
.B(n_1733),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2634),
.Y(n_2985)
);

INVx4_ASAP7_75t_L g2986 ( 
.A(n_2747),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2635),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_SL g2988 ( 
.A(n_2773),
.B(n_1742),
.Y(n_2988)
);

NOR2xp33_ASAP7_75t_L g2989 ( 
.A(n_2727),
.B(n_1822),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2636),
.Y(n_2990)
);

AND2x6_ASAP7_75t_L g2991 ( 
.A(n_2840),
.B(n_1868),
.Y(n_2991)
);

INVx4_ASAP7_75t_L g2992 ( 
.A(n_2749),
.Y(n_2992)
);

AOI22xp33_ASAP7_75t_L g2993 ( 
.A1(n_2608),
.A2(n_1293),
.B1(n_1548),
.B2(n_1540),
.Y(n_2993)
);

INVx3_ASAP7_75t_L g2994 ( 
.A(n_2649),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2704),
.B(n_1748),
.Y(n_2995)
);

INVx3_ASAP7_75t_L g2996 ( 
.A(n_2649),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2765),
.Y(n_2997)
);

OR2x6_ASAP7_75t_L g2998 ( 
.A(n_2657),
.B(n_1355),
.Y(n_2998)
);

XNOR2xp5_ASAP7_75t_L g2999 ( 
.A(n_2654),
.B(n_1983),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2767),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2638),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2774),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2641),
.Y(n_3003)
);

INVx3_ASAP7_75t_L g3004 ( 
.A(n_2665),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2794),
.B(n_1749),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2779),
.Y(n_3006)
);

BUFx10_ASAP7_75t_L g3007 ( 
.A(n_2639),
.Y(n_3007)
);

INVx3_ASAP7_75t_L g3008 ( 
.A(n_2665),
.Y(n_3008)
);

INVxp67_ASAP7_75t_SL g3009 ( 
.A(n_2890),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2811),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2710),
.B(n_1833),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_SL g3012 ( 
.A(n_2712),
.B(n_1751),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_SL g3013 ( 
.A(n_2865),
.B(n_1757),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_2802),
.B(n_2667),
.Y(n_3014)
);

INVxp33_ASAP7_75t_L g3015 ( 
.A(n_2742),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2786),
.Y(n_3016)
);

BUFx10_ASAP7_75t_L g3017 ( 
.A(n_2643),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2813),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2754),
.B(n_1855),
.Y(n_3019)
);

OR2x6_ASAP7_75t_L g3020 ( 
.A(n_2612),
.B(n_1358),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_SL g3021 ( 
.A(n_2808),
.B(n_1769),
.Y(n_3021)
);

BUFx6f_ASAP7_75t_L g3022 ( 
.A(n_2692),
.Y(n_3022)
);

HB1xp67_ASAP7_75t_L g3023 ( 
.A(n_2852),
.Y(n_3023)
);

BUFx3_ASAP7_75t_L g3024 ( 
.A(n_2726),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2618),
.B(n_1772),
.Y(n_3025)
);

BUFx10_ASAP7_75t_L g3026 ( 
.A(n_2646),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2626),
.B(n_1779),
.Y(n_3027)
);

INVx3_ASAP7_75t_L g3028 ( 
.A(n_2692),
.Y(n_3028)
);

BUFx6f_ASAP7_75t_SL g3029 ( 
.A(n_2680),
.Y(n_3029)
);

BUFx10_ASAP7_75t_L g3030 ( 
.A(n_2647),
.Y(n_3030)
);

OR2x6_ASAP7_75t_L g3031 ( 
.A(n_2868),
.B(n_1376),
.Y(n_3031)
);

OR2x2_ASAP7_75t_L g3032 ( 
.A(n_2807),
.B(n_1900),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2788),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2796),
.Y(n_3034)
);

BUFx4f_ASAP7_75t_L g3035 ( 
.A(n_2664),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2799),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_SL g3037 ( 
.A(n_2831),
.B(n_2893),
.Y(n_3037)
);

INVx5_ASAP7_75t_L g3038 ( 
.A(n_2749),
.Y(n_3038)
);

AOI22xp33_ASAP7_75t_L g3039 ( 
.A1(n_2630),
.A2(n_1293),
.B1(n_1592),
.B2(n_1550),
.Y(n_3039)
);

INVxp67_ASAP7_75t_SL g3040 ( 
.A(n_2897),
.Y(n_3040)
);

BUFx6f_ASAP7_75t_L g3041 ( 
.A(n_2697),
.Y(n_3041)
);

AND2x6_ASAP7_75t_L g3042 ( 
.A(n_2843),
.B(n_1868),
.Y(n_3042)
);

AND2x6_ASAP7_75t_L g3043 ( 
.A(n_2691),
.B(n_1377),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_SL g3044 ( 
.A(n_2896),
.B(n_1790),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2806),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2817),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2828),
.Y(n_3047)
);

BUFx10_ASAP7_75t_L g3048 ( 
.A(n_2651),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2830),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2837),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_2632),
.A2(n_1696),
.B1(n_1722),
.B2(n_1652),
.Y(n_3051)
);

INVx3_ASAP7_75t_L g3052 ( 
.A(n_2697),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2839),
.Y(n_3053)
);

BUFx10_ASAP7_75t_L g3054 ( 
.A(n_2588),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2681),
.Y(n_3055)
);

NOR2xp33_ASAP7_75t_L g3056 ( 
.A(n_2755),
.B(n_1919),
.Y(n_3056)
);

BUFx3_ASAP7_75t_L g3057 ( 
.A(n_2797),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2687),
.Y(n_3058)
);

AND2x4_ASAP7_75t_L g3059 ( 
.A(n_2633),
.B(n_2478),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2882),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2733),
.B(n_1792),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2883),
.Y(n_3062)
);

AOI22xp33_ASAP7_75t_L g3063 ( 
.A1(n_2847),
.A2(n_1838),
.B1(n_1854),
.B2(n_1768),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2889),
.Y(n_3064)
);

AOI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_2887),
.A2(n_1929),
.B1(n_1964),
.B2(n_1871),
.Y(n_3065)
);

INVx3_ASAP7_75t_L g3066 ( 
.A(n_2715),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2733),
.B(n_1799),
.Y(n_3067)
);

INVx3_ASAP7_75t_L g3068 ( 
.A(n_2715),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2891),
.Y(n_3069)
);

AO21x2_ASAP7_75t_L g3070 ( 
.A1(n_2844),
.A2(n_1386),
.B(n_1383),
.Y(n_3070)
);

BUFx3_ASAP7_75t_L g3071 ( 
.A(n_2797),
.Y(n_3071)
);

INVx3_ASAP7_75t_L g3072 ( 
.A(n_2800),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2848),
.Y(n_3073)
);

INVx2_ASAP7_75t_SL g3074 ( 
.A(n_2706),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2898),
.B(n_2876),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2849),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2855),
.Y(n_3077)
);

NOR2xp33_ASAP7_75t_L g3078 ( 
.A(n_2757),
.B(n_1973),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2733),
.B(n_1800),
.Y(n_3079)
);

AOI22xp5_ASAP7_75t_L g3080 ( 
.A1(n_2820),
.A2(n_1807),
.B1(n_1815),
.B2(n_1806),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2857),
.Y(n_3081)
);

AOI22xp33_ASAP7_75t_L g3082 ( 
.A1(n_2879),
.A2(n_2034),
.B1(n_2080),
.B2(n_2006),
.Y(n_3082)
);

XOR2x2_ASAP7_75t_L g3083 ( 
.A(n_2825),
.B(n_1),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2709),
.B(n_1816),
.Y(n_3084)
);

AOI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_2795),
.A2(n_1859),
.B1(n_1881),
.B2(n_1853),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2664),
.B(n_1882),
.Y(n_3086)
);

AOI22xp5_ASAP7_75t_L g3087 ( 
.A1(n_2899),
.A2(n_1893),
.B1(n_1905),
.B2(n_1890),
.Y(n_3087)
);

AOI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_2884),
.A2(n_1950),
.B1(n_1957),
.B2(n_1912),
.Y(n_3088)
);

INVx4_ASAP7_75t_L g3089 ( 
.A(n_2800),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2858),
.Y(n_3090)
);

OA22x2_ASAP7_75t_L g3091 ( 
.A1(n_2814),
.A2(n_1371),
.B1(n_1372),
.B2(n_1366),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2860),
.Y(n_3092)
);

BUFx4f_ASAP7_75t_L g3093 ( 
.A(n_2606),
.Y(n_3093)
);

INVx2_ASAP7_75t_SL g3094 ( 
.A(n_2758),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2866),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2867),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2874),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_2810),
.B(n_1375),
.Y(n_3098)
);

CKINVDCx5p33_ASAP7_75t_R g3099 ( 
.A(n_2593),
.Y(n_3099)
);

NOR2xp33_ASAP7_75t_L g3100 ( 
.A(n_2818),
.B(n_1379),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2875),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2597),
.B(n_2600),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2880),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2881),
.Y(n_3104)
);

AOI22xp5_ASAP7_75t_L g3105 ( 
.A1(n_2624),
.A2(n_1974),
.B1(n_1982),
.B2(n_1969),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_SL g3106 ( 
.A(n_2877),
.B(n_1985),
.Y(n_3106)
);

BUFx6f_ASAP7_75t_L g3107 ( 
.A(n_2809),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_2901),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_SL g3109 ( 
.A(n_2619),
.B(n_1988),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2690),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_SL g3111 ( 
.A(n_2766),
.B(n_1996),
.Y(n_3111)
);

INVx1_ASAP7_75t_SL g3112 ( 
.A(n_2743),
.Y(n_3112)
);

NOR2x1p5_ASAP7_75t_L g3113 ( 
.A(n_2714),
.B(n_1380),
.Y(n_3113)
);

BUFx3_ASAP7_75t_L g3114 ( 
.A(n_2809),
.Y(n_3114)
);

OR2x2_ASAP7_75t_L g3115 ( 
.A(n_2693),
.B(n_2483),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_SL g3116 ( 
.A(n_2653),
.B(n_2001),
.Y(n_3116)
);

NOR2x1p5_ASAP7_75t_L g3117 ( 
.A(n_2835),
.B(n_1384),
.Y(n_3117)
);

INVx3_ASAP7_75t_L g3118 ( 
.A(n_2594),
.Y(n_3118)
);

INVx2_ASAP7_75t_SL g3119 ( 
.A(n_2614),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2694),
.Y(n_3120)
);

BUFx3_ASAP7_75t_L g3121 ( 
.A(n_2628),
.Y(n_3121)
);

BUFx8_ASAP7_75t_SL g3122 ( 
.A(n_2659),
.Y(n_3122)
);

BUFx2_ASAP7_75t_L g3123 ( 
.A(n_2769),
.Y(n_3123)
);

BUFx10_ASAP7_75t_L g3124 ( 
.A(n_2625),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2698),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2702),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2705),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2713),
.Y(n_3128)
);

AND2x2_ASAP7_75t_L g3129 ( 
.A(n_2833),
.B(n_2487),
.Y(n_3129)
);

INVx2_ASAP7_75t_SL g3130 ( 
.A(n_2696),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2661),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2607),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2663),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2669),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2670),
.B(n_2002),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2738),
.A2(n_1389),
.B1(n_1391),
.B2(n_1390),
.Y(n_3136)
);

BUFx3_ASAP7_75t_L g3137 ( 
.A(n_2751),
.Y(n_3137)
);

INVx1_ASAP7_75t_SL g3138 ( 
.A(n_2720),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2610),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_SL g3140 ( 
.A(n_2674),
.B(n_2024),
.Y(n_3140)
);

INVx3_ASAP7_75t_L g3141 ( 
.A(n_2611),
.Y(n_3141)
);

AOI22xp33_ASAP7_75t_L g3142 ( 
.A1(n_2609),
.A2(n_2707),
.B1(n_1397),
.B2(n_1406),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2906),
.B(n_2871),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2945),
.B(n_2873),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_2982),
.B(n_2596),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2989),
.B(n_2602),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2902),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2922),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_2910),
.B(n_2762),
.Y(n_3149)
);

BUFx3_ASAP7_75t_L g3150 ( 
.A(n_3107),
.Y(n_3150)
);

INVx4_ASAP7_75t_SL g3151 ( 
.A(n_3029),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2905),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_SL g3153 ( 
.A(n_3014),
.B(n_2629),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_3011),
.B(n_2759),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2927),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2929),
.Y(n_3156)
);

AND2x4_ASAP7_75t_L g3157 ( 
.A(n_2925),
.B(n_2617),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2911),
.Y(n_3158)
);

INVx4_ASAP7_75t_L g3159 ( 
.A(n_2925),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2931),
.Y(n_3160)
);

AND2x4_ASAP7_75t_L g3161 ( 
.A(n_3038),
.B(n_2916),
.Y(n_3161)
);

INVxp67_ASAP7_75t_L g3162 ( 
.A(n_3032),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2937),
.Y(n_3163)
);

BUFx6f_ASAP7_75t_L g3164 ( 
.A(n_3107),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2912),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2914),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_SL g3167 ( 
.A(n_2938),
.B(n_2684),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2941),
.Y(n_3168)
);

AND2x2_ASAP7_75t_L g3169 ( 
.A(n_2903),
.B(n_2836),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_2919),
.Y(n_3170)
);

AOI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_3078),
.A2(n_2804),
.B1(n_2730),
.B2(n_2775),
.Y(n_3171)
);

AND2x2_ASAP7_75t_L g3172 ( 
.A(n_2904),
.B(n_2716),
.Y(n_3172)
);

OR2x2_ASAP7_75t_L g3173 ( 
.A(n_2942),
.B(n_2966),
.Y(n_3173)
);

AND2x4_ASAP7_75t_L g3174 ( 
.A(n_3038),
.B(n_3024),
.Y(n_3174)
);

OAI22xp5_ASAP7_75t_L g3175 ( 
.A1(n_2936),
.A2(n_2845),
.B1(n_2689),
.B2(n_2708),
.Y(n_3175)
);

NOR2xp33_ASAP7_75t_L g3176 ( 
.A(n_2908),
.B(n_2823),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_3100),
.B(n_2685),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_L g3178 ( 
.A(n_2909),
.B(n_2678),
.Y(n_3178)
);

BUFx3_ASAP7_75t_L g3179 ( 
.A(n_2960),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_3019),
.B(n_2627),
.Y(n_3180)
);

BUFx3_ASAP7_75t_L g3181 ( 
.A(n_2960),
.Y(n_3181)
);

AND2x2_ASAP7_75t_L g3182 ( 
.A(n_3056),
.B(n_2637),
.Y(n_3182)
);

AND2x4_ASAP7_75t_L g3183 ( 
.A(n_3121),
.B(n_2642),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2944),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2932),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2939),
.Y(n_3186)
);

AND2x4_ASAP7_75t_L g3187 ( 
.A(n_3137),
.B(n_2650),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2948),
.Y(n_3188)
);

AND2x2_ASAP7_75t_L g3189 ( 
.A(n_2947),
.B(n_2655),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2954),
.Y(n_3190)
);

AO22x2_ASAP7_75t_L g3191 ( 
.A1(n_3112),
.A2(n_2772),
.B1(n_2763),
.B2(n_2792),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2949),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2950),
.Y(n_3193)
);

INVx4_ASAP7_75t_SL g3194 ( 
.A(n_3043),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2968),
.Y(n_3195)
);

BUFx6f_ASAP7_75t_L g3196 ( 
.A(n_3022),
.Y(n_3196)
);

INVxp67_ASAP7_75t_L g3197 ( 
.A(n_2976),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2924),
.B(n_2035),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2973),
.Y(n_3199)
);

OAI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_2920),
.A2(n_2067),
.B1(n_2076),
.B2(n_1997),
.Y(n_3200)
);

NAND2x1p5_ASAP7_75t_L g3201 ( 
.A(n_2986),
.B(n_2645),
.Y(n_3201)
);

CKINVDCx20_ASAP7_75t_R g3202 ( 
.A(n_2923),
.Y(n_3202)
);

INVx3_ASAP7_75t_L g3203 ( 
.A(n_3022),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2962),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3040),
.B(n_2064),
.Y(n_3205)
);

INVxp67_ASAP7_75t_L g3206 ( 
.A(n_3098),
.Y(n_3206)
);

HB1xp67_ASAP7_75t_L g3207 ( 
.A(n_3023),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2915),
.B(n_2668),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2974),
.Y(n_3209)
);

AND2x4_ASAP7_75t_L g3210 ( 
.A(n_3057),
.B(n_2673),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2979),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_3123),
.B(n_2675),
.Y(n_3212)
);

NOR2xp33_ASAP7_75t_L g3213 ( 
.A(n_3015),
.B(n_2958),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_2964),
.Y(n_3214)
);

NOR2xp33_ASAP7_75t_L g3215 ( 
.A(n_2983),
.B(n_2652),
.Y(n_3215)
);

BUFx6f_ASAP7_75t_L g3216 ( 
.A(n_3041),
.Y(n_3216)
);

BUFx6f_ASAP7_75t_L g3217 ( 
.A(n_3041),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_3119),
.B(n_2676),
.Y(n_3218)
);

NAND2x1p5_ASAP7_75t_L g3219 ( 
.A(n_2992),
.B(n_2699),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2995),
.B(n_2065),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2997),
.Y(n_3221)
);

BUFx6f_ASAP7_75t_L g3222 ( 
.A(n_3071),
.Y(n_3222)
);

BUFx6f_ASAP7_75t_L g3223 ( 
.A(n_3114),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_3130),
.B(n_2688),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_SL g3225 ( 
.A(n_2940),
.B(n_2656),
.Y(n_3225)
);

INVx1_ASAP7_75t_SL g3226 ( 
.A(n_3138),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3000),
.Y(n_3227)
);

BUFx2_ASAP7_75t_L g3228 ( 
.A(n_2917),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3002),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3006),
.Y(n_3230)
);

HB1xp67_ASAP7_75t_L g3231 ( 
.A(n_3031),
.Y(n_3231)
);

BUFx6f_ASAP7_75t_L g3232 ( 
.A(n_3089),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3016),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3033),
.Y(n_3234)
);

BUFx3_ASAP7_75t_L g3235 ( 
.A(n_3122),
.Y(n_3235)
);

A2O1A1Ixp33_ASAP7_75t_L g3236 ( 
.A1(n_3034),
.A2(n_2878),
.B(n_1415),
.C(n_1424),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3036),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_2967),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_2907),
.B(n_2703),
.Y(n_3239)
);

INVxp67_ASAP7_75t_L g3240 ( 
.A(n_3115),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_SL g3241 ( 
.A(n_3108),
.B(n_2658),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3045),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_SL g3243 ( 
.A(n_3074),
.B(n_2662),
.Y(n_3243)
);

AOI22xp33_ASAP7_75t_L g3244 ( 
.A1(n_3060),
.A2(n_1430),
.B1(n_1441),
.B2(n_1395),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3064),
.Y(n_3245)
);

INVxp67_ASAP7_75t_L g3246 ( 
.A(n_3094),
.Y(n_3246)
);

CKINVDCx5p33_ASAP7_75t_R g3247 ( 
.A(n_3099),
.Y(n_3247)
);

INVx8_ASAP7_75t_L g3248 ( 
.A(n_3043),
.Y(n_3248)
);

AND2x6_ASAP7_75t_L g3249 ( 
.A(n_3087),
.B(n_2732),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3069),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3046),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3049),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_SL g3253 ( 
.A(n_2930),
.B(n_2666),
.Y(n_3253)
);

NOR2xp33_ASAP7_75t_L g3254 ( 
.A(n_2913),
.B(n_2803),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_L g3255 ( 
.A(n_3009),
.B(n_3080),
.Y(n_3255)
);

AOI22xp5_ASAP7_75t_L g3256 ( 
.A1(n_2956),
.A2(n_2073),
.B1(n_2089),
.B2(n_2068),
.Y(n_3256)
);

INVx3_ASAP7_75t_L g3257 ( 
.A(n_3072),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3050),
.Y(n_3258)
);

AND2x2_ASAP7_75t_L g3259 ( 
.A(n_3129),
.B(n_2737),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_2969),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_2963),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3058),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3076),
.Y(n_3263)
);

AND2x6_ASAP7_75t_L g3264 ( 
.A(n_3131),
.B(n_2745),
.Y(n_3264)
);

INVx3_ASAP7_75t_L g3265 ( 
.A(n_2955),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_3010),
.Y(n_3266)
);

CKINVDCx20_ASAP7_75t_R g3267 ( 
.A(n_3054),
.Y(n_3267)
);

INVx3_ASAP7_75t_L g3268 ( 
.A(n_2972),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_SL g3269 ( 
.A(n_3062),
.B(n_2671),
.Y(n_3269)
);

NOR2xp33_ASAP7_75t_L g3270 ( 
.A(n_3044),
.B(n_2660),
.Y(n_3270)
);

OR2x2_ASAP7_75t_SL g3271 ( 
.A(n_3083),
.B(n_2888),
.Y(n_3271)
);

AND2x4_ASAP7_75t_L g3272 ( 
.A(n_2977),
.B(n_2701),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3077),
.Y(n_3273)
);

INVx4_ASAP7_75t_L g3274 ( 
.A(n_2994),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3081),
.Y(n_3275)
);

INVx4_ASAP7_75t_L g3276 ( 
.A(n_2996),
.Y(n_3276)
);

OR2x6_ASAP7_75t_L g3277 ( 
.A(n_3031),
.B(n_2589),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3082),
.B(n_2592),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3090),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3092),
.Y(n_3280)
);

INVx3_ASAP7_75t_L g3281 ( 
.A(n_3004),
.Y(n_3281)
);

AOI22xp5_ASAP7_75t_L g3282 ( 
.A1(n_3133),
.A2(n_2604),
.B1(n_2595),
.B2(n_2863),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_3075),
.B(n_2729),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3095),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3096),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_2971),
.B(n_2489),
.Y(n_3286)
);

AND2x4_ASAP7_75t_L g3287 ( 
.A(n_3008),
.B(n_2739),
.Y(n_3287)
);

AO22x2_ASAP7_75t_L g3288 ( 
.A1(n_3037),
.A2(n_1446),
.B1(n_1455),
.B2(n_1443),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3018),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_SL g3290 ( 
.A(n_3084),
.B(n_3025),
.Y(n_3290)
);

NOR2xp33_ASAP7_75t_L g3291 ( 
.A(n_2953),
.B(n_2841),
.Y(n_3291)
);

NOR2xp33_ASAP7_75t_L g3292 ( 
.A(n_2965),
.B(n_2842),
.Y(n_3292)
);

AND2x4_ASAP7_75t_L g3293 ( 
.A(n_3028),
.B(n_2760),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3047),
.Y(n_3294)
);

INVx5_ASAP7_75t_L g3295 ( 
.A(n_2970),
.Y(n_3295)
);

NOR2xp33_ASAP7_75t_L g3296 ( 
.A(n_2975),
.B(n_2846),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3097),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_3065),
.B(n_2850),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3104),
.Y(n_3299)
);

NAND2xp33_ASAP7_75t_L g3300 ( 
.A(n_3143),
.B(n_3043),
.Y(n_3300)
);

NOR2xp33_ASAP7_75t_L g3301 ( 
.A(n_3206),
.B(n_2999),
.Y(n_3301)
);

NOR2xp33_ASAP7_75t_L g3302 ( 
.A(n_3145),
.B(n_2935),
.Y(n_3302)
);

OAI22xp5_ASAP7_75t_L g3303 ( 
.A1(n_3255),
.A2(n_3142),
.B1(n_3013),
.B2(n_3136),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3154),
.B(n_2946),
.Y(n_3304)
);

NAND2x1_ASAP7_75t_L g3305 ( 
.A(n_3147),
.B(n_2985),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_3146),
.B(n_2981),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3180),
.B(n_2952),
.Y(n_3307)
);

AOI22xp33_ASAP7_75t_L g3308 ( 
.A1(n_3148),
.A2(n_3091),
.B1(n_2987),
.B2(n_3001),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3155),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_3177),
.B(n_2957),
.Y(n_3310)
);

OAI22xp5_ASAP7_75t_L g3311 ( 
.A1(n_3144),
.A2(n_2918),
.B1(n_3134),
.B2(n_3027),
.Y(n_3311)
);

CKINVDCx5p33_ASAP7_75t_R g3312 ( 
.A(n_3247),
.Y(n_3312)
);

INVx2_ASAP7_75t_SL g3313 ( 
.A(n_3164),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_SL g3314 ( 
.A(n_3172),
.B(n_3035),
.Y(n_3314)
);

AND2x4_ASAP7_75t_L g3315 ( 
.A(n_3161),
.B(n_3052),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3156),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3160),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3163),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3168),
.Y(n_3319)
);

INVxp67_ASAP7_75t_L g3320 ( 
.A(n_3207),
.Y(n_3320)
);

AND2x4_ASAP7_75t_L g3321 ( 
.A(n_3174),
.B(n_3066),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3182),
.B(n_3053),
.Y(n_3322)
);

NAND2xp33_ASAP7_75t_L g3323 ( 
.A(n_3248),
.B(n_2991),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_3162),
.B(n_3093),
.Y(n_3324)
);

A2O1A1Ixp33_ASAP7_75t_L g3325 ( 
.A1(n_3290),
.A2(n_3126),
.B(n_3127),
.C(n_3125),
.Y(n_3325)
);

AOI22xp33_ASAP7_75t_L g3326 ( 
.A1(n_3184),
.A2(n_3003),
.B1(n_3055),
.B2(n_2990),
.Y(n_3326)
);

AOI22xp5_ASAP7_75t_L g3327 ( 
.A1(n_3213),
.A2(n_2943),
.B1(n_2980),
.B2(n_2961),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_SL g3328 ( 
.A(n_3226),
.B(n_3135),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3188),
.B(n_3073),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3152),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3192),
.B(n_3101),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3158),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3193),
.B(n_3103),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_3198),
.A2(n_3128),
.B(n_3012),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_SL g3335 ( 
.A(n_3153),
.B(n_3088),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3195),
.B(n_3110),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_SL g3337 ( 
.A(n_3176),
.B(n_3007),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_SL g3338 ( 
.A(n_3298),
.B(n_3120),
.Y(n_3338)
);

AOI22xp33_ASAP7_75t_L g3339 ( 
.A1(n_3199),
.A2(n_3070),
.B1(n_2978),
.B2(n_3005),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3209),
.Y(n_3340)
);

INVx2_ASAP7_75t_SL g3341 ( 
.A(n_3164),
.Y(n_3341)
);

INVxp67_ASAP7_75t_L g3342 ( 
.A(n_3173),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_3169),
.B(n_3085),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_3165),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3166),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3211),
.B(n_2988),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3221),
.Y(n_3347)
);

INVx2_ASAP7_75t_SL g3348 ( 
.A(n_3196),
.Y(n_3348)
);

AOI22xp33_ASAP7_75t_L g3349 ( 
.A1(n_3227),
.A2(n_2959),
.B1(n_2984),
.B2(n_3102),
.Y(n_3349)
);

NOR2xp33_ASAP7_75t_L g3350 ( 
.A(n_3200),
.B(n_3106),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3229),
.B(n_2951),
.Y(n_3351)
);

INVx4_ASAP7_75t_L g3352 ( 
.A(n_3232),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3170),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3230),
.B(n_3111),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3233),
.B(n_3105),
.Y(n_3355)
);

AOI22xp33_ASAP7_75t_L g3356 ( 
.A1(n_3234),
.A2(n_3140),
.B1(n_3116),
.B2(n_2993),
.Y(n_3356)
);

AND2x4_ASAP7_75t_L g3357 ( 
.A(n_3232),
.B(n_3068),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3237),
.B(n_2934),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3242),
.B(n_3021),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3245),
.B(n_3109),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_L g3361 ( 
.A(n_3167),
.B(n_3197),
.Y(n_3361)
);

BUFx3_ASAP7_75t_L g3362 ( 
.A(n_3150),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3250),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3251),
.B(n_3063),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3252),
.B(n_3132),
.Y(n_3365)
);

BUFx12f_ASAP7_75t_L g3366 ( 
.A(n_3222),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3258),
.B(n_3139),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3262),
.Y(n_3368)
);

OAI22xp5_ASAP7_75t_L g3369 ( 
.A1(n_3220),
.A2(n_3086),
.B1(n_3061),
.B2(n_3079),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3263),
.Y(n_3370)
);

AOI21xp5_ASAP7_75t_L g3371 ( 
.A1(n_3205),
.A2(n_3067),
.B(n_2926),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_3240),
.B(n_2998),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3273),
.B(n_3020),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3275),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_3185),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3279),
.B(n_3020),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3280),
.B(n_3284),
.Y(n_3377)
);

AOI22xp33_ASAP7_75t_L g3378 ( 
.A1(n_3261),
.A2(n_3039),
.B1(n_2998),
.B2(n_2991),
.Y(n_3378)
);

INVxp33_ASAP7_75t_L g3379 ( 
.A(n_3212),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_3285),
.B(n_2921),
.Y(n_3380)
);

NAND3xp33_ASAP7_75t_L g3381 ( 
.A(n_3171),
.B(n_3051),
.C(n_2812),
.Y(n_3381)
);

INVx2_ASAP7_75t_SL g3382 ( 
.A(n_3196),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_SL g3383 ( 
.A(n_3175),
.B(n_3017),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3297),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3299),
.Y(n_3385)
);

NOR2xp33_ASAP7_75t_L g3386 ( 
.A(n_3149),
.B(n_3124),
.Y(n_3386)
);

AOI22xp33_ASAP7_75t_L g3387 ( 
.A1(n_3266),
.A2(n_3042),
.B1(n_2991),
.B2(n_3117),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_3278),
.B(n_3042),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3289),
.B(n_3042),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3294),
.B(n_3059),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3186),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3190),
.B(n_3118),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3204),
.B(n_3141),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3286),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3214),
.B(n_2928),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3238),
.B(n_2933),
.Y(n_3396)
);

OR2x6_ASAP7_75t_L g3397 ( 
.A(n_3248),
.B(n_2970),
.Y(n_3397)
);

OAI22xp5_ASAP7_75t_L g3398 ( 
.A1(n_3260),
.A2(n_3113),
.B1(n_2805),
.B2(n_2853),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3259),
.B(n_3026),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_3239),
.B(n_3030),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_3249),
.A2(n_1467),
.B1(n_1470),
.B2(n_1457),
.Y(n_3401)
);

AOI22xp33_ASAP7_75t_L g3402 ( 
.A1(n_3249),
.A2(n_1480),
.B1(n_1491),
.B2(n_1473),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3208),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_L g3404 ( 
.A(n_3178),
.B(n_3048),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3288),
.B(n_2491),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3256),
.B(n_2494),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3189),
.Y(n_3407)
);

OAI22xp5_ASAP7_75t_L g3408 ( 
.A1(n_3246),
.A2(n_1393),
.B1(n_1400),
.B2(n_1396),
.Y(n_3408)
);

HB1xp67_ASAP7_75t_L g3409 ( 
.A(n_3216),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3264),
.B(n_2496),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_3264),
.B(n_2499),
.Y(n_3411)
);

AND2x4_ASAP7_75t_L g3412 ( 
.A(n_3293),
.B(n_3272),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3264),
.B(n_2519),
.Y(n_3413)
);

AOI22xp33_ASAP7_75t_L g3414 ( 
.A1(n_3249),
.A2(n_1493),
.B1(n_1504),
.B2(n_1492),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3291),
.B(n_2547),
.Y(n_3415)
);

CKINVDCx5p33_ASAP7_75t_R g3416 ( 
.A(n_3202),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_SL g3417 ( 
.A(n_3194),
.B(n_2768),
.Y(n_3417)
);

NOR2xp33_ASAP7_75t_L g3418 ( 
.A(n_3215),
.B(n_2782),
.Y(n_3418)
);

INVx2_ASAP7_75t_SL g3419 ( 
.A(n_3216),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3292),
.B(n_2564),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3218),
.Y(n_3421)
);

AND2x2_ASAP7_75t_L g3422 ( 
.A(n_3224),
.B(n_2791),
.Y(n_3422)
);

INVx3_ASAP7_75t_L g3423 ( 
.A(n_3222),
.Y(n_3423)
);

BUFx6f_ASAP7_75t_L g3424 ( 
.A(n_3217),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3244),
.B(n_2584),
.Y(n_3425)
);

AOI22xp5_ASAP7_75t_L g3426 ( 
.A1(n_3254),
.A2(n_2826),
.B1(n_2819),
.B2(n_1401),
.Y(n_3426)
);

CKINVDCx5p33_ASAP7_75t_R g3427 ( 
.A(n_3235),
.Y(n_3427)
);

INVx2_ASAP7_75t_SL g3428 ( 
.A(n_3217),
.Y(n_3428)
);

OR2x6_ASAP7_75t_L g3429 ( 
.A(n_3159),
.B(n_2821),
.Y(n_3429)
);

INVxp67_ASAP7_75t_SL g3430 ( 
.A(n_3179),
.Y(n_3430)
);

BUFx6f_ASAP7_75t_L g3431 ( 
.A(n_3366),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3309),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3307),
.B(n_3270),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3316),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3394),
.B(n_3296),
.Y(n_3435)
);

BUFx4f_ASAP7_75t_L g3436 ( 
.A(n_3424),
.Y(n_3436)
);

NOR2xp33_ASAP7_75t_R g3437 ( 
.A(n_3416),
.B(n_3267),
.Y(n_3437)
);

INVx3_ASAP7_75t_L g3438 ( 
.A(n_3352),
.Y(n_3438)
);

INVx3_ASAP7_75t_L g3439 ( 
.A(n_3362),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3317),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3318),
.Y(n_3441)
);

BUFx3_ASAP7_75t_L g3442 ( 
.A(n_3424),
.Y(n_3442)
);

NOR2xp33_ASAP7_75t_L g3443 ( 
.A(n_3379),
.B(n_3228),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3319),
.Y(n_3444)
);

OR2x6_ASAP7_75t_L g3445 ( 
.A(n_3397),
.B(n_3223),
.Y(n_3445)
);

INVx3_ASAP7_75t_L g3446 ( 
.A(n_3357),
.Y(n_3446)
);

CKINVDCx6p67_ASAP7_75t_R g3447 ( 
.A(n_3397),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_L g3448 ( 
.A1(n_3350),
.A2(n_3253),
.B1(n_3231),
.B2(n_3283),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3340),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3347),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3363),
.Y(n_3451)
);

HB1xp67_ASAP7_75t_L g3452 ( 
.A(n_3320),
.Y(n_3452)
);

HB1xp67_ASAP7_75t_L g3453 ( 
.A(n_3342),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3368),
.Y(n_3454)
);

BUFx2_ASAP7_75t_L g3455 ( 
.A(n_3409),
.Y(n_3455)
);

OR2x2_ASAP7_75t_L g3456 ( 
.A(n_3322),
.B(n_3271),
.Y(n_3456)
);

BUFx6f_ASAP7_75t_L g3457 ( 
.A(n_3313),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3370),
.Y(n_3458)
);

OR2x2_ASAP7_75t_L g3459 ( 
.A(n_3421),
.B(n_3223),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3374),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3384),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3385),
.Y(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_3301),
.B(n_3225),
.Y(n_3463)
);

NOR2xp33_ASAP7_75t_L g3464 ( 
.A(n_3306),
.B(n_3274),
.Y(n_3464)
);

INVx3_ASAP7_75t_L g3465 ( 
.A(n_3423),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3330),
.Y(n_3466)
);

NAND2xp33_ASAP7_75t_SL g3467 ( 
.A(n_3312),
.B(n_3276),
.Y(n_3467)
);

OAI22xp5_ASAP7_75t_SL g3468 ( 
.A1(n_3381),
.A2(n_2700),
.B1(n_2686),
.B2(n_3295),
.Y(n_3468)
);

BUFx6f_ASAP7_75t_SL g3469 ( 
.A(n_3412),
.Y(n_3469)
);

OR2x6_ASAP7_75t_L g3470 ( 
.A(n_3341),
.B(n_3181),
.Y(n_3470)
);

INVx4_ASAP7_75t_L g3471 ( 
.A(n_3315),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3332),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3377),
.Y(n_3473)
);

BUFx3_ASAP7_75t_L g3474 ( 
.A(n_3321),
.Y(n_3474)
);

NOR3xp33_ASAP7_75t_SL g3475 ( 
.A(n_3302),
.B(n_3335),
.C(n_3398),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3329),
.Y(n_3476)
);

BUFx6f_ASAP7_75t_L g3477 ( 
.A(n_3348),
.Y(n_3477)
);

HB1xp67_ASAP7_75t_L g3478 ( 
.A(n_3382),
.Y(n_3478)
);

AND2x4_ASAP7_75t_L g3479 ( 
.A(n_3430),
.B(n_3287),
.Y(n_3479)
);

HB1xp67_ASAP7_75t_L g3480 ( 
.A(n_3419),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3331),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3304),
.B(n_3257),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_SL g3483 ( 
.A(n_3310),
.B(n_3295),
.Y(n_3483)
);

INVx3_ASAP7_75t_L g3484 ( 
.A(n_3400),
.Y(n_3484)
);

INVx4_ASAP7_75t_L g3485 ( 
.A(n_3427),
.Y(n_3485)
);

BUFx8_ASAP7_75t_L g3486 ( 
.A(n_3399),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_SL g3487 ( 
.A(n_3361),
.B(n_3282),
.Y(n_3487)
);

INVx2_ASAP7_75t_SL g3488 ( 
.A(n_3428),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3333),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3403),
.B(n_3265),
.Y(n_3490)
);

AND2x4_ASAP7_75t_L g3491 ( 
.A(n_3422),
.B(n_3210),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3336),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3407),
.B(n_3268),
.Y(n_3493)
);

BUFx6f_ASAP7_75t_L g3494 ( 
.A(n_3429),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3365),
.Y(n_3495)
);

INVx2_ASAP7_75t_SL g3496 ( 
.A(n_3429),
.Y(n_3496)
);

NAND2x1p5_ASAP7_75t_L g3497 ( 
.A(n_3324),
.B(n_3203),
.Y(n_3497)
);

AO22x1_ASAP7_75t_L g3498 ( 
.A1(n_3404),
.A2(n_3418),
.B1(n_3386),
.B2(n_3372),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3344),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3367),
.Y(n_3500)
);

CKINVDCx11_ASAP7_75t_R g3501 ( 
.A(n_3345),
.Y(n_3501)
);

CKINVDCx5p33_ASAP7_75t_R g3502 ( 
.A(n_3383),
.Y(n_3502)
);

NOR3xp33_ASAP7_75t_SL g3503 ( 
.A(n_3314),
.B(n_3269),
.C(n_3241),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3354),
.B(n_3281),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3358),
.B(n_3183),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3353),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_SL g3507 ( 
.A(n_3337),
.B(n_3243),
.Y(n_3507)
);

NOR2x1_ASAP7_75t_L g3508 ( 
.A(n_3328),
.B(n_3277),
.Y(n_3508)
);

XNOR2xp5_ASAP7_75t_L g3509 ( 
.A(n_3327),
.B(n_3191),
.Y(n_3509)
);

NOR3xp33_ASAP7_75t_SL g3510 ( 
.A(n_3343),
.B(n_2892),
.C(n_1405),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3375),
.Y(n_3511)
);

NOR2xp33_ASAP7_75t_L g3512 ( 
.A(n_3359),
.B(n_3351),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3391),
.Y(n_3513)
);

INVx3_ASAP7_75t_L g3514 ( 
.A(n_3305),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3392),
.Y(n_3515)
);

AND2x4_ASAP7_75t_L g3516 ( 
.A(n_3417),
.B(n_3187),
.Y(n_3516)
);

AND2x4_ASAP7_75t_L g3517 ( 
.A(n_3390),
.B(n_3157),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3393),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3415),
.B(n_3236),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3395),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3396),
.Y(n_3521)
);

NOR2xp33_ASAP7_75t_R g3522 ( 
.A(n_3300),
.B(n_2603),
.Y(n_3522)
);

AND2x4_ASAP7_75t_L g3523 ( 
.A(n_3373),
.B(n_3151),
.Y(n_3523)
);

AND2x6_ASAP7_75t_L g3524 ( 
.A(n_3388),
.B(n_1510),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3420),
.B(n_3201),
.Y(n_3525)
);

AND2x4_ASAP7_75t_L g3526 ( 
.A(n_3376),
.B(n_3219),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3364),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3410),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3346),
.B(n_1523),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3338),
.B(n_1526),
.Y(n_3530)
);

INVx3_ASAP7_75t_L g3531 ( 
.A(n_3380),
.Y(n_3531)
);

NAND2x1p5_ASAP7_75t_L g3532 ( 
.A(n_3360),
.B(n_1546),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3405),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3411),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3413),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3355),
.B(n_3401),
.Y(n_3536)
);

INVx6_ASAP7_75t_L g3537 ( 
.A(n_3308),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3325),
.Y(n_3538)
);

BUFx6f_ASAP7_75t_L g3539 ( 
.A(n_3436),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3433),
.B(n_3402),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3512),
.B(n_3414),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3473),
.B(n_3311),
.Y(n_3542)
);

AND2x4_ASAP7_75t_L g3543 ( 
.A(n_3439),
.B(n_3326),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3456),
.B(n_3426),
.Y(n_3544)
);

BUFx12f_ASAP7_75t_L g3545 ( 
.A(n_3431),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_SL g3546 ( 
.A(n_3435),
.B(n_3303),
.Y(n_3546)
);

NOR2xp33_ASAP7_75t_L g3547 ( 
.A(n_3463),
.B(n_3408),
.Y(n_3547)
);

OAI21x1_ASAP7_75t_SL g3548 ( 
.A1(n_3536),
.A2(n_3371),
.B(n_3339),
.Y(n_3548)
);

AOI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_3519),
.A2(n_3334),
.B(n_3369),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3476),
.B(n_3349),
.Y(n_3550)
);

OAI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_3487),
.A2(n_3406),
.B(n_3356),
.Y(n_3551)
);

A2O1A1Ixp33_ASAP7_75t_L g3552 ( 
.A1(n_3475),
.A2(n_3387),
.B(n_3378),
.C(n_3389),
.Y(n_3552)
);

CKINVDCx6p67_ASAP7_75t_R g3553 ( 
.A(n_3442),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3481),
.B(n_3425),
.Y(n_3554)
);

AOI21xp5_ASAP7_75t_SL g3555 ( 
.A1(n_3525),
.A2(n_3323),
.B(n_1313),
.Y(n_3555)
);

BUFx2_ASAP7_75t_L g3556 ( 
.A(n_3484),
.Y(n_3556)
);

OAI21x1_ASAP7_75t_L g3557 ( 
.A1(n_3538),
.A2(n_1551),
.B(n_1549),
.Y(n_3557)
);

A2O1A1Ixp33_ASAP7_75t_L g3558 ( 
.A1(n_3503),
.A2(n_1560),
.B(n_1570),
.C(n_1557),
.Y(n_3558)
);

NAND3xp33_ASAP7_75t_L g3559 ( 
.A(n_3448),
.B(n_3509),
.C(n_3510),
.Y(n_3559)
);

AOI22xp5_ASAP7_75t_L g3560 ( 
.A1(n_3502),
.A2(n_1407),
.B1(n_1409),
.B2(n_1402),
.Y(n_3560)
);

BUFx2_ASAP7_75t_SL g3561 ( 
.A(n_3469),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_3535),
.A2(n_1575),
.B(n_1573),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3489),
.B(n_1410),
.Y(n_3563)
);

AND2x2_ASAP7_75t_L g3564 ( 
.A(n_3531),
.B(n_1842),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3492),
.B(n_1413),
.Y(n_3565)
);

OAI21x1_ASAP7_75t_L g3566 ( 
.A1(n_3514),
.A2(n_1589),
.B(n_1586),
.Y(n_3566)
);

OAI21x1_ASAP7_75t_L g3567 ( 
.A1(n_3528),
.A2(n_1600),
.B(n_1591),
.Y(n_3567)
);

AOI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_3482),
.A2(n_1612),
.B(n_1610),
.Y(n_3568)
);

A2O1A1Ixp33_ASAP7_75t_L g3569 ( 
.A1(n_3533),
.A2(n_1621),
.B(n_1624),
.C(n_1620),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3495),
.B(n_1414),
.Y(n_3570)
);

A2O1A1Ixp33_ASAP7_75t_L g3571 ( 
.A1(n_3527),
.A2(n_1640),
.B(n_1641),
.C(n_1625),
.Y(n_3571)
);

AO31x2_ASAP7_75t_L g3572 ( 
.A1(n_3534),
.A2(n_1648),
.A3(n_1656),
.B(n_1643),
.Y(n_3572)
);

OAI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_3529),
.A2(n_3532),
.B(n_3464),
.Y(n_3573)
);

NAND2x1p5_ASAP7_75t_L g3574 ( 
.A(n_3485),
.B(n_1657),
.Y(n_3574)
);

AO31x2_ASAP7_75t_L g3575 ( 
.A1(n_3432),
.A2(n_1668),
.A3(n_1673),
.B(n_1661),
.Y(n_3575)
);

OAI21x1_ASAP7_75t_SL g3576 ( 
.A1(n_3530),
.A2(n_1683),
.B(n_1681),
.Y(n_3576)
);

INVx3_ASAP7_75t_L g3577 ( 
.A(n_3471),
.Y(n_3577)
);

NAND2x1p5_ASAP7_75t_L g3578 ( 
.A(n_3438),
.B(n_1710),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_3500),
.A2(n_1719),
.B(n_1712),
.Y(n_3579)
);

O2A1O1Ixp5_ASAP7_75t_L g3580 ( 
.A1(n_3498),
.A2(n_1725),
.B(n_1732),
.C(n_1721),
.Y(n_3580)
);

BUFx12f_ASAP7_75t_L g3581 ( 
.A(n_3431),
.Y(n_3581)
);

INVx3_ASAP7_75t_L g3582 ( 
.A(n_3457),
.Y(n_3582)
);

CKINVDCx6p67_ASAP7_75t_R g3583 ( 
.A(n_3445),
.Y(n_3583)
);

AOI21x1_ASAP7_75t_L g3584 ( 
.A1(n_3507),
.A2(n_1743),
.B(n_1736),
.Y(n_3584)
);

OAI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_3505),
.A2(n_1758),
.B(n_1750),
.Y(n_3585)
);

BUFx6f_ASAP7_75t_L g3586 ( 
.A(n_3501),
.Y(n_3586)
);

AO31x2_ASAP7_75t_L g3587 ( 
.A1(n_3440),
.A2(n_1764),
.A3(n_1775),
.B(n_1761),
.Y(n_3587)
);

INVx2_ASAP7_75t_SL g3588 ( 
.A(n_3457),
.Y(n_3588)
);

OAI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3504),
.A2(n_1794),
.B(n_1788),
.Y(n_3589)
);

AOI21xp33_ASAP7_75t_L g3590 ( 
.A1(n_3520),
.A2(n_1803),
.B(n_1801),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3515),
.B(n_1416),
.Y(n_3591)
);

INVx2_ASAP7_75t_L g3592 ( 
.A(n_3434),
.Y(n_3592)
);

AO31x2_ASAP7_75t_L g3593 ( 
.A1(n_3441),
.A2(n_1824),
.A3(n_1827),
.B(n_1805),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3518),
.A2(n_1840),
.B(n_1834),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_SL g3595 ( 
.A1(n_3521),
.A2(n_1846),
.B(n_1845),
.Y(n_3595)
);

AOI21x1_ASAP7_75t_L g3596 ( 
.A1(n_3444),
.A2(n_1848),
.B(n_1847),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3450),
.A2(n_1858),
.B(n_1856),
.Y(n_3597)
);

OAI21x1_ASAP7_75t_L g3598 ( 
.A1(n_3449),
.A2(n_1865),
.B(n_1861),
.Y(n_3598)
);

AOI21x1_ASAP7_75t_L g3599 ( 
.A1(n_3454),
.A2(n_1883),
.B(n_1872),
.Y(n_3599)
);

OAI21x1_ASAP7_75t_L g3600 ( 
.A1(n_3461),
.A2(n_1888),
.B(n_1887),
.Y(n_3600)
);

AND2x2_ASAP7_75t_L g3601 ( 
.A(n_3491),
.B(n_1842),
.Y(n_3601)
);

AOI21xp5_ASAP7_75t_L g3602 ( 
.A1(n_3451),
.A2(n_1897),
.B(n_1896),
.Y(n_3602)
);

AOI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_3458),
.A2(n_1922),
.B(n_1903),
.Y(n_3603)
);

INVxp67_ASAP7_75t_SL g3604 ( 
.A(n_3453),
.Y(n_3604)
);

AOI21x1_ASAP7_75t_L g3605 ( 
.A1(n_3462),
.A2(n_1925),
.B(n_1923),
.Y(n_3605)
);

A2O1A1Ixp33_ASAP7_75t_L g3606 ( 
.A1(n_3508),
.A2(n_1939),
.B(n_1942),
.C(n_1932),
.Y(n_3606)
);

NOR2xp33_ASAP7_75t_L g3607 ( 
.A(n_3443),
.B(n_1417),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3537),
.B(n_1419),
.Y(n_3608)
);

OAI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3460),
.A2(n_1954),
.B(n_1946),
.Y(n_3609)
);

OAI21x1_ASAP7_75t_L g3610 ( 
.A1(n_3506),
.A2(n_1967),
.B(n_1955),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_3483),
.A2(n_1975),
.B(n_1971),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_3467),
.A2(n_1984),
.B(n_1979),
.Y(n_3612)
);

OAI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3524),
.A2(n_1995),
.B(n_1993),
.Y(n_3613)
);

AOI21x1_ASAP7_75t_L g3614 ( 
.A1(n_3490),
.A2(n_2009),
.B(n_2004),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3524),
.B(n_1422),
.Y(n_3615)
);

AOI21xp33_ASAP7_75t_SL g3616 ( 
.A1(n_3468),
.A2(n_3497),
.B(n_3496),
.Y(n_3616)
);

NAND2x1p5_ASAP7_75t_L g3617 ( 
.A(n_3494),
.B(n_2015),
.Y(n_3617)
);

OAI22xp5_ASAP7_75t_L g3618 ( 
.A1(n_3459),
.A2(n_1426),
.B1(n_1431),
.B2(n_1425),
.Y(n_3618)
);

OR2x2_ASAP7_75t_L g3619 ( 
.A(n_3452),
.B(n_2016),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3466),
.Y(n_3620)
);

INVx4_ASAP7_75t_L g3621 ( 
.A(n_3477),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3524),
.B(n_1433),
.Y(n_3622)
);

A2O1A1Ixp33_ASAP7_75t_L g3623 ( 
.A1(n_3526),
.A2(n_2021),
.B(n_2022),
.C(n_2018),
.Y(n_3623)
);

AO31x2_ASAP7_75t_L g3624 ( 
.A1(n_3472),
.A2(n_2030),
.A3(n_2044),
.B(n_2025),
.Y(n_3624)
);

BUFx6f_ASAP7_75t_L g3625 ( 
.A(n_3477),
.Y(n_3625)
);

OAI21x1_ASAP7_75t_L g3626 ( 
.A1(n_3499),
.A2(n_3513),
.B(n_3511),
.Y(n_3626)
);

OAI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3493),
.A2(n_2046),
.B(n_2045),
.Y(n_3627)
);

OAI21x1_ASAP7_75t_L g3628 ( 
.A1(n_3465),
.A2(n_2051),
.B(n_2047),
.Y(n_3628)
);

OAI21xp5_ASAP7_75t_L g3629 ( 
.A1(n_3517),
.A2(n_3516),
.B(n_3523),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3455),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_3479),
.A2(n_3446),
.B(n_3470),
.Y(n_3631)
);

BUFx2_ASAP7_75t_L g3632 ( 
.A(n_3478),
.Y(n_3632)
);

AOI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_3522),
.A2(n_2063),
.B(n_2056),
.Y(n_3633)
);

AOI21x1_ASAP7_75t_L g3634 ( 
.A1(n_3480),
.A2(n_2070),
.B(n_1057),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_SL g3635 ( 
.A(n_3437),
.B(n_1878),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_3488),
.A2(n_3494),
.B(n_3474),
.Y(n_3636)
);

OAI21x1_ASAP7_75t_L g3637 ( 
.A1(n_3447),
.A2(n_1058),
.B(n_1056),
.Y(n_3637)
);

NOR2xp67_ASAP7_75t_L g3638 ( 
.A(n_3486),
.B(n_1059),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3519),
.A2(n_1062),
.B(n_1061),
.Y(n_3639)
);

OAI21x1_ASAP7_75t_L g3640 ( 
.A1(n_3538),
.A2(n_1065),
.B(n_1063),
.Y(n_3640)
);

OAI21x1_ASAP7_75t_L g3641 ( 
.A1(n_3538),
.A2(n_1068),
.B(n_1066),
.Y(n_3641)
);

AND2x2_ASAP7_75t_SL g3642 ( 
.A(n_3464),
.B(n_1878),
.Y(n_3642)
);

OAI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3435),
.A2(n_1436),
.B(n_1434),
.Y(n_3643)
);

OAI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_3435),
.A2(n_1440),
.B(n_1437),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3434),
.Y(n_3645)
);

AOI21xp33_ASAP7_75t_L g3646 ( 
.A1(n_3536),
.A2(n_1448),
.B(n_1442),
.Y(n_3646)
);

O2A1O1Ixp5_ASAP7_75t_L g3647 ( 
.A1(n_3487),
.A2(n_1998),
.B(n_2059),
.C(n_1970),
.Y(n_3647)
);

CKINVDCx5p33_ASAP7_75t_R g3648 ( 
.A(n_3437),
.Y(n_3648)
);

NOR2xp67_ASAP7_75t_L g3649 ( 
.A(n_3484),
.B(n_1070),
.Y(n_3649)
);

BUFx4f_ASAP7_75t_L g3650 ( 
.A(n_3431),
.Y(n_3650)
);

BUFx12f_ASAP7_75t_L g3651 ( 
.A(n_3545),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3540),
.B(n_1449),
.Y(n_3652)
);

AOI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3547),
.A2(n_1453),
.B1(n_1454),
.B2(n_1452),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3645),
.Y(n_3654)
);

AND2x4_ASAP7_75t_L g3655 ( 
.A(n_3629),
.B(n_1071),
.Y(n_3655)
);

INVx6_ASAP7_75t_L g3656 ( 
.A(n_3539),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3592),
.Y(n_3657)
);

BUFx3_ASAP7_75t_L g3658 ( 
.A(n_3539),
.Y(n_3658)
);

AND2x4_ASAP7_75t_L g3659 ( 
.A(n_3632),
.B(n_1072),
.Y(n_3659)
);

AOI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3642),
.A2(n_1463),
.B1(n_1464),
.B2(n_1458),
.Y(n_3660)
);

BUFx4_ASAP7_75t_SL g3661 ( 
.A(n_3648),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3551),
.A2(n_1469),
.B(n_1466),
.Y(n_3662)
);

AOI22xp33_ASAP7_75t_L g3663 ( 
.A1(n_3559),
.A2(n_1998),
.B1(n_2059),
.B2(n_1970),
.Y(n_3663)
);

AND2x4_ASAP7_75t_L g3664 ( 
.A(n_3604),
.B(n_1073),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_SL g3665 ( 
.A(n_3573),
.B(n_1472),
.Y(n_3665)
);

INVx2_ASAP7_75t_SL g3666 ( 
.A(n_3625),
.Y(n_3666)
);

INVx3_ASAP7_75t_L g3667 ( 
.A(n_3625),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3626),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3620),
.Y(n_3669)
);

BUFx12f_ASAP7_75t_L g3670 ( 
.A(n_3581),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3575),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_SL g3672 ( 
.A(n_3541),
.B(n_1474),
.Y(n_3672)
);

AND2x4_ASAP7_75t_L g3673 ( 
.A(n_3556),
.B(n_1074),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3572),
.Y(n_3674)
);

CKINVDCx20_ASAP7_75t_R g3675 ( 
.A(n_3583),
.Y(n_3675)
);

AND2x4_ASAP7_75t_L g3676 ( 
.A(n_3582),
.B(n_1075),
.Y(n_3676)
);

AOI21xp5_ASAP7_75t_SL g3677 ( 
.A1(n_3546),
.A2(n_1479),
.B(n_1475),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_SL g3678 ( 
.A(n_3550),
.B(n_1482),
.Y(n_3678)
);

BUFx3_ASAP7_75t_L g3679 ( 
.A(n_3650),
.Y(n_3679)
);

INVxp67_ASAP7_75t_L g3680 ( 
.A(n_3630),
.Y(n_3680)
);

HB1xp67_ASAP7_75t_L g3681 ( 
.A(n_3543),
.Y(n_3681)
);

AOI22xp33_ASAP7_75t_L g3682 ( 
.A1(n_3646),
.A2(n_3544),
.B1(n_3585),
.B2(n_3590),
.Y(n_3682)
);

OR2x2_ASAP7_75t_SL g3683 ( 
.A(n_3586),
.B(n_1483),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3572),
.Y(n_3684)
);

CKINVDCx5p33_ASAP7_75t_R g3685 ( 
.A(n_3553),
.Y(n_3685)
);

AOI21xp5_ASAP7_75t_L g3686 ( 
.A1(n_3549),
.A2(n_1487),
.B(n_1486),
.Y(n_3686)
);

AOI22xp33_ASAP7_75t_L g3687 ( 
.A1(n_3589),
.A2(n_1490),
.B1(n_1494),
.B2(n_1488),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3558),
.B(n_1077),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_3542),
.A2(n_1496),
.B(n_1495),
.Y(n_3689)
);

AOI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_3635),
.A2(n_1500),
.B1(n_1501),
.B2(n_1497),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3575),
.Y(n_3691)
);

BUFx2_ASAP7_75t_L g3692 ( 
.A(n_3588),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3554),
.B(n_1507),
.Y(n_3693)
);

OR2x2_ASAP7_75t_L g3694 ( 
.A(n_3619),
.B(n_2),
.Y(n_3694)
);

NAND2xp33_ASAP7_75t_L g3695 ( 
.A(n_3552),
.B(n_1509),
.Y(n_3695)
);

BUFx2_ASAP7_75t_L g3696 ( 
.A(n_3577),
.Y(n_3696)
);

BUFx3_ASAP7_75t_L g3697 ( 
.A(n_3621),
.Y(n_3697)
);

OAI22xp5_ASAP7_75t_L g3698 ( 
.A1(n_3608),
.A2(n_1512),
.B1(n_1514),
.B2(n_1511),
.Y(n_3698)
);

OR2x6_ASAP7_75t_L g3699 ( 
.A(n_3561),
.B(n_1079),
.Y(n_3699)
);

AOI22xp5_ASAP7_75t_L g3700 ( 
.A1(n_3607),
.A2(n_1517),
.B1(n_1518),
.B2(n_1515),
.Y(n_3700)
);

INVx3_ASAP7_75t_SL g3701 ( 
.A(n_3586),
.Y(n_3701)
);

AND2x2_ASAP7_75t_L g3702 ( 
.A(n_3587),
.B(n_3593),
.Y(n_3702)
);

INVx3_ASAP7_75t_SL g3703 ( 
.A(n_3601),
.Y(n_3703)
);

AOI22xp5_ASAP7_75t_L g3704 ( 
.A1(n_3615),
.A2(n_1521),
.B1(n_1528),
.B2(n_1520),
.Y(n_3704)
);

AOI22xp33_ASAP7_75t_L g3705 ( 
.A1(n_3622),
.A2(n_1534),
.B1(n_1535),
.B2(n_1529),
.Y(n_3705)
);

BUFx3_ASAP7_75t_L g3706 ( 
.A(n_3617),
.Y(n_3706)
);

INVx4_ASAP7_75t_L g3707 ( 
.A(n_3578),
.Y(n_3707)
);

OAI22xp5_ASAP7_75t_L g3708 ( 
.A1(n_3616),
.A2(n_1539),
.B1(n_1542),
.B2(n_1537),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3563),
.B(n_1545),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3587),
.Y(n_3710)
);

AOI22xp33_ASAP7_75t_SL g3711 ( 
.A1(n_3627),
.A2(n_1561),
.B1(n_1562),
.B2(n_1552),
.Y(n_3711)
);

CKINVDCx11_ASAP7_75t_R g3712 ( 
.A(n_3618),
.Y(n_3712)
);

INVx3_ASAP7_75t_L g3713 ( 
.A(n_3584),
.Y(n_3713)
);

AND2x4_ASAP7_75t_L g3714 ( 
.A(n_3631),
.B(n_1081),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3593),
.B(n_1082),
.Y(n_3715)
);

BUFx3_ASAP7_75t_L g3716 ( 
.A(n_3564),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3624),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_3548),
.A2(n_1565),
.B(n_1563),
.Y(n_3718)
);

AND2x4_ASAP7_75t_L g3719 ( 
.A(n_3636),
.B(n_1083),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_SL g3720 ( 
.A(n_3647),
.B(n_1566),
.Y(n_3720)
);

INVx3_ASAP7_75t_SL g3721 ( 
.A(n_3638),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3624),
.Y(n_3722)
);

OR2x2_ASAP7_75t_L g3723 ( 
.A(n_3591),
.B(n_2),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3567),
.Y(n_3724)
);

AND2x4_ASAP7_75t_L g3725 ( 
.A(n_3649),
.B(n_1085),
.Y(n_3725)
);

OR2x6_ASAP7_75t_L g3726 ( 
.A(n_3595),
.B(n_1086),
.Y(n_3726)
);

NAND2x1p5_ASAP7_75t_L g3727 ( 
.A(n_3637),
.B(n_1087),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3609),
.Y(n_3728)
);

INVx2_ASAP7_75t_SL g3729 ( 
.A(n_3574),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3598),
.Y(n_3730)
);

BUFx2_ASAP7_75t_L g3731 ( 
.A(n_3610),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3580),
.B(n_1090),
.Y(n_3732)
);

O2A1O1Ixp33_ASAP7_75t_SL g3733 ( 
.A1(n_3606),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3596),
.Y(n_3734)
);

OAI22xp5_ASAP7_75t_L g3735 ( 
.A1(n_3560),
.A2(n_1568),
.B1(n_1578),
.B2(n_1567),
.Y(n_3735)
);

AND2x4_ASAP7_75t_L g3736 ( 
.A(n_3628),
.B(n_1093),
.Y(n_3736)
);

AOI22xp5_ASAP7_75t_L g3737 ( 
.A1(n_3643),
.A2(n_1582),
.B1(n_1583),
.B2(n_1579),
.Y(n_3737)
);

AOI21xp5_ASAP7_75t_L g3738 ( 
.A1(n_3555),
.A2(n_1593),
.B(n_1590),
.Y(n_3738)
);

INVxp67_ASAP7_75t_L g3739 ( 
.A(n_3565),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3600),
.Y(n_3740)
);

CKINVDCx5p33_ASAP7_75t_R g3741 ( 
.A(n_3633),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3599),
.Y(n_3742)
);

OR2x2_ASAP7_75t_L g3743 ( 
.A(n_3570),
.B(n_6),
.Y(n_3743)
);

BUFx2_ASAP7_75t_L g3744 ( 
.A(n_3566),
.Y(n_3744)
);

AND2x2_ASAP7_75t_L g3745 ( 
.A(n_3681),
.B(n_3613),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3654),
.Y(n_3746)
);

INVx2_ASAP7_75t_L g3747 ( 
.A(n_3669),
.Y(n_3747)
);

CKINVDCx5p33_ASAP7_75t_R g3748 ( 
.A(n_3661),
.Y(n_3748)
);

BUFx3_ASAP7_75t_L g3749 ( 
.A(n_3656),
.Y(n_3749)
);

NOR2xp33_ASAP7_75t_SL g3750 ( 
.A(n_3685),
.B(n_3707),
.Y(n_3750)
);

OAI22xp33_ASAP7_75t_L g3751 ( 
.A1(n_3741),
.A2(n_3639),
.B1(n_3644),
.B2(n_3612),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_3657),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3680),
.B(n_3568),
.Y(n_3753)
);

INVxp67_ASAP7_75t_L g3754 ( 
.A(n_3692),
.Y(n_3754)
);

OAI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_3682),
.A2(n_3594),
.B(n_3562),
.Y(n_3755)
);

CKINVDCx8_ASAP7_75t_R g3756 ( 
.A(n_3696),
.Y(n_3756)
);

INVxp67_ASAP7_75t_SL g3757 ( 
.A(n_3668),
.Y(n_3757)
);

BUFx3_ASAP7_75t_L g3758 ( 
.A(n_3656),
.Y(n_3758)
);

BUFx2_ASAP7_75t_L g3759 ( 
.A(n_3716),
.Y(n_3759)
);

AO21x2_ASAP7_75t_L g3760 ( 
.A1(n_3671),
.A2(n_3634),
.B(n_3605),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3691),
.Y(n_3761)
);

AOI221xp5_ASAP7_75t_L g3762 ( 
.A1(n_3733),
.A2(n_1602),
.B1(n_1603),
.B2(n_1599),
.C(n_1596),
.Y(n_3762)
);

OAI21x1_ASAP7_75t_SL g3763 ( 
.A1(n_3718),
.A2(n_3614),
.B(n_3576),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3710),
.Y(n_3764)
);

OAI21x1_ASAP7_75t_L g3765 ( 
.A1(n_3674),
.A2(n_3557),
.B(n_3640),
.Y(n_3765)
);

INVx1_ASAP7_75t_SL g3766 ( 
.A(n_3703),
.Y(n_3766)
);

OAI21x1_ASAP7_75t_L g3767 ( 
.A1(n_3684),
.A2(n_3641),
.B(n_3602),
.Y(n_3767)
);

CKINVDCx6p67_ASAP7_75t_R g3768 ( 
.A(n_3701),
.Y(n_3768)
);

AOI21xp5_ASAP7_75t_L g3769 ( 
.A1(n_3665),
.A2(n_3695),
.B(n_3678),
.Y(n_3769)
);

AOI21x1_ASAP7_75t_L g3770 ( 
.A1(n_3720),
.A2(n_3579),
.B(n_3597),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3722),
.Y(n_3771)
);

OAI21x1_ASAP7_75t_L g3772 ( 
.A1(n_3717),
.A2(n_3603),
.B(n_3611),
.Y(n_3772)
);

INVxp67_ASAP7_75t_SL g3773 ( 
.A(n_3734),
.Y(n_3773)
);

AND2x4_ASAP7_75t_L g3774 ( 
.A(n_3667),
.B(n_3569),
.Y(n_3774)
);

OR2x2_ASAP7_75t_L g3775 ( 
.A(n_3652),
.B(n_3623),
.Y(n_3775)
);

AO21x2_ASAP7_75t_L g3776 ( 
.A1(n_3702),
.A2(n_3571),
.B(n_1608),
.Y(n_3776)
);

OA21x2_ASAP7_75t_L g3777 ( 
.A1(n_3742),
.A2(n_1609),
.B(n_1606),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3728),
.Y(n_3778)
);

OAI21x1_ASAP7_75t_SL g3779 ( 
.A1(n_3686),
.A2(n_6),
.B(n_7),
.Y(n_3779)
);

OAI21x1_ASAP7_75t_L g3780 ( 
.A1(n_3730),
.A2(n_1097),
.B(n_1094),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3739),
.B(n_1611),
.Y(n_3781)
);

AO21x2_ASAP7_75t_L g3782 ( 
.A1(n_3740),
.A2(n_1617),
.B(n_1616),
.Y(n_3782)
);

BUFx2_ASAP7_75t_L g3783 ( 
.A(n_3697),
.Y(n_3783)
);

AOI22xp5_ASAP7_75t_L g3784 ( 
.A1(n_3712),
.A2(n_1623),
.B1(n_1626),
.B2(n_1622),
.Y(n_3784)
);

AOI222xp33_ASAP7_75t_L g3785 ( 
.A1(n_3663),
.A2(n_1634),
.B1(n_1631),
.B2(n_1638),
.C1(n_1633),
.C2(n_1628),
.Y(n_3785)
);

O2A1O1Ixp33_ASAP7_75t_L g3786 ( 
.A1(n_3672),
.A2(n_1647),
.B(n_1651),
.C(n_1642),
.Y(n_3786)
);

OAI21x1_ASAP7_75t_L g3787 ( 
.A1(n_3724),
.A2(n_1099),
.B(n_1098),
.Y(n_3787)
);

O2A1O1Ixp33_ASAP7_75t_SL g3788 ( 
.A1(n_3729),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_3788)
);

BUFx2_ASAP7_75t_R g3789 ( 
.A(n_3679),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3731),
.Y(n_3790)
);

OAI21x1_ASAP7_75t_L g3791 ( 
.A1(n_3713),
.A2(n_1102),
.B(n_1100),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3664),
.Y(n_3792)
);

CKINVDCx20_ASAP7_75t_R g3793 ( 
.A(n_3675),
.Y(n_3793)
);

OAI21x1_ASAP7_75t_L g3794 ( 
.A1(n_3727),
.A2(n_1104),
.B(n_1103),
.Y(n_3794)
);

AO21x2_ASAP7_75t_L g3795 ( 
.A1(n_3662),
.A2(n_1659),
.B(n_1658),
.Y(n_3795)
);

NAND2x1p5_ASAP7_75t_L g3796 ( 
.A(n_3714),
.B(n_3655),
.Y(n_3796)
);

AOI22xp33_ASAP7_75t_L g3797 ( 
.A1(n_3688),
.A2(n_1662),
.B1(n_1666),
.B2(n_1660),
.Y(n_3797)
);

INVx3_ASAP7_75t_L g3798 ( 
.A(n_3658),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3744),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3715),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3723),
.Y(n_3801)
);

AOI22xp5_ASAP7_75t_L g3802 ( 
.A1(n_3726),
.A2(n_1670),
.B1(n_1671),
.B2(n_1669),
.Y(n_3802)
);

OAI21x1_ASAP7_75t_L g3803 ( 
.A1(n_3732),
.A2(n_1106),
.B(n_1105),
.Y(n_3803)
);

OAI22xp5_ASAP7_75t_L g3804 ( 
.A1(n_3660),
.A2(n_1678),
.B1(n_1680),
.B2(n_1674),
.Y(n_3804)
);

AOI22xp5_ASAP7_75t_L g3805 ( 
.A1(n_3726),
.A2(n_3719),
.B1(n_3699),
.B2(n_3653),
.Y(n_3805)
);

AOI22xp33_ASAP7_75t_L g3806 ( 
.A1(n_3689),
.A2(n_1686),
.B1(n_1687),
.B2(n_1685),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3743),
.Y(n_3807)
);

OAI21x1_ASAP7_75t_L g3808 ( 
.A1(n_3738),
.A2(n_1109),
.B(n_1108),
.Y(n_3808)
);

AOI21xp33_ASAP7_75t_L g3809 ( 
.A1(n_3693),
.A2(n_1691),
.B(n_1688),
.Y(n_3809)
);

OAI21x1_ASAP7_75t_L g3810 ( 
.A1(n_3677),
.A2(n_1111),
.B(n_1110),
.Y(n_3810)
);

OA21x2_ASAP7_75t_L g3811 ( 
.A1(n_3736),
.A2(n_3709),
.B(n_3725),
.Y(n_3811)
);

HB1xp67_ASAP7_75t_L g3812 ( 
.A(n_3666),
.Y(n_3812)
);

OAI21x1_ASAP7_75t_L g3813 ( 
.A1(n_3708),
.A2(n_1115),
.B(n_1114),
.Y(n_3813)
);

O2A1O1Ixp33_ASAP7_75t_SL g3814 ( 
.A1(n_3694),
.A2(n_18),
.B(n_30),
.C(n_8),
.Y(n_3814)
);

AO31x2_ASAP7_75t_L g3815 ( 
.A1(n_3698),
.A2(n_12),
.A3(n_10),
.B(n_11),
.Y(n_3815)
);

AO21x2_ASAP7_75t_L g3816 ( 
.A1(n_3737),
.A2(n_1694),
.B(n_1692),
.Y(n_3816)
);

AND2x2_ASAP7_75t_L g3817 ( 
.A(n_3659),
.B(n_11),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3673),
.Y(n_3818)
);

OAI21x1_ASAP7_75t_L g3819 ( 
.A1(n_3705),
.A2(n_1117),
.B(n_1116),
.Y(n_3819)
);

AND2x2_ASAP7_75t_L g3820 ( 
.A(n_3676),
.B(n_12),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3706),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3759),
.B(n_3766),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_SL g3823 ( 
.A(n_3751),
.B(n_3721),
.Y(n_3823)
);

OAI21x1_ASAP7_75t_L g3824 ( 
.A1(n_3765),
.A2(n_3704),
.B(n_3735),
.Y(n_3824)
);

OAI22xp5_ASAP7_75t_L g3825 ( 
.A1(n_3797),
.A2(n_3699),
.B1(n_3683),
.B2(n_3711),
.Y(n_3825)
);

INVx3_ASAP7_75t_L g3826 ( 
.A(n_3756),
.Y(n_3826)
);

AOI221xp5_ASAP7_75t_L g3827 ( 
.A1(n_3814),
.A2(n_3687),
.B1(n_1701),
.B2(n_1702),
.C(n_1698),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3801),
.B(n_3651),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3746),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3761),
.Y(n_3830)
);

NAND3xp33_ASAP7_75t_L g3831 ( 
.A(n_3755),
.B(n_3700),
.C(n_3690),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3764),
.Y(n_3832)
);

BUFx6f_ASAP7_75t_L g3833 ( 
.A(n_3749),
.Y(n_3833)
);

OAI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3769),
.A2(n_1705),
.B(n_1695),
.Y(n_3834)
);

OR2x2_ASAP7_75t_L g3835 ( 
.A(n_3799),
.B(n_13),
.Y(n_3835)
);

OAI22xp5_ASAP7_75t_L g3836 ( 
.A1(n_3805),
.A2(n_3670),
.B1(n_1708),
.B2(n_1709),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3807),
.B(n_3783),
.Y(n_3837)
);

OAI22xp5_ASAP7_75t_L g3838 ( 
.A1(n_3802),
.A2(n_1714),
.B1(n_1715),
.B2(n_1707),
.Y(n_3838)
);

OAI22xp33_ASAP7_75t_L g3839 ( 
.A1(n_3750),
.A2(n_2083),
.B1(n_2084),
.B2(n_2082),
.Y(n_3839)
);

CKINVDCx14_ASAP7_75t_R g3840 ( 
.A(n_3748),
.Y(n_3840)
);

INVx3_ASAP7_75t_L g3841 ( 
.A(n_3798),
.Y(n_3841)
);

AOI222xp33_ASAP7_75t_L g3842 ( 
.A1(n_3762),
.A2(n_1728),
.B1(n_1726),
.B2(n_1730),
.C1(n_1727),
.C2(n_1716),
.Y(n_3842)
);

AOI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_3811),
.A2(n_1735),
.B1(n_1737),
.B2(n_1731),
.Y(n_3843)
);

AOI22xp33_ASAP7_75t_L g3844 ( 
.A1(n_3795),
.A2(n_1741),
.B1(n_1747),
.B2(n_1738),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_3754),
.B(n_3821),
.Y(n_3845)
);

AOI22xp33_ASAP7_75t_L g3846 ( 
.A1(n_3816),
.A2(n_1759),
.B1(n_1760),
.B2(n_1754),
.Y(n_3846)
);

INVx2_ASAP7_75t_L g3847 ( 
.A(n_3752),
.Y(n_3847)
);

INVx2_ASAP7_75t_SL g3848 ( 
.A(n_3812),
.Y(n_3848)
);

OAI22xp5_ASAP7_75t_L g3849 ( 
.A1(n_3775),
.A2(n_1770),
.B1(n_1773),
.B2(n_1762),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_SL g3850 ( 
.A(n_3753),
.B(n_1774),
.Y(n_3850)
);

INVxp33_ASAP7_75t_SL g3851 ( 
.A(n_3784),
.Y(n_3851)
);

NAND2xp33_ASAP7_75t_SL g3852 ( 
.A(n_3793),
.B(n_1777),
.Y(n_3852)
);

BUFx2_ASAP7_75t_L g3853 ( 
.A(n_3768),
.Y(n_3853)
);

AOI222xp33_ASAP7_75t_L g3854 ( 
.A1(n_3804),
.A2(n_1785),
.B1(n_1783),
.B2(n_1786),
.C1(n_1784),
.C2(n_1781),
.Y(n_3854)
);

AOI221xp5_ASAP7_75t_L g3855 ( 
.A1(n_3788),
.A2(n_2066),
.B1(n_2069),
.B2(n_2058),
.C(n_2057),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3745),
.B(n_13),
.Y(n_3856)
);

OAI22xp5_ASAP7_75t_L g3857 ( 
.A1(n_3796),
.A2(n_1791),
.B1(n_1793),
.B2(n_1789),
.Y(n_3857)
);

AND2x2_ASAP7_75t_L g3858 ( 
.A(n_3747),
.B(n_14),
.Y(n_3858)
);

AND2x6_ASAP7_75t_L g3859 ( 
.A(n_3774),
.B(n_1118),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3778),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3800),
.B(n_14),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3771),
.Y(n_3862)
);

AOI22xp33_ASAP7_75t_L g3863 ( 
.A1(n_3776),
.A2(n_1798),
.B1(n_1804),
.B2(n_1796),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3773),
.B(n_1808),
.Y(n_3864)
);

HB1xp67_ASAP7_75t_L g3865 ( 
.A(n_3790),
.Y(n_3865)
);

INVx4_ASAP7_75t_L g3866 ( 
.A(n_3758),
.Y(n_3866)
);

BUFx2_ASAP7_75t_L g3867 ( 
.A(n_3792),
.Y(n_3867)
);

OR2x2_ASAP7_75t_L g3868 ( 
.A(n_3757),
.B(n_16),
.Y(n_3868)
);

NAND3xp33_ASAP7_75t_SL g3869 ( 
.A(n_3785),
.B(n_1810),
.C(n_1809),
.Y(n_3869)
);

AOI22xp5_ASAP7_75t_L g3870 ( 
.A1(n_3782),
.A2(n_1817),
.B1(n_1819),
.B2(n_1814),
.Y(n_3870)
);

AO31x2_ASAP7_75t_L g3871 ( 
.A1(n_3760),
.A2(n_3818),
.A3(n_3781),
.B(n_3767),
.Y(n_3871)
);

AO31x2_ASAP7_75t_L g3872 ( 
.A1(n_3815),
.A2(n_18),
.A3(n_16),
.B(n_17),
.Y(n_3872)
);

CKINVDCx8_ASAP7_75t_R g3873 ( 
.A(n_3789),
.Y(n_3873)
);

AO31x2_ASAP7_75t_L g3874 ( 
.A1(n_3815),
.A2(n_21),
.A3(n_17),
.B(n_19),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3777),
.B(n_1826),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3817),
.B(n_1828),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3772),
.Y(n_3877)
);

OAI222xp33_ASAP7_75t_L g3878 ( 
.A1(n_3806),
.A2(n_1841),
.B1(n_1836),
.B2(n_1843),
.C1(n_1839),
.C2(n_1829),
.Y(n_3878)
);

OAI22xp5_ASAP7_75t_L g3879 ( 
.A1(n_3770),
.A2(n_1849),
.B1(n_1851),
.B2(n_1844),
.Y(n_3879)
);

AND2x4_ASAP7_75t_SL g3880 ( 
.A(n_3820),
.B(n_1119),
.Y(n_3880)
);

NAND3xp33_ASAP7_75t_L g3881 ( 
.A(n_3809),
.B(n_1860),
.C(n_1857),
.Y(n_3881)
);

HB1xp67_ASAP7_75t_L g3882 ( 
.A(n_3803),
.Y(n_3882)
);

OR2x2_ASAP7_75t_L g3883 ( 
.A(n_3791),
.B(n_19),
.Y(n_3883)
);

AND2x4_ASAP7_75t_L g3884 ( 
.A(n_3794),
.B(n_1120),
.Y(n_3884)
);

NOR2xp33_ASAP7_75t_L g3885 ( 
.A(n_3786),
.B(n_1864),
.Y(n_3885)
);

AOI22xp33_ASAP7_75t_SL g3886 ( 
.A1(n_3779),
.A2(n_1869),
.B1(n_1870),
.B2(n_1867),
.Y(n_3886)
);

NAND2xp33_ASAP7_75t_SL g3887 ( 
.A(n_3810),
.B(n_1873),
.Y(n_3887)
);

OR2x2_ASAP7_75t_L g3888 ( 
.A(n_3813),
.B(n_22),
.Y(n_3888)
);

AND2x6_ASAP7_75t_L g3889 ( 
.A(n_3819),
.B(n_22),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3787),
.Y(n_3890)
);

BUFx12f_ASAP7_75t_L g3891 ( 
.A(n_3808),
.Y(n_3891)
);

AOI22xp33_ASAP7_75t_L g3892 ( 
.A1(n_3763),
.A2(n_1879),
.B1(n_1880),
.B2(n_1876),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3780),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_L g3894 ( 
.A(n_3752),
.B(n_1884),
.Y(n_3894)
);

INVx3_ASAP7_75t_L g3895 ( 
.A(n_3841),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3829),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3847),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3848),
.Y(n_3898)
);

AND2x2_ASAP7_75t_L g3899 ( 
.A(n_3822),
.B(n_23),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3830),
.Y(n_3900)
);

AOI22xp33_ASAP7_75t_L g3901 ( 
.A1(n_3831),
.A2(n_2054),
.B1(n_2055),
.B2(n_2053),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3832),
.Y(n_3902)
);

AO21x2_ASAP7_75t_L g3903 ( 
.A1(n_3877),
.A2(n_25),
.B(n_27),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_3865),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3860),
.Y(n_3905)
);

INVx3_ASAP7_75t_L g3906 ( 
.A(n_3866),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3862),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3837),
.B(n_1885),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3867),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_3845),
.B(n_25),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3871),
.Y(n_3911)
);

INVx2_ASAP7_75t_L g3912 ( 
.A(n_3871),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3828),
.B(n_27),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3868),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3890),
.Y(n_3915)
);

OA21x2_ASAP7_75t_L g3916 ( 
.A1(n_3824),
.A2(n_3823),
.B(n_3864),
.Y(n_3916)
);

AND2x2_ASAP7_75t_L g3917 ( 
.A(n_3826),
.B(n_29),
.Y(n_3917)
);

INVx3_ASAP7_75t_L g3918 ( 
.A(n_3833),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3853),
.B(n_30),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3893),
.Y(n_3920)
);

AND2x2_ASAP7_75t_L g3921 ( 
.A(n_3833),
.B(n_31),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3835),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3882),
.Y(n_3923)
);

BUFx3_ASAP7_75t_L g3924 ( 
.A(n_3873),
.Y(n_3924)
);

INVx2_ASAP7_75t_SL g3925 ( 
.A(n_3858),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3883),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3872),
.Y(n_3927)
);

INVx5_ASAP7_75t_L g3928 ( 
.A(n_3859),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3856),
.B(n_32),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3872),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3888),
.Y(n_3931)
);

HB1xp67_ASAP7_75t_L g3932 ( 
.A(n_3874),
.Y(n_3932)
);

OAI21x1_ASAP7_75t_L g3933 ( 
.A1(n_3879),
.A2(n_32),
.B(n_33),
.Y(n_3933)
);

AND2x4_ASAP7_75t_L g3934 ( 
.A(n_3861),
.B(n_34),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3874),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3894),
.Y(n_3936)
);

AND2x2_ASAP7_75t_L g3937 ( 
.A(n_3840),
.B(n_34),
.Y(n_3937)
);

INVx2_ASAP7_75t_L g3938 ( 
.A(n_3891),
.Y(n_3938)
);

O2A1O1Ixp5_ASAP7_75t_L g3939 ( 
.A1(n_3887),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_3939)
);

INVx6_ASAP7_75t_L g3940 ( 
.A(n_3859),
.Y(n_3940)
);

HB1xp67_ASAP7_75t_L g3941 ( 
.A(n_3875),
.Y(n_3941)
);

OR2x2_ASAP7_75t_L g3942 ( 
.A(n_3876),
.B(n_3836),
.Y(n_3942)
);

NOR2xp33_ASAP7_75t_L g3943 ( 
.A(n_3851),
.B(n_3850),
.Y(n_3943)
);

BUFx2_ASAP7_75t_L g3944 ( 
.A(n_3859),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3843),
.Y(n_3945)
);

INVxp67_ASAP7_75t_L g3946 ( 
.A(n_3889),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3889),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3884),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3870),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3880),
.Y(n_3950)
);

OA21x2_ASAP7_75t_L g3951 ( 
.A1(n_3863),
.A2(n_1889),
.B(n_1886),
.Y(n_3951)
);

OAI21xp5_ASAP7_75t_L g3952 ( 
.A1(n_3834),
.A2(n_3825),
.B(n_3846),
.Y(n_3952)
);

INVx5_ASAP7_75t_L g3953 ( 
.A(n_3852),
.Y(n_3953)
);

OAI21x1_ASAP7_75t_L g3954 ( 
.A1(n_3857),
.A2(n_37),
.B(n_38),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3849),
.Y(n_3955)
);

NOR2xp33_ASAP7_75t_L g3956 ( 
.A(n_3839),
.B(n_1891),
.Y(n_3956)
);

BUFx3_ASAP7_75t_L g3957 ( 
.A(n_3881),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3892),
.Y(n_3958)
);

AOI21x1_ASAP7_75t_L g3959 ( 
.A1(n_3838),
.A2(n_1898),
.B(n_1892),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3886),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3896),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3923),
.Y(n_3962)
);

HB1xp67_ASAP7_75t_L g3963 ( 
.A(n_3920),
.Y(n_3963)
);

INVx2_ASAP7_75t_L g3964 ( 
.A(n_3931),
.Y(n_3964)
);

OA21x2_ASAP7_75t_L g3965 ( 
.A1(n_3911),
.A2(n_3844),
.B(n_3855),
.Y(n_3965)
);

AOI22xp33_ASAP7_75t_L g3966 ( 
.A1(n_3952),
.A2(n_3869),
.B1(n_3827),
.B2(n_3885),
.Y(n_3966)
);

BUFx2_ASAP7_75t_L g3967 ( 
.A(n_3944),
.Y(n_3967)
);

OAI21x1_ASAP7_75t_L g3968 ( 
.A1(n_3912),
.A2(n_3878),
.B(n_3842),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3900),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3909),
.B(n_39),
.Y(n_3970)
);

OAI221xp5_ASAP7_75t_L g3971 ( 
.A1(n_3901),
.A2(n_3854),
.B1(n_1902),
.B2(n_1910),
.C(n_1901),
.Y(n_3971)
);

AND2x2_ASAP7_75t_L g3972 ( 
.A(n_3895),
.B(n_39),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3926),
.B(n_40),
.Y(n_3973)
);

OAI221xp5_ASAP7_75t_L g3974 ( 
.A1(n_3945),
.A2(n_3949),
.B1(n_3946),
.B2(n_3941),
.C(n_3958),
.Y(n_3974)
);

AOI22xp33_ASAP7_75t_L g3975 ( 
.A1(n_3957),
.A2(n_1913),
.B1(n_1915),
.B2(n_1899),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3902),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3904),
.B(n_1916),
.Y(n_3977)
);

INVx3_ASAP7_75t_L g3978 ( 
.A(n_3906),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3922),
.B(n_40),
.Y(n_3979)
);

AOI22xp33_ASAP7_75t_L g3980 ( 
.A1(n_3960),
.A2(n_1921),
.B1(n_1924),
.B2(n_1917),
.Y(n_3980)
);

AOI22xp33_ASAP7_75t_L g3981 ( 
.A1(n_3916),
.A2(n_1933),
.B1(n_1935),
.B2(n_1928),
.Y(n_3981)
);

NAND4xp25_ASAP7_75t_L g3982 ( 
.A(n_3956),
.B(n_44),
.C(n_42),
.D(n_43),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3905),
.Y(n_3983)
);

AOI33xp33_ASAP7_75t_L g3984 ( 
.A1(n_3955),
.A2(n_1941),
.A3(n_1937),
.B1(n_1947),
.B2(n_1938),
.B3(n_1936),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3915),
.Y(n_3985)
);

AOI22xp33_ASAP7_75t_L g3986 ( 
.A1(n_3947),
.A2(n_1956),
.B1(n_1959),
.B2(n_1948),
.Y(n_3986)
);

OAI221xp5_ASAP7_75t_L g3987 ( 
.A1(n_3943),
.A2(n_1963),
.B1(n_1977),
.B2(n_1961),
.C(n_1960),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3936),
.B(n_1980),
.Y(n_3988)
);

AOI22xp33_ASAP7_75t_SL g3989 ( 
.A1(n_3928),
.A2(n_1989),
.B1(n_1990),
.B2(n_1986),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3914),
.B(n_1992),
.Y(n_3990)
);

AOI21xp5_ASAP7_75t_L g3991 ( 
.A1(n_3939),
.A2(n_2014),
.B(n_2000),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3951),
.A2(n_1999),
.B1(n_2005),
.B2(n_1994),
.Y(n_3992)
);

AOI22xp5_ASAP7_75t_L g3993 ( 
.A1(n_3928),
.A2(n_2008),
.B1(n_2010),
.B2(n_2007),
.Y(n_3993)
);

AOI221xp5_ASAP7_75t_SL g3994 ( 
.A1(n_3927),
.A2(n_3930),
.B1(n_3935),
.B2(n_3942),
.C(n_3938),
.Y(n_3994)
);

INVx3_ASAP7_75t_L g3995 ( 
.A(n_3918),
.Y(n_3995)
);

AND2x2_ASAP7_75t_L g3996 ( 
.A(n_3898),
.B(n_42),
.Y(n_3996)
);

OAI211xp5_ASAP7_75t_L g3997 ( 
.A1(n_3932),
.A2(n_2012),
.B(n_2013),
.C(n_2011),
.Y(n_3997)
);

OAI22xp5_ASAP7_75t_L g3998 ( 
.A1(n_3940),
.A2(n_2020),
.B1(n_2028),
.B2(n_2017),
.Y(n_3998)
);

OAI211xp5_ASAP7_75t_L g3999 ( 
.A1(n_3959),
.A2(n_2031),
.B(n_2032),
.C(n_2029),
.Y(n_3999)
);

AOI221xp5_ASAP7_75t_L g4000 ( 
.A1(n_3908),
.A2(n_2040),
.B1(n_2041),
.B2(n_2039),
.C(n_2037),
.Y(n_4000)
);

OAI22xp5_ASAP7_75t_L g4001 ( 
.A1(n_3948),
.A2(n_2048),
.B1(n_2050),
.B2(n_2042),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3907),
.Y(n_4002)
);

AOI21xp5_ASAP7_75t_L g4003 ( 
.A1(n_3903),
.A2(n_2078),
.B(n_2072),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3925),
.B(n_43),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3897),
.Y(n_4005)
);

AOI222xp33_ASAP7_75t_L g4006 ( 
.A1(n_3953),
.A2(n_3933),
.B1(n_3954),
.B2(n_3919),
.C1(n_3917),
.C2(n_3937),
.Y(n_4006)
);

AOI221xp5_ASAP7_75t_L g4007 ( 
.A1(n_3910),
.A2(n_2079),
.B1(n_2085),
.B2(n_2077),
.C(n_2052),
.Y(n_4007)
);

AOI22xp33_ASAP7_75t_L g4008 ( 
.A1(n_3953),
.A2(n_2088),
.B1(n_2087),
.B2(n_46),
.Y(n_4008)
);

NAND3xp33_ASAP7_75t_L g4009 ( 
.A(n_3899),
.B(n_44),
.C(n_45),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3929),
.B(n_3934),
.Y(n_4010)
);

AOI221xp5_ASAP7_75t_L g4011 ( 
.A1(n_3921),
.A2(n_48),
.B1(n_45),
.B2(n_47),
.C(n_49),
.Y(n_4011)
);

AOI221xp5_ASAP7_75t_L g4012 ( 
.A1(n_3913),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.C(n_50),
.Y(n_4012)
);

AOI221xp5_ASAP7_75t_L g4013 ( 
.A1(n_3924),
.A2(n_53),
.B1(n_50),
.B2(n_51),
.C(n_54),
.Y(n_4013)
);

OAI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_3950),
.A2(n_51),
.B(n_53),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3923),
.Y(n_4015)
);

OAI22xp5_ASAP7_75t_L g4016 ( 
.A1(n_3928),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_4016)
);

OAI211xp5_ASAP7_75t_L g4017 ( 
.A1(n_3952),
.A2(n_58),
.B(n_55),
.C(n_57),
.Y(n_4017)
);

AOI21xp5_ASAP7_75t_L g4018 ( 
.A1(n_3952),
.A2(n_57),
.B(n_61),
.Y(n_4018)
);

OR2x2_ASAP7_75t_L g4019 ( 
.A(n_3904),
.B(n_61),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3923),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3941),
.B(n_63),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3923),
.Y(n_4022)
);

OAI22xp5_ASAP7_75t_L g4023 ( 
.A1(n_3928),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_3909),
.B(n_64),
.Y(n_4024)
);

OR2x2_ASAP7_75t_L g4025 ( 
.A(n_3904),
.B(n_65),
.Y(n_4025)
);

BUFx6f_ASAP7_75t_L g4026 ( 
.A(n_3918),
.Y(n_4026)
);

AOI221xp5_ASAP7_75t_L g4027 ( 
.A1(n_3952),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.C(n_69),
.Y(n_4027)
);

OAI21x1_ASAP7_75t_L g4028 ( 
.A1(n_3912),
.A2(n_66),
.B(n_69),
.Y(n_4028)
);

OAI22xp5_ASAP7_75t_L g4029 ( 
.A1(n_3928),
.A2(n_74),
.B1(n_71),
.B2(n_72),
.Y(n_4029)
);

AOI22xp33_ASAP7_75t_L g4030 ( 
.A1(n_3952),
.A2(n_76),
.B1(n_72),
.B2(n_75),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3909),
.B(n_75),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3923),
.Y(n_4032)
);

AO21x2_ASAP7_75t_L g4033 ( 
.A1(n_3911),
.A2(n_76),
.B(n_77),
.Y(n_4033)
);

NAND3xp33_ASAP7_75t_L g4034 ( 
.A(n_3952),
.B(n_77),
.C(n_78),
.Y(n_4034)
);

AOI22xp33_ASAP7_75t_SL g4035 ( 
.A1(n_3952),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3896),
.Y(n_4036)
);

HB1xp67_ASAP7_75t_L g4037 ( 
.A(n_3920),
.Y(n_4037)
);

OR2x2_ASAP7_75t_L g4038 ( 
.A(n_3904),
.B(n_79),
.Y(n_4038)
);

NAND4xp25_ASAP7_75t_L g4039 ( 
.A(n_3952),
.B(n_83),
.C(n_80),
.D(n_82),
.Y(n_4039)
);

AOI22xp33_ASAP7_75t_L g4040 ( 
.A1(n_3952),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_4040)
);

AOI21xp5_ASAP7_75t_L g4041 ( 
.A1(n_3952),
.A2(n_84),
.B(n_85),
.Y(n_4041)
);

OA21x2_ASAP7_75t_L g4042 ( 
.A1(n_3911),
.A2(n_86),
.B(n_87),
.Y(n_4042)
);

AOI221xp5_ASAP7_75t_L g4043 ( 
.A1(n_3952),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.C(n_92),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3896),
.Y(n_4044)
);

OAI21x1_ASAP7_75t_L g4045 ( 
.A1(n_3912),
.A2(n_89),
.B(n_91),
.Y(n_4045)
);

NAND3xp33_ASAP7_75t_L g4046 ( 
.A(n_3952),
.B(n_93),
.C(n_94),
.Y(n_4046)
);

OAI21x1_ASAP7_75t_L g4047 ( 
.A1(n_3912),
.A2(n_93),
.B(n_95),
.Y(n_4047)
);

AOI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3952),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_4048)
);

AOI22xp33_ASAP7_75t_SL g4049 ( 
.A1(n_3952),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_4049)
);

AOI322xp5_ASAP7_75t_L g4050 ( 
.A1(n_3960),
.A2(n_104),
.A3(n_103),
.B1(n_101),
.B2(n_99),
.C1(n_100),
.C2(n_102),
.Y(n_4050)
);

AOI21x1_ASAP7_75t_L g4051 ( 
.A1(n_3941),
.A2(n_100),
.B(n_104),
.Y(n_4051)
);

AOI222xp33_ASAP7_75t_L g4052 ( 
.A1(n_3952),
.A2(n_107),
.B1(n_109),
.B2(n_105),
.C1(n_106),
.C2(n_108),
.Y(n_4052)
);

INVx2_ASAP7_75t_L g4053 ( 
.A(n_3923),
.Y(n_4053)
);

OAI211xp5_ASAP7_75t_L g4054 ( 
.A1(n_3952),
.A2(n_109),
.B(n_106),
.C(n_108),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3941),
.B(n_110),
.Y(n_4055)
);

OA21x2_ASAP7_75t_L g4056 ( 
.A1(n_3911),
.A2(n_110),
.B(n_111),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3896),
.Y(n_4057)
);

OAI211xp5_ASAP7_75t_L g4058 ( 
.A1(n_3952),
.A2(n_114),
.B(n_112),
.C(n_113),
.Y(n_4058)
);

OAI22xp5_ASAP7_75t_L g4059 ( 
.A1(n_3928),
.A2(n_115),
.B1(n_112),
.B2(n_113),
.Y(n_4059)
);

AND2x2_ASAP7_75t_L g4060 ( 
.A(n_3909),
.B(n_116),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3896),
.Y(n_4061)
);

AOI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_3952),
.A2(n_116),
.B(n_117),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3896),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3941),
.B(n_117),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3896),
.Y(n_4065)
);

OAI221xp5_ASAP7_75t_L g4066 ( 
.A1(n_3952),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.C(n_121),
.Y(n_4066)
);

OAI221xp5_ASAP7_75t_L g4067 ( 
.A1(n_3952),
.A2(n_123),
.B1(n_118),
.B2(n_122),
.C(n_124),
.Y(n_4067)
);

OAI21x1_ASAP7_75t_L g4068 ( 
.A1(n_3912),
.A2(n_123),
.B(n_125),
.Y(n_4068)
);

AOI222xp33_ASAP7_75t_L g4069 ( 
.A1(n_3952),
.A2(n_127),
.B1(n_129),
.B2(n_125),
.C1(n_126),
.C2(n_128),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3896),
.Y(n_4070)
);

AOI22xp33_ASAP7_75t_L g4071 ( 
.A1(n_3952),
.A2(n_130),
.B1(n_127),
.B2(n_128),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_3923),
.Y(n_4072)
);

AOI221xp5_ASAP7_75t_L g4073 ( 
.A1(n_3952),
.A2(n_133),
.B1(n_130),
.B2(n_132),
.C(n_134),
.Y(n_4073)
);

INVx2_ASAP7_75t_L g4074 ( 
.A(n_3923),
.Y(n_4074)
);

OR2x2_ASAP7_75t_L g4075 ( 
.A(n_3904),
.B(n_132),
.Y(n_4075)
);

AND2x2_ASAP7_75t_L g4076 ( 
.A(n_3909),
.B(n_133),
.Y(n_4076)
);

AOI22xp5_ASAP7_75t_L g4077 ( 
.A1(n_3952),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_4077)
);

AOI22xp5_ASAP7_75t_L g4078 ( 
.A1(n_3952),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_4078)
);

HB1xp67_ASAP7_75t_L g4079 ( 
.A(n_3963),
.Y(n_4079)
);

AND2x2_ASAP7_75t_L g4080 ( 
.A(n_3967),
.B(n_138),
.Y(n_4080)
);

AND2x2_ASAP7_75t_L g4081 ( 
.A(n_3978),
.B(n_138),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_3995),
.B(n_139),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3961),
.Y(n_4083)
);

NOR2x1_ASAP7_75t_L g4084 ( 
.A(n_3974),
.B(n_139),
.Y(n_4084)
);

NAND2x1_ASAP7_75t_L g4085 ( 
.A(n_3962),
.B(n_141),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_3964),
.B(n_140),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_3976),
.Y(n_4087)
);

OR2x2_ASAP7_75t_L g4088 ( 
.A(n_4002),
.B(n_141),
.Y(n_4088)
);

NAND2x1p5_ASAP7_75t_L g4089 ( 
.A(n_4026),
.B(n_142),
.Y(n_4089)
);

INVx2_ASAP7_75t_SL g4090 ( 
.A(n_4026),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3994),
.B(n_143),
.Y(n_4091)
);

AND2x2_ASAP7_75t_L g4092 ( 
.A(n_4015),
.B(n_143),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_3969),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_4020),
.B(n_144),
.Y(n_4094)
);

INVx2_ASAP7_75t_L g4095 ( 
.A(n_4022),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3983),
.Y(n_4096)
);

OR2x2_ASAP7_75t_L g4097 ( 
.A(n_4005),
.B(n_4019),
.Y(n_4097)
);

INVxp33_ASAP7_75t_L g4098 ( 
.A(n_3968),
.Y(n_4098)
);

INVxp67_ASAP7_75t_SL g4099 ( 
.A(n_4037),
.Y(n_4099)
);

AND2x2_ASAP7_75t_L g4100 ( 
.A(n_4032),
.B(n_144),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_4036),
.Y(n_4101)
);

INVx4_ASAP7_75t_L g4102 ( 
.A(n_3972),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4044),
.Y(n_4103)
);

AOI22xp33_ASAP7_75t_L g4104 ( 
.A1(n_3966),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_4053),
.B(n_4072),
.Y(n_4105)
);

INVx4_ASAP7_75t_L g4106 ( 
.A(n_4004),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_4074),
.B(n_145),
.Y(n_4107)
);

OR2x2_ASAP7_75t_L g4108 ( 
.A(n_4025),
.B(n_146),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_4006),
.B(n_147),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_3970),
.B(n_148),
.Y(n_4110)
);

BUFx6f_ASAP7_75t_L g4111 ( 
.A(n_4024),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_4057),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4061),
.Y(n_4113)
);

AND2x4_ASAP7_75t_L g4114 ( 
.A(n_4031),
.B(n_149),
.Y(n_4114)
);

NOR2xp33_ASAP7_75t_L g4115 ( 
.A(n_4021),
.B(n_150),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_4063),
.Y(n_4116)
);

INVxp67_ASAP7_75t_L g4117 ( 
.A(n_3990),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_4065),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_4060),
.B(n_4076),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_4070),
.Y(n_4120)
);

AND2x4_ASAP7_75t_L g4121 ( 
.A(n_3996),
.B(n_150),
.Y(n_4121)
);

AND2x2_ASAP7_75t_L g4122 ( 
.A(n_3979),
.B(n_151),
.Y(n_4122)
);

NOR2xp33_ASAP7_75t_L g4123 ( 
.A(n_4055),
.B(n_151),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3985),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4042),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4042),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_4038),
.B(n_152),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_4056),
.Y(n_4128)
);

INVxp67_ASAP7_75t_SL g4129 ( 
.A(n_4056),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_4075),
.B(n_152),
.Y(n_4130)
);

OR2x2_ASAP7_75t_L g4131 ( 
.A(n_4064),
.B(n_153),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3977),
.Y(n_4132)
);

AND2x4_ASAP7_75t_L g4133 ( 
.A(n_3973),
.B(n_154),
.Y(n_4133)
);

AND2x4_ASAP7_75t_L g4134 ( 
.A(n_4010),
.B(n_154),
.Y(n_4134)
);

AOI22xp5_ASAP7_75t_L g4135 ( 
.A1(n_4039),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_4135)
);

AND2x2_ASAP7_75t_L g4136 ( 
.A(n_3965),
.B(n_3981),
.Y(n_4136)
);

INVxp67_ASAP7_75t_SL g4137 ( 
.A(n_4051),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_3965),
.B(n_155),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_4018),
.B(n_156),
.Y(n_4139)
);

OR2x2_ASAP7_75t_L g4140 ( 
.A(n_4009),
.B(n_157),
.Y(n_4140)
);

HB1xp67_ASAP7_75t_L g4141 ( 
.A(n_4033),
.Y(n_4141)
);

AOI22xp33_ASAP7_75t_L g4142 ( 
.A1(n_4041),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4028),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4045),
.Y(n_4144)
);

NAND2x1_ASAP7_75t_L g4145 ( 
.A(n_4034),
.B(n_160),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_4047),
.Y(n_4146)
);

INVx1_ASAP7_75t_SL g4147 ( 
.A(n_3988),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_4068),
.Y(n_4148)
);

INVx2_ASAP7_75t_L g4149 ( 
.A(n_4001),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_4014),
.B(n_159),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_4062),
.B(n_163),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_4046),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_4077),
.B(n_164),
.Y(n_4153)
);

INVxp67_ASAP7_75t_L g4154 ( 
.A(n_4016),
.Y(n_4154)
);

BUFx3_ASAP7_75t_L g4155 ( 
.A(n_3993),
.Y(n_4155)
);

INVxp67_ASAP7_75t_L g4156 ( 
.A(n_4023),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_4078),
.Y(n_4157)
);

OR2x2_ASAP7_75t_L g4158 ( 
.A(n_3982),
.B(n_164),
.Y(n_4158)
);

AND2x4_ASAP7_75t_L g4159 ( 
.A(n_4003),
.B(n_165),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_4029),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_4052),
.B(n_166),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_3980),
.B(n_166),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_4066),
.Y(n_4163)
);

INVx2_ASAP7_75t_SL g4164 ( 
.A(n_4059),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4067),
.Y(n_4165)
);

HB1xp67_ASAP7_75t_L g4166 ( 
.A(n_4017),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_3998),
.Y(n_4167)
);

AND2x2_ASAP7_75t_L g4168 ( 
.A(n_3986),
.B(n_167),
.Y(n_4168)
);

INVx2_ASAP7_75t_L g4169 ( 
.A(n_3987),
.Y(n_4169)
);

INVxp67_ASAP7_75t_SL g4170 ( 
.A(n_4069),
.Y(n_4170)
);

INVx4_ASAP7_75t_L g4171 ( 
.A(n_3989),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_3971),
.Y(n_4172)
);

AOI22xp33_ASAP7_75t_L g4173 ( 
.A1(n_4027),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_4173)
);

INVx2_ASAP7_75t_L g4174 ( 
.A(n_4054),
.Y(n_4174)
);

AND2x2_ASAP7_75t_L g4175 ( 
.A(n_4035),
.B(n_168),
.Y(n_4175)
);

HB1xp67_ASAP7_75t_L g4176 ( 
.A(n_4058),
.Y(n_4176)
);

OAI22xp5_ASAP7_75t_L g4177 ( 
.A1(n_4049),
.A2(n_4030),
.B1(n_4040),
.B2(n_4048),
.Y(n_4177)
);

AND2x2_ASAP7_75t_L g4178 ( 
.A(n_4007),
.B(n_4008),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4043),
.B(n_169),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_4073),
.B(n_170),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3991),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3997),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4011),
.Y(n_4183)
);

OR2x2_ASAP7_75t_L g4184 ( 
.A(n_4071),
.B(n_170),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3999),
.Y(n_4185)
);

AND2x2_ASAP7_75t_L g4186 ( 
.A(n_4012),
.B(n_171),
.Y(n_4186)
);

OR2x2_ASAP7_75t_L g4187 ( 
.A(n_3975),
.B(n_171),
.Y(n_4187)
);

INVx3_ASAP7_75t_L g4188 ( 
.A(n_3984),
.Y(n_4188)
);

AND2x2_ASAP7_75t_L g4189 ( 
.A(n_3992),
.B(n_172),
.Y(n_4189)
);

INVxp67_ASAP7_75t_SL g4190 ( 
.A(n_4013),
.Y(n_4190)
);

AND2x2_ASAP7_75t_L g4191 ( 
.A(n_4050),
.B(n_173),
.Y(n_4191)
);

AND2x2_ASAP7_75t_L g4192 ( 
.A(n_4000),
.B(n_174),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_3961),
.Y(n_4193)
);

HB1xp67_ASAP7_75t_L g4194 ( 
.A(n_3963),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_3967),
.B(n_174),
.Y(n_4195)
);

AND2x4_ASAP7_75t_L g4196 ( 
.A(n_3967),
.B(n_175),
.Y(n_4196)
);

OR2x2_ASAP7_75t_L g4197 ( 
.A(n_3964),
.B(n_176),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_3967),
.Y(n_4198)
);

AND2x2_ASAP7_75t_L g4199 ( 
.A(n_3967),
.B(n_177),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3961),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_3967),
.B(n_177),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_3994),
.B(n_178),
.Y(n_4202)
);

AND2x4_ASAP7_75t_SL g4203 ( 
.A(n_4026),
.B(n_178),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_3967),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_3967),
.B(n_179),
.Y(n_4205)
);

AOI22xp33_ASAP7_75t_L g4206 ( 
.A1(n_3966),
.A2(n_182),
.B1(n_179),
.B2(n_181),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_3967),
.B(n_181),
.Y(n_4207)
);

NAND2x1p5_ASAP7_75t_L g4208 ( 
.A(n_3967),
.B(n_183),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_3994),
.B(n_185),
.Y(n_4209)
);

BUFx6f_ASAP7_75t_L g4210 ( 
.A(n_3972),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3961),
.Y(n_4211)
);

BUFx2_ASAP7_75t_L g4212 ( 
.A(n_3967),
.Y(n_4212)
);

AND2x4_ASAP7_75t_L g4213 ( 
.A(n_3967),
.B(n_186),
.Y(n_4213)
);

AND2x2_ASAP7_75t_L g4214 ( 
.A(n_3967),
.B(n_187),
.Y(n_4214)
);

INVx2_ASAP7_75t_L g4215 ( 
.A(n_3967),
.Y(n_4215)
);

INVx5_ASAP7_75t_L g4216 ( 
.A(n_3972),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_3967),
.Y(n_4217)
);

NOR2xp33_ASAP7_75t_L g4218 ( 
.A(n_3974),
.B(n_187),
.Y(n_4218)
);

OR2x2_ASAP7_75t_L g4219 ( 
.A(n_3964),
.B(n_188),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_3961),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_3967),
.Y(n_4221)
);

INVxp67_ASAP7_75t_SL g4222 ( 
.A(n_3967),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_3967),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_3967),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3961),
.Y(n_4225)
);

OR2x2_ASAP7_75t_L g4226 ( 
.A(n_3964),
.B(n_188),
.Y(n_4226)
);

AND2x4_ASAP7_75t_L g4227 ( 
.A(n_3967),
.B(n_189),
.Y(n_4227)
);

AND2x2_ASAP7_75t_L g4228 ( 
.A(n_3967),
.B(n_190),
.Y(n_4228)
);

AND2x4_ASAP7_75t_L g4229 ( 
.A(n_3967),
.B(n_191),
.Y(n_4229)
);

INVx6_ASAP7_75t_L g4230 ( 
.A(n_4026),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_3961),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_3994),
.B(n_191),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_3994),
.B(n_192),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_3961),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_3967),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_3961),
.Y(n_4236)
);

AOI22xp33_ASAP7_75t_L g4237 ( 
.A1(n_3966),
.A2(n_195),
.B1(n_192),
.B2(n_194),
.Y(n_4237)
);

INVx2_ASAP7_75t_SL g4238 ( 
.A(n_4026),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_3994),
.B(n_194),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_4212),
.B(n_195),
.Y(n_4240)
);

OAI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_4084),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_4170),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4138),
.B(n_199),
.Y(n_4243)
);

OAI221xp5_ASAP7_75t_L g4244 ( 
.A1(n_4190),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.C(n_202),
.Y(n_4244)
);

NOR2xp33_ASAP7_75t_L g4245 ( 
.A(n_4171),
.B(n_200),
.Y(n_4245)
);

AOI22xp33_ASAP7_75t_L g4246 ( 
.A1(n_4136),
.A2(n_204),
.B1(n_201),
.B2(n_203),
.Y(n_4246)
);

AOI21xp33_ASAP7_75t_SL g4247 ( 
.A1(n_4166),
.A2(n_205),
.B(n_206),
.Y(n_4247)
);

OAI31xp33_ASAP7_75t_L g4248 ( 
.A1(n_4176),
.A2(n_209),
.A3(n_207),
.B(n_208),
.Y(n_4248)
);

NAND3xp33_ASAP7_75t_L g4249 ( 
.A(n_4141),
.B(n_207),
.C(n_210),
.Y(n_4249)
);

OAI221xp5_ASAP7_75t_L g4250 ( 
.A1(n_4165),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.C(n_214),
.Y(n_4250)
);

OAI22xp5_ASAP7_75t_L g4251 ( 
.A1(n_4091),
.A2(n_215),
.B1(n_212),
.B2(n_214),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4083),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4222),
.B(n_215),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4230),
.Y(n_4254)
);

OAI22xp5_ASAP7_75t_L g4255 ( 
.A1(n_4202),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_4255)
);

OAI22xp5_ASAP7_75t_L g4256 ( 
.A1(n_4209),
.A2(n_219),
.B1(n_216),
.B2(n_218),
.Y(n_4256)
);

AO21x1_ASAP7_75t_SL g4257 ( 
.A1(n_4232),
.A2(n_219),
.B(n_220),
.Y(n_4257)
);

NOR2xp33_ASAP7_75t_R g4258 ( 
.A(n_4182),
.B(n_220),
.Y(n_4258)
);

AND2x2_ASAP7_75t_L g4259 ( 
.A(n_4198),
.B(n_224),
.Y(n_4259)
);

AND2x4_ASAP7_75t_L g4260 ( 
.A(n_4216),
.B(n_224),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4093),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_4204),
.B(n_225),
.Y(n_4262)
);

AOI22xp33_ASAP7_75t_L g4263 ( 
.A1(n_4163),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_4263)
);

AND2x2_ASAP7_75t_L g4264 ( 
.A(n_4215),
.B(n_226),
.Y(n_4264)
);

INVx3_ASAP7_75t_L g4265 ( 
.A(n_4230),
.Y(n_4265)
);

AOI22xp33_ASAP7_75t_SL g4266 ( 
.A1(n_4109),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_4266)
);

OAI22xp5_ASAP7_75t_L g4267 ( 
.A1(n_4233),
.A2(n_4239),
.B1(n_4135),
.B2(n_4098),
.Y(n_4267)
);

AOI21xp5_ASAP7_75t_L g4268 ( 
.A1(n_4139),
.A2(n_230),
.B(n_231),
.Y(n_4268)
);

OR2x2_ASAP7_75t_L g4269 ( 
.A(n_4217),
.B(n_231),
.Y(n_4269)
);

INVx2_ASAP7_75t_R g4270 ( 
.A(n_4125),
.Y(n_4270)
);

OR2x2_ASAP7_75t_L g4271 ( 
.A(n_4221),
.B(n_4235),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4096),
.Y(n_4272)
);

OA21x2_ASAP7_75t_L g4273 ( 
.A1(n_4129),
.A2(n_4128),
.B(n_4126),
.Y(n_4273)
);

AOI211xp5_ASAP7_75t_L g4274 ( 
.A1(n_4177),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4101),
.Y(n_4275)
);

NOR2xp33_ASAP7_75t_R g4276 ( 
.A(n_4155),
.B(n_232),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_4216),
.Y(n_4277)
);

OAI211xp5_ASAP7_75t_L g4278 ( 
.A1(n_4161),
.A2(n_236),
.B(n_233),
.C(n_235),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_4223),
.B(n_235),
.Y(n_4279)
);

AND2x2_ASAP7_75t_L g4280 ( 
.A(n_4224),
.B(n_236),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_4210),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4103),
.Y(n_4282)
);

OR2x2_ASAP7_75t_L g4283 ( 
.A(n_4097),
.B(n_237),
.Y(n_4283)
);

HB1xp67_ASAP7_75t_L g4284 ( 
.A(n_4079),
.Y(n_4284)
);

OAI211xp5_ASAP7_75t_L g4285 ( 
.A1(n_4145),
.A2(n_239),
.B(n_237),
.C(n_238),
.Y(n_4285)
);

AOI22xp33_ASAP7_75t_L g4286 ( 
.A1(n_4183),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_4286)
);

INVx4_ASAP7_75t_L g4287 ( 
.A(n_4203),
.Y(n_4287)
);

AND2x2_ASAP7_75t_L g4288 ( 
.A(n_4090),
.B(n_241),
.Y(n_4288)
);

CKINVDCx5p33_ASAP7_75t_R g4289 ( 
.A(n_4238),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4112),
.Y(n_4290)
);

OA21x2_ASAP7_75t_L g4291 ( 
.A1(n_4137),
.A2(n_242),
.B(n_243),
.Y(n_4291)
);

BUFx10_ASAP7_75t_L g4292 ( 
.A(n_4196),
.Y(n_4292)
);

AND2x2_ASAP7_75t_L g4293 ( 
.A(n_4105),
.B(n_242),
.Y(n_4293)
);

A2O1A1Ixp33_ASAP7_75t_L g4294 ( 
.A1(n_4218),
.A2(n_246),
.B(n_244),
.C(n_245),
.Y(n_4294)
);

BUFx3_ASAP7_75t_L g4295 ( 
.A(n_4213),
.Y(n_4295)
);

OAI21x1_ASAP7_75t_L g4296 ( 
.A1(n_4099),
.A2(n_244),
.B(n_246),
.Y(n_4296)
);

OR2x2_ASAP7_75t_L g4297 ( 
.A(n_4095),
.B(n_247),
.Y(n_4297)
);

OAI22xp5_ASAP7_75t_L g4298 ( 
.A1(n_4152),
.A2(n_251),
.B1(n_248),
.B2(n_250),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4113),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4116),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4118),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4120),
.Y(n_4302)
);

NOR3xp33_ASAP7_75t_L g4303 ( 
.A(n_4151),
.B(n_250),
.C(n_251),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4124),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4193),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4200),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4211),
.Y(n_4307)
);

OAI22xp33_ASAP7_75t_L g4308 ( 
.A1(n_4174),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4210),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_4157),
.B(n_4143),
.Y(n_4310)
);

OR2x2_ASAP7_75t_L g4311 ( 
.A(n_4194),
.B(n_252),
.Y(n_4311)
);

NOR4xp25_ASAP7_75t_SL g4312 ( 
.A(n_4144),
.B(n_257),
.C(n_253),
.D(n_254),
.Y(n_4312)
);

OR2x2_ASAP7_75t_L g4313 ( 
.A(n_4087),
.B(n_257),
.Y(n_4313)
);

AOI22xp33_ASAP7_75t_SL g4314 ( 
.A1(n_4191),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_4314)
);

OAI22xp5_ASAP7_75t_L g4315 ( 
.A1(n_4154),
.A2(n_263),
.B1(n_260),
.B2(n_262),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_L g4316 ( 
.A(n_4146),
.B(n_262),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_4111),
.B(n_264),
.Y(n_4317)
);

OA21x2_ASAP7_75t_L g4318 ( 
.A1(n_4156),
.A2(n_264),
.B(n_265),
.Y(n_4318)
);

AOI22xp5_ASAP7_75t_L g4319 ( 
.A1(n_4164),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_4319)
);

BUFx2_ASAP7_75t_SL g4320 ( 
.A(n_4227),
.Y(n_4320)
);

HB1xp67_ASAP7_75t_L g4321 ( 
.A(n_4148),
.Y(n_4321)
);

NOR4xp25_ASAP7_75t_SL g4322 ( 
.A(n_4160),
.B(n_270),
.C(n_267),
.D(n_269),
.Y(n_4322)
);

CKINVDCx20_ASAP7_75t_R g4323 ( 
.A(n_4102),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4220),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4225),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_4181),
.B(n_269),
.Y(n_4326)
);

INVx2_ASAP7_75t_L g4327 ( 
.A(n_4111),
.Y(n_4327)
);

INVx2_ASAP7_75t_SL g4328 ( 
.A(n_4229),
.Y(n_4328)
);

OR2x2_ASAP7_75t_L g4329 ( 
.A(n_4197),
.B(n_270),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_4132),
.B(n_271),
.Y(n_4330)
);

INVx1_ASAP7_75t_SL g4331 ( 
.A(n_4080),
.Y(n_4331)
);

AO21x2_ASAP7_75t_L g4332 ( 
.A1(n_4195),
.A2(n_271),
.B(n_272),
.Y(n_4332)
);

NOR2xp33_ASAP7_75t_L g4333 ( 
.A(n_4147),
.B(n_272),
.Y(n_4333)
);

AOI31xp33_ASAP7_75t_L g4334 ( 
.A1(n_4208),
.A2(n_275),
.A3(n_273),
.B(n_274),
.Y(n_4334)
);

AOI221xp5_ASAP7_75t_L g4335 ( 
.A1(n_4179),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.C(n_277),
.Y(n_4335)
);

AND2x2_ASAP7_75t_L g4336 ( 
.A(n_4119),
.B(n_276),
.Y(n_4336)
);

NAND3xp33_ASAP7_75t_L g4337 ( 
.A(n_4142),
.B(n_277),
.C(n_278),
.Y(n_4337)
);

NOR2xp33_ASAP7_75t_R g4338 ( 
.A(n_4140),
.B(n_4158),
.Y(n_4338)
);

INVx3_ASAP7_75t_L g4339 ( 
.A(n_4106),
.Y(n_4339)
);

AOI22xp33_ASAP7_75t_L g4340 ( 
.A1(n_4172),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4231),
.Y(n_4341)
);

OR2x6_ASAP7_75t_L g4342 ( 
.A(n_4089),
.B(n_279),
.Y(n_4342)
);

BUFx2_ASAP7_75t_L g4343 ( 
.A(n_4199),
.Y(n_4343)
);

OAI31xp33_ASAP7_75t_L g4344 ( 
.A1(n_4153),
.A2(n_283),
.A3(n_280),
.B(n_281),
.Y(n_4344)
);

AOI22xp5_ASAP7_75t_L g4345 ( 
.A1(n_4173),
.A2(n_284),
.B1(n_281),
.B2(n_283),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4201),
.B(n_285),
.Y(n_4346)
);

OAI22xp5_ASAP7_75t_L g4347 ( 
.A1(n_4104),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_4347)
);

OAI211xp5_ASAP7_75t_L g4348 ( 
.A1(n_4180),
.A2(n_290),
.B(n_287),
.C(n_288),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_4186),
.A2(n_288),
.B(n_290),
.Y(n_4349)
);

OAI22xp5_ASAP7_75t_L g4350 ( 
.A1(n_4206),
.A2(n_295),
.B1(n_291),
.B2(n_293),
.Y(n_4350)
);

AND3x1_ASAP7_75t_L g4351 ( 
.A(n_4178),
.B(n_291),
.C(n_293),
.Y(n_4351)
);

OR2x2_ASAP7_75t_L g4352 ( 
.A(n_4219),
.B(n_4226),
.Y(n_4352)
);

NOR2x1_ASAP7_75t_SL g4353 ( 
.A(n_4205),
.B(n_4207),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4117),
.B(n_295),
.Y(n_4354)
);

OAI33xp33_ASAP7_75t_L g4355 ( 
.A1(n_4234),
.A2(n_4236),
.A3(n_4088),
.B1(n_4184),
.B2(n_4131),
.B3(n_4108),
.Y(n_4355)
);

OA21x2_ASAP7_75t_L g4356 ( 
.A1(n_4214),
.A2(n_296),
.B(n_297),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4092),
.Y(n_4357)
);

AOI221xp5_ASAP7_75t_L g4358 ( 
.A1(n_4188),
.A2(n_299),
.B1(n_296),
.B2(n_298),
.C(n_300),
.Y(n_4358)
);

AOI22xp33_ASAP7_75t_L g4359 ( 
.A1(n_4169),
.A2(n_301),
.B1(n_298),
.B2(n_300),
.Y(n_4359)
);

NAND3xp33_ASAP7_75t_L g4360 ( 
.A(n_4237),
.B(n_301),
.C(n_302),
.Y(n_4360)
);

INVxp67_ASAP7_75t_L g4361 ( 
.A(n_4228),
.Y(n_4361)
);

INVx3_ASAP7_75t_L g4362 ( 
.A(n_4082),
.Y(n_4362)
);

HB1xp67_ASAP7_75t_L g4363 ( 
.A(n_4085),
.Y(n_4363)
);

HB1xp67_ASAP7_75t_L g4364 ( 
.A(n_4127),
.Y(n_4364)
);

BUFx2_ASAP7_75t_L g4365 ( 
.A(n_4134),
.Y(n_4365)
);

AND2x2_ASAP7_75t_L g4366 ( 
.A(n_4081),
.B(n_303),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4094),
.Y(n_4367)
);

NOR2xp33_ASAP7_75t_R g4368 ( 
.A(n_4175),
.B(n_303),
.Y(n_4368)
);

AOI22xp33_ASAP7_75t_L g4369 ( 
.A1(n_4185),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_4369)
);

INVx2_ASAP7_75t_SL g4370 ( 
.A(n_4100),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4107),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_4086),
.B(n_304),
.Y(n_4372)
);

AOI22xp33_ASAP7_75t_L g4373 ( 
.A1(n_4150),
.A2(n_308),
.B1(n_305),
.B2(n_307),
.Y(n_4373)
);

AOI21xp5_ASAP7_75t_L g4374 ( 
.A1(n_4159),
.A2(n_309),
.B(n_310),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_4130),
.B(n_309),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4167),
.B(n_311),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4122),
.Y(n_4377)
);

OR2x2_ASAP7_75t_L g4378 ( 
.A(n_4149),
.B(n_311),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4110),
.Y(n_4379)
);

AOI221xp5_ASAP7_75t_L g4380 ( 
.A1(n_4115),
.A2(n_315),
.B1(n_312),
.B2(n_313),
.C(n_316),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4133),
.Y(n_4381)
);

OAI332xp33_ASAP7_75t_SL g4382 ( 
.A1(n_4123),
.A2(n_319),
.A3(n_318),
.B1(n_315),
.B2(n_320),
.B3(n_312),
.C1(n_313),
.C2(n_316),
.Y(n_4382)
);

OAI22xp33_ASAP7_75t_L g4383 ( 
.A1(n_4187),
.A2(n_322),
.B1(n_318),
.B2(n_319),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4121),
.Y(n_4384)
);

AO21x2_ASAP7_75t_L g4385 ( 
.A1(n_4114),
.A2(n_4192),
.B(n_4162),
.Y(n_4385)
);

CKINVDCx5p33_ASAP7_75t_R g4386 ( 
.A(n_4168),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4189),
.Y(n_4387)
);

OA21x2_ASAP7_75t_L g4388 ( 
.A1(n_4129),
.A2(n_323),
.B(n_324),
.Y(n_4388)
);

OR2x2_ASAP7_75t_L g4389 ( 
.A(n_4198),
.B(n_323),
.Y(n_4389)
);

OAI21xp5_ASAP7_75t_L g4390 ( 
.A1(n_4084),
.A2(n_324),
.B(n_325),
.Y(n_4390)
);

AND2x2_ASAP7_75t_L g4391 ( 
.A(n_4212),
.B(n_325),
.Y(n_4391)
);

OAI33xp33_ASAP7_75t_L g4392 ( 
.A1(n_4091),
.A2(n_328),
.A3(n_330),
.B1(n_326),
.B2(n_327),
.B3(n_329),
.Y(n_4392)
);

OAI221xp5_ASAP7_75t_L g4393 ( 
.A1(n_4170),
.A2(n_330),
.B1(n_327),
.B2(n_329),
.C(n_331),
.Y(n_4393)
);

OAI221xp5_ASAP7_75t_SL g4394 ( 
.A1(n_4170),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_4394)
);

INVx2_ASAP7_75t_SL g4395 ( 
.A(n_4230),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4212),
.B(n_334),
.Y(n_4396)
);

OAI332xp33_ASAP7_75t_L g4397 ( 
.A1(n_4170),
.A2(n_341),
.A3(n_340),
.B1(n_337),
.B2(n_343),
.B3(n_335),
.C1(n_336),
.C2(n_338),
.Y(n_4397)
);

OA21x2_ASAP7_75t_L g4398 ( 
.A1(n_4129),
.A2(n_336),
.B(n_338),
.Y(n_4398)
);

AOI22xp33_ASAP7_75t_L g4399 ( 
.A1(n_4170),
.A2(n_345),
.B1(n_341),
.B2(n_343),
.Y(n_4399)
);

INVx2_ASAP7_75t_L g4400 ( 
.A(n_4212),
.Y(n_4400)
);

BUFx3_ASAP7_75t_L g4401 ( 
.A(n_4230),
.Y(n_4401)
);

CKINVDCx16_ASAP7_75t_R g4402 ( 
.A(n_4084),
.Y(n_4402)
);

AOI22xp33_ASAP7_75t_L g4403 ( 
.A1(n_4170),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_4403)
);

AND2x2_ASAP7_75t_SL g4404 ( 
.A(n_4136),
.B(n_346),
.Y(n_4404)
);

OR2x2_ASAP7_75t_L g4405 ( 
.A(n_4198),
.B(n_348),
.Y(n_4405)
);

OAI22xp33_ASAP7_75t_L g4406 ( 
.A1(n_4098),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4083),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4083),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4083),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4083),
.Y(n_4410)
);

HB1xp67_ASAP7_75t_L g4411 ( 
.A(n_4212),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4083),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4083),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4212),
.B(n_350),
.Y(n_4414)
);

INVx2_ASAP7_75t_L g4415 ( 
.A(n_4212),
.Y(n_4415)
);

BUFx3_ASAP7_75t_L g4416 ( 
.A(n_4230),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4083),
.Y(n_4417)
);

AOI22xp33_ASAP7_75t_L g4418 ( 
.A1(n_4170),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_4418)
);

NOR2xp33_ASAP7_75t_L g4419 ( 
.A(n_4171),
.B(n_352),
.Y(n_4419)
);

NOR2x1p5_ASAP7_75t_L g4420 ( 
.A(n_4171),
.B(n_354),
.Y(n_4420)
);

HB1xp67_ASAP7_75t_L g4421 ( 
.A(n_4212),
.Y(n_4421)
);

INVx4_ASAP7_75t_L g4422 ( 
.A(n_4203),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4083),
.Y(n_4423)
);

OAI21xp33_ASAP7_75t_L g4424 ( 
.A1(n_4170),
.A2(n_355),
.B(n_356),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4083),
.Y(n_4425)
);

OA21x2_ASAP7_75t_L g4426 ( 
.A1(n_4129),
.A2(n_355),
.B(n_356),
.Y(n_4426)
);

BUFx3_ASAP7_75t_L g4427 ( 
.A(n_4230),
.Y(n_4427)
);

OAI221xp5_ASAP7_75t_L g4428 ( 
.A1(n_4170),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.C(n_360),
.Y(n_4428)
);

A2O1A1Ixp33_ASAP7_75t_L g4429 ( 
.A1(n_4084),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_4429)
);

BUFx3_ASAP7_75t_L g4430 ( 
.A(n_4230),
.Y(n_4430)
);

AOI221xp5_ASAP7_75t_L g4431 ( 
.A1(n_4170),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.C(n_363),
.Y(n_4431)
);

AND2x4_ASAP7_75t_L g4432 ( 
.A(n_4216),
.B(n_361),
.Y(n_4432)
);

AOI33xp33_ASAP7_75t_L g4433 ( 
.A1(n_4191),
.A2(n_364),
.A3(n_366),
.B1(n_362),
.B2(n_363),
.B3(n_365),
.Y(n_4433)
);

OR2x2_ASAP7_75t_L g4434 ( 
.A(n_4198),
.B(n_364),
.Y(n_4434)
);

NAND3xp33_ASAP7_75t_L g4435 ( 
.A(n_4402),
.B(n_366),
.C(n_367),
.Y(n_4435)
);

AOI22xp5_ASAP7_75t_SL g4436 ( 
.A1(n_4241),
.A2(n_369),
.B1(n_370),
.B2(n_368),
.Y(n_4436)
);

NAND2xp5_ASAP7_75t_SL g4437 ( 
.A(n_4265),
.B(n_367),
.Y(n_4437)
);

NAND3xp33_ASAP7_75t_L g4438 ( 
.A(n_4274),
.B(n_368),
.C(n_369),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4411),
.B(n_371),
.Y(n_4439)
);

AO21x2_ASAP7_75t_L g4440 ( 
.A1(n_4276),
.A2(n_371),
.B(n_372),
.Y(n_4440)
);

NAND4xp75_ASAP7_75t_L g4441 ( 
.A(n_4351),
.B(n_374),
.C(n_372),
.D(n_373),
.Y(n_4441)
);

AND2x2_ASAP7_75t_L g4442 ( 
.A(n_4401),
.B(n_375),
.Y(n_4442)
);

NOR3xp33_ASAP7_75t_L g4443 ( 
.A(n_4397),
.B(n_376),
.C(n_377),
.Y(n_4443)
);

OR2x2_ASAP7_75t_L g4444 ( 
.A(n_4364),
.B(n_376),
.Y(n_4444)
);

AO22x1_ASAP7_75t_L g4445 ( 
.A1(n_4390),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4416),
.B(n_378),
.Y(n_4446)
);

AND2x2_ASAP7_75t_L g4447 ( 
.A(n_4427),
.B(n_379),
.Y(n_4447)
);

XOR2x2_ASAP7_75t_L g4448 ( 
.A(n_4394),
.B(n_380),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_4430),
.B(n_380),
.Y(n_4449)
);

AOI22xp33_ASAP7_75t_SL g4450 ( 
.A1(n_4353),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_4450)
);

NOR2x1_ASAP7_75t_L g4451 ( 
.A(n_4388),
.B(n_4398),
.Y(n_4451)
);

AND2x2_ASAP7_75t_L g4452 ( 
.A(n_4395),
.B(n_381),
.Y(n_4452)
);

AO21x2_ASAP7_75t_L g4453 ( 
.A1(n_4277),
.A2(n_382),
.B(n_384),
.Y(n_4453)
);

NOR3xp33_ASAP7_75t_L g4454 ( 
.A(n_4267),
.B(n_384),
.C(n_385),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4284),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_L g4456 ( 
.A(n_4421),
.B(n_386),
.Y(n_4456)
);

NAND4xp75_ASAP7_75t_L g4457 ( 
.A(n_4273),
.B(n_388),
.C(n_386),
.D(n_387),
.Y(n_4457)
);

OR2x2_ASAP7_75t_L g4458 ( 
.A(n_4400),
.B(n_387),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4343),
.B(n_388),
.Y(n_4459)
);

NOR3xp33_ASAP7_75t_L g4460 ( 
.A(n_4278),
.B(n_389),
.C(n_390),
.Y(n_4460)
);

AOI211xp5_ASAP7_75t_L g4461 ( 
.A1(n_4429),
.A2(n_394),
.B(n_392),
.C(n_393),
.Y(n_4461)
);

NAND3xp33_ASAP7_75t_L g4462 ( 
.A(n_4431),
.B(n_392),
.C(n_393),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4273),
.Y(n_4463)
);

INVx2_ASAP7_75t_SL g4464 ( 
.A(n_4292),
.Y(n_4464)
);

BUFx2_ASAP7_75t_L g4465 ( 
.A(n_4323),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4331),
.B(n_4415),
.Y(n_4466)
);

NOR3xp33_ASAP7_75t_L g4467 ( 
.A(n_4355),
.B(n_394),
.C(n_396),
.Y(n_4467)
);

BUFx2_ASAP7_75t_L g4468 ( 
.A(n_4363),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_4252),
.Y(n_4469)
);

AOI22xp33_ASAP7_75t_L g4470 ( 
.A1(n_4303),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_4470)
);

NAND3xp33_ASAP7_75t_L g4471 ( 
.A(n_4358),
.B(n_397),
.C(n_398),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4365),
.B(n_399),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_L g4473 ( 
.A(n_4404),
.B(n_400),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4261),
.Y(n_4474)
);

OR2x2_ASAP7_75t_L g4475 ( 
.A(n_4352),
.B(n_4310),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_4370),
.B(n_400),
.Y(n_4476)
);

OR2x2_ASAP7_75t_L g4477 ( 
.A(n_4271),
.B(n_401),
.Y(n_4477)
);

NOR2xp33_ASAP7_75t_L g4478 ( 
.A(n_4287),
.B(n_402),
.Y(n_4478)
);

AND2x4_ASAP7_75t_L g4479 ( 
.A(n_4254),
.B(n_403),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4385),
.B(n_404),
.Y(n_4480)
);

NAND3xp33_ASAP7_75t_L g4481 ( 
.A(n_4248),
.B(n_404),
.C(n_405),
.Y(n_4481)
);

INVx2_ASAP7_75t_L g4482 ( 
.A(n_4295),
.Y(n_4482)
);

NAND2x1_ASAP7_75t_L g4483 ( 
.A(n_4339),
.B(n_405),
.Y(n_4483)
);

NOR2xp33_ASAP7_75t_L g4484 ( 
.A(n_4422),
.B(n_406),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_4377),
.B(n_407),
.Y(n_4485)
);

NOR2xp33_ASAP7_75t_L g4486 ( 
.A(n_4289),
.B(n_409),
.Y(n_4486)
);

NAND3xp33_ASAP7_75t_L g4487 ( 
.A(n_4335),
.B(n_410),
.C(n_411),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_SL g4488 ( 
.A(n_4362),
.B(n_410),
.Y(n_4488)
);

NOR3xp33_ASAP7_75t_L g4489 ( 
.A(n_4251),
.B(n_411),
.C(n_412),
.Y(n_4489)
);

AOI211xp5_ASAP7_75t_L g4490 ( 
.A1(n_4406),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_4490)
);

NAND3xp33_ASAP7_75t_L g4491 ( 
.A(n_4380),
.B(n_413),
.C(n_414),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4379),
.B(n_415),
.Y(n_4492)
);

AOI22xp33_ASAP7_75t_SL g4493 ( 
.A1(n_4338),
.A2(n_418),
.B1(n_416),
.B2(n_417),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4327),
.B(n_416),
.Y(n_4494)
);

NAND4xp25_ASAP7_75t_L g4495 ( 
.A(n_4314),
.B(n_419),
.C(n_417),
.D(n_418),
.Y(n_4495)
);

AOI22xp33_ASAP7_75t_L g4496 ( 
.A1(n_4270),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_4496)
);

AND2x4_ASAP7_75t_L g4497 ( 
.A(n_4281),
.B(n_420),
.Y(n_4497)
);

NOR3xp33_ASAP7_75t_L g4498 ( 
.A(n_4255),
.B(n_423),
.C(n_425),
.Y(n_4498)
);

NAND3xp33_ASAP7_75t_L g4499 ( 
.A(n_4249),
.B(n_423),
.C(n_425),
.Y(n_4499)
);

INVx2_ASAP7_75t_L g4500 ( 
.A(n_4260),
.Y(n_4500)
);

AOI22xp5_ASAP7_75t_L g4501 ( 
.A1(n_4256),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_4501)
);

OR2x2_ASAP7_75t_L g4502 ( 
.A(n_4361),
.B(n_426),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_L g4503 ( 
.A(n_4357),
.B(n_427),
.Y(n_4503)
);

AO21x2_ASAP7_75t_L g4504 ( 
.A1(n_4316),
.A2(n_428),
.B(n_429),
.Y(n_4504)
);

OAI211xp5_ASAP7_75t_L g4505 ( 
.A1(n_4247),
.A2(n_437),
.B(n_447),
.C(n_429),
.Y(n_4505)
);

AND2x2_ASAP7_75t_L g4506 ( 
.A(n_4309),
.B(n_430),
.Y(n_4506)
);

OR2x2_ASAP7_75t_L g4507 ( 
.A(n_4367),
.B(n_431),
.Y(n_4507)
);

NOR3xp33_ASAP7_75t_L g4508 ( 
.A(n_4393),
.B(n_431),
.C(n_432),
.Y(n_4508)
);

OR2x2_ASAP7_75t_L g4509 ( 
.A(n_4371),
.B(n_433),
.Y(n_4509)
);

BUFx2_ASAP7_75t_L g4510 ( 
.A(n_4432),
.Y(n_4510)
);

NOR2xp33_ASAP7_75t_L g4511 ( 
.A(n_4424),
.B(n_433),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_4387),
.B(n_434),
.Y(n_4512)
);

INVx2_ASAP7_75t_SL g4513 ( 
.A(n_4328),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4381),
.B(n_434),
.Y(n_4514)
);

NAND4xp75_ASAP7_75t_L g4515 ( 
.A(n_4291),
.B(n_438),
.C(n_435),
.D(n_436),
.Y(n_4515)
);

OR2x2_ASAP7_75t_L g4516 ( 
.A(n_4283),
.B(n_435),
.Y(n_4516)
);

INVx2_ASAP7_75t_L g4517 ( 
.A(n_4384),
.Y(n_4517)
);

OAI21xp5_ASAP7_75t_L g4518 ( 
.A1(n_4294),
.A2(n_438),
.B(n_439),
.Y(n_4518)
);

INVxp33_ASAP7_75t_SL g4519 ( 
.A(n_4368),
.Y(n_4519)
);

AND2x2_ASAP7_75t_L g4520 ( 
.A(n_4320),
.B(n_4336),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4272),
.Y(n_4521)
);

OAI211xp5_ASAP7_75t_L g4522 ( 
.A1(n_4348),
.A2(n_450),
.B(n_459),
.C(n_439),
.Y(n_4522)
);

NAND3xp33_ASAP7_75t_L g4523 ( 
.A(n_4433),
.B(n_441),
.C(n_442),
.Y(n_4523)
);

OAI211xp5_ASAP7_75t_L g4524 ( 
.A1(n_4285),
.A2(n_453),
.B(n_461),
.C(n_442),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_4268),
.B(n_444),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4275),
.Y(n_4526)
);

INVxp67_ASAP7_75t_L g4527 ( 
.A(n_4257),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_4297),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4282),
.Y(n_4529)
);

OR2x2_ASAP7_75t_L g4530 ( 
.A(n_4269),
.B(n_444),
.Y(n_4530)
);

AND2x4_ASAP7_75t_L g4531 ( 
.A(n_4321),
.B(n_445),
.Y(n_4531)
);

AOI22xp5_ASAP7_75t_L g4532 ( 
.A1(n_4245),
.A2(n_448),
.B1(n_445),
.B2(n_446),
.Y(n_4532)
);

BUFx3_ASAP7_75t_L g4533 ( 
.A(n_4288),
.Y(n_4533)
);

NAND3xp33_ASAP7_75t_L g4534 ( 
.A(n_4344),
.B(n_449),
.C(n_450),
.Y(n_4534)
);

BUFx2_ASAP7_75t_L g4535 ( 
.A(n_4342),
.Y(n_4535)
);

NAND4xp75_ASAP7_75t_L g4536 ( 
.A(n_4291),
.B(n_4398),
.C(n_4426),
.D(n_4388),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_4356),
.B(n_449),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_4313),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4356),
.B(n_451),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4290),
.Y(n_4540)
);

NAND3xp33_ASAP7_75t_L g4541 ( 
.A(n_4419),
.B(n_451),
.C(n_454),
.Y(n_4541)
);

AOI22xp5_ASAP7_75t_L g4542 ( 
.A1(n_4392),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_4542)
);

NOR3xp33_ASAP7_75t_L g4543 ( 
.A(n_4428),
.B(n_455),
.C(n_457),
.Y(n_4543)
);

AO21x2_ASAP7_75t_L g4544 ( 
.A1(n_4258),
.A2(n_4253),
.B(n_4243),
.Y(n_4544)
);

NAND3xp33_ASAP7_75t_L g4545 ( 
.A(n_4266),
.B(n_458),
.C(n_459),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4376),
.B(n_458),
.Y(n_4546)
);

NOR3xp33_ASAP7_75t_L g4547 ( 
.A(n_4349),
.B(n_460),
.C(n_461),
.Y(n_4547)
);

NOR3xp33_ASAP7_75t_L g4548 ( 
.A(n_4244),
.B(n_4250),
.C(n_4337),
.Y(n_4548)
);

OR2x2_ASAP7_75t_L g4549 ( 
.A(n_4434),
.B(n_460),
.Y(n_4549)
);

NOR3xp33_ASAP7_75t_L g4550 ( 
.A(n_4360),
.B(n_462),
.C(n_464),
.Y(n_4550)
);

OR2x2_ASAP7_75t_L g4551 ( 
.A(n_4389),
.B(n_466),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_4240),
.B(n_467),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4391),
.B(n_467),
.Y(n_4553)
);

NAND3xp33_ASAP7_75t_L g4554 ( 
.A(n_4242),
.B(n_468),
.C(n_469),
.Y(n_4554)
);

OAI211xp5_ASAP7_75t_SL g4555 ( 
.A1(n_4399),
.A2(n_471),
.B(n_468),
.C(n_469),
.Y(n_4555)
);

NOR2xp33_ASAP7_75t_L g4556 ( 
.A(n_4378),
.B(n_471),
.Y(n_4556)
);

NAND2xp5_ASAP7_75t_L g4557 ( 
.A(n_4318),
.B(n_472),
.Y(n_4557)
);

INVx1_ASAP7_75t_SL g4558 ( 
.A(n_4396),
.Y(n_4558)
);

NAND3xp33_ASAP7_75t_L g4559 ( 
.A(n_4403),
.B(n_473),
.C(n_474),
.Y(n_4559)
);

AND2x2_ASAP7_75t_L g4560 ( 
.A(n_4414),
.B(n_473),
.Y(n_4560)
);

OR2x2_ASAP7_75t_L g4561 ( 
.A(n_4405),
.B(n_4326),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_4318),
.B(n_4332),
.Y(n_4562)
);

OA21x2_ASAP7_75t_L g4563 ( 
.A1(n_4299),
.A2(n_474),
.B(n_475),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_4386),
.B(n_475),
.Y(n_4564)
);

INVxp67_ASAP7_75t_SL g4565 ( 
.A(n_4420),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4319),
.B(n_476),
.Y(n_4566)
);

AND2x2_ASAP7_75t_L g4567 ( 
.A(n_4293),
.B(n_476),
.Y(n_4567)
);

OA211x2_ASAP7_75t_L g4568 ( 
.A1(n_4317),
.A2(n_479),
.B(n_477),
.C(n_478),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_4259),
.B(n_477),
.Y(n_4569)
);

NAND3xp33_ASAP7_75t_L g4570 ( 
.A(n_4418),
.B(n_478),
.C(n_479),
.Y(n_4570)
);

AND2x2_ASAP7_75t_L g4571 ( 
.A(n_4262),
.B(n_482),
.Y(n_4571)
);

AOI33xp33_ASAP7_75t_L g4572 ( 
.A1(n_4450),
.A2(n_4246),
.A3(n_4308),
.B1(n_4373),
.B2(n_4263),
.B3(n_4383),
.Y(n_4572)
);

OR2x2_ASAP7_75t_L g4573 ( 
.A(n_4558),
.B(n_4466),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4465),
.Y(n_4574)
);

AOI33xp33_ASAP7_75t_L g4575 ( 
.A1(n_4493),
.A2(n_4369),
.A3(n_4340),
.B1(n_4286),
.B2(n_4359),
.B3(n_4322),
.Y(n_4575)
);

OR2x2_ASAP7_75t_L g4576 ( 
.A(n_4468),
.B(n_4330),
.Y(n_4576)
);

AND2x2_ASAP7_75t_L g4577 ( 
.A(n_4520),
.B(n_4264),
.Y(n_4577)
);

NAND4xp25_ASAP7_75t_L g4578 ( 
.A(n_4443),
.B(n_4345),
.C(n_4333),
.D(n_4374),
.Y(n_4578)
);

OAI211xp5_ASAP7_75t_L g4579 ( 
.A1(n_4467),
.A2(n_4312),
.B(n_4426),
.C(n_4315),
.Y(n_4579)
);

HB1xp67_ASAP7_75t_L g4580 ( 
.A(n_4510),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4565),
.B(n_4535),
.Y(n_4581)
);

NOR2xp33_ASAP7_75t_L g4582 ( 
.A(n_4519),
.B(n_4354),
.Y(n_4582)
);

OAI31xp33_ASAP7_75t_L g4583 ( 
.A1(n_4438),
.A2(n_4298),
.A3(n_4350),
.B(n_4347),
.Y(n_4583)
);

AOI22xp33_ASAP7_75t_L g4584 ( 
.A1(n_4548),
.A2(n_4464),
.B1(n_4543),
.B2(n_4508),
.Y(n_4584)
);

OR2x2_ASAP7_75t_L g4585 ( 
.A(n_4562),
.B(n_4311),
.Y(n_4585)
);

INVx2_ASAP7_75t_L g4586 ( 
.A(n_4533),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4483),
.Y(n_4587)
);

OAI221xp5_ASAP7_75t_L g4588 ( 
.A1(n_4451),
.A2(n_4334),
.B1(n_4342),
.B2(n_4300),
.C(n_4304),
.Y(n_4588)
);

AOI322xp5_ASAP7_75t_L g4589 ( 
.A1(n_4460),
.A2(n_4375),
.A3(n_4346),
.B1(n_4372),
.B2(n_4280),
.C1(n_4279),
.C2(n_4302),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4463),
.Y(n_4590)
);

AND2x2_ASAP7_75t_L g4591 ( 
.A(n_4500),
.B(n_4366),
.Y(n_4591)
);

AOI22xp33_ASAP7_75t_L g4592 ( 
.A1(n_4454),
.A2(n_4301),
.B1(n_4306),
.B2(n_4305),
.Y(n_4592)
);

OR2x2_ASAP7_75t_L g4593 ( 
.A(n_4475),
.B(n_4307),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4513),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4482),
.B(n_4324),
.Y(n_4595)
);

INVx4_ASAP7_75t_L g4596 ( 
.A(n_4479),
.Y(n_4596)
);

BUFx2_ASAP7_75t_L g4597 ( 
.A(n_4544),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4455),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_4527),
.B(n_4325),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_4497),
.Y(n_4600)
);

INVx1_ASAP7_75t_SL g4601 ( 
.A(n_4459),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_SL g4602 ( 
.A(n_4542),
.B(n_4531),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4507),
.Y(n_4603)
);

INVx2_ASAP7_75t_L g4604 ( 
.A(n_4497),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_4440),
.B(n_4341),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4509),
.Y(n_4606)
);

OAI33xp33_ASAP7_75t_L g4607 ( 
.A1(n_4480),
.A2(n_4407),
.A3(n_4409),
.B1(n_4412),
.B2(n_4410),
.B3(n_4408),
.Y(n_4607)
);

INVx2_ASAP7_75t_SL g4608 ( 
.A(n_4479),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_4517),
.B(n_4413),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4504),
.B(n_4528),
.Y(n_4610)
);

BUFx3_ASAP7_75t_L g4611 ( 
.A(n_4442),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4538),
.B(n_4417),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4444),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_4556),
.B(n_4423),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4502),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4531),
.Y(n_4616)
);

INVx2_ASAP7_75t_L g4617 ( 
.A(n_4458),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4476),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_4453),
.B(n_4425),
.Y(n_4619)
);

NAND3xp33_ASAP7_75t_L g4620 ( 
.A(n_4462),
.B(n_4329),
.C(n_4382),
.Y(n_4620)
);

AND2x2_ASAP7_75t_L g4621 ( 
.A(n_4478),
.B(n_4484),
.Y(n_4621)
);

AND2x4_ASAP7_75t_L g4622 ( 
.A(n_4452),
.B(n_4296),
.Y(n_4622)
);

NOR2xp33_ASAP7_75t_L g4623 ( 
.A(n_4561),
.B(n_482),
.Y(n_4623)
);

AND2x2_ASAP7_75t_L g4624 ( 
.A(n_4546),
.B(n_483),
.Y(n_4624)
);

OAI21xp5_ASAP7_75t_L g4625 ( 
.A1(n_4536),
.A2(n_487),
.B(n_488),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4446),
.B(n_488),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4469),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4447),
.B(n_489),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4474),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4441),
.B(n_490),
.Y(n_4630)
);

HB1xp67_ASAP7_75t_L g4631 ( 
.A(n_4563),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4521),
.Y(n_4632)
);

NAND4xp25_ASAP7_75t_L g4633 ( 
.A(n_4523),
.B(n_494),
.C(n_491),
.D(n_493),
.Y(n_4633)
);

HB1xp67_ASAP7_75t_L g4634 ( 
.A(n_4563),
.Y(n_4634)
);

INVx2_ASAP7_75t_SL g4635 ( 
.A(n_4449),
.Y(n_4635)
);

OAI31xp33_ASAP7_75t_L g4636 ( 
.A1(n_4522),
.A2(n_4524),
.A3(n_4491),
.B(n_4487),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4526),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_4477),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4529),
.Y(n_4639)
);

AOI21xp33_ASAP7_75t_L g4640 ( 
.A1(n_4525),
.A2(n_491),
.B(n_494),
.Y(n_4640)
);

NOR3xp33_ASAP7_75t_SL g4641 ( 
.A(n_4471),
.B(n_495),
.C(n_496),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_4494),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4567),
.B(n_496),
.Y(n_4643)
);

OAI221xp5_ASAP7_75t_L g4644 ( 
.A1(n_4489),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.C(n_501),
.Y(n_4644)
);

AOI22xp33_ASAP7_75t_L g4645 ( 
.A1(n_4547),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4537),
.B(n_501),
.Y(n_4646)
);

NOR3xp33_ASAP7_75t_L g4647 ( 
.A(n_4481),
.B(n_502),
.C(n_503),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4540),
.Y(n_4648)
);

BUFx2_ASAP7_75t_L g4649 ( 
.A(n_4439),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4472),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4506),
.Y(n_4651)
);

AOI33xp33_ASAP7_75t_L g4652 ( 
.A1(n_4470),
.A2(n_505),
.A3(n_507),
.B1(n_503),
.B2(n_504),
.B3(n_506),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4456),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_4530),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4516),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4552),
.B(n_4553),
.Y(n_4656)
);

OR2x2_ASAP7_75t_L g4657 ( 
.A(n_4512),
.B(n_504),
.Y(n_4657)
);

NAND2x1p5_ASAP7_75t_L g4658 ( 
.A(n_4488),
.B(n_506),
.Y(n_4658)
);

OAI31xp33_ASAP7_75t_L g4659 ( 
.A1(n_4505),
.A2(n_508),
.A3(n_505),
.B(n_507),
.Y(n_4659)
);

AOI22xp33_ASAP7_75t_L g4660 ( 
.A1(n_4498),
.A2(n_511),
.B1(n_509),
.B2(n_510),
.Y(n_4660)
);

INVx3_ASAP7_75t_L g4661 ( 
.A(n_4549),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4503),
.Y(n_4662)
);

NAND4xp25_ASAP7_75t_L g4663 ( 
.A(n_4461),
.B(n_512),
.C(n_510),
.D(n_511),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_4551),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4580),
.Y(n_4665)
);

INVx3_ASAP7_75t_L g4666 ( 
.A(n_4596),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_4590),
.Y(n_4667)
);

INVx2_ASAP7_75t_SL g4668 ( 
.A(n_4608),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4631),
.Y(n_4669)
);

AOI22xp5_ASAP7_75t_L g4670 ( 
.A1(n_4579),
.A2(n_4550),
.B1(n_4457),
.B2(n_4534),
.Y(n_4670)
);

INVxp67_ASAP7_75t_SL g4671 ( 
.A(n_4658),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_4634),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4581),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4661),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4597),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4655),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4574),
.B(n_4539),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_4601),
.B(n_4557),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4577),
.B(n_4560),
.Y(n_4679)
);

INVxp67_ASAP7_75t_L g4680 ( 
.A(n_4587),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_4656),
.B(n_4600),
.Y(n_4681)
);

NAND2x1_ASAP7_75t_SL g4682 ( 
.A(n_4622),
.B(n_4569),
.Y(n_4682)
);

NOR2xp33_ASAP7_75t_L g4683 ( 
.A(n_4611),
.B(n_4485),
.Y(n_4683)
);

AOI22xp5_ASAP7_75t_L g4684 ( 
.A1(n_4625),
.A2(n_4545),
.B1(n_4448),
.B2(n_4515),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_4604),
.Y(n_4685)
);

INVx1_ASAP7_75t_SL g4686 ( 
.A(n_4573),
.Y(n_4686)
);

NAND4xp75_ASAP7_75t_SL g4687 ( 
.A(n_4636),
.B(n_4511),
.C(n_4486),
.D(n_4571),
.Y(n_4687)
);

A2O1A1Ixp33_ASAP7_75t_L g4688 ( 
.A1(n_4659),
.A2(n_4436),
.B(n_4435),
.C(n_4518),
.Y(n_4688)
);

INVx3_ASAP7_75t_L g4689 ( 
.A(n_4616),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4664),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_4594),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_L g4692 ( 
.A(n_4635),
.B(n_4492),
.Y(n_4692)
);

NOR2xp33_ASAP7_75t_SL g4693 ( 
.A(n_4588),
.B(n_4495),
.Y(n_4693)
);

INVx2_ASAP7_75t_L g4694 ( 
.A(n_4591),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4654),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4638),
.Y(n_4696)
);

INVx2_ASAP7_75t_L g4697 ( 
.A(n_4586),
.Y(n_4697)
);

AND2x4_ASAP7_75t_L g4698 ( 
.A(n_4642),
.B(n_4514),
.Y(n_4698)
);

INVx4_ASAP7_75t_L g4699 ( 
.A(n_4626),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_4622),
.B(n_4564),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4603),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4606),
.Y(n_4702)
);

AOI22xp33_ASAP7_75t_L g4703 ( 
.A1(n_4584),
.A2(n_4555),
.B1(n_4559),
.B2(n_4554),
.Y(n_4703)
);

OAI22xp5_ASAP7_75t_L g4704 ( 
.A1(n_4641),
.A2(n_4496),
.B1(n_4501),
.B2(n_4499),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4617),
.Y(n_4705)
);

AND2x2_ASAP7_75t_L g4706 ( 
.A(n_4651),
.B(n_4437),
.Y(n_4706)
);

AOI22xp5_ASAP7_75t_L g4707 ( 
.A1(n_4578),
.A2(n_4647),
.B1(n_4602),
.B2(n_4633),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4615),
.Y(n_4708)
);

AND2x2_ASAP7_75t_L g4709 ( 
.A(n_4621),
.B(n_4473),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4613),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4612),
.Y(n_4711)
);

AND2x2_ASAP7_75t_L g4712 ( 
.A(n_4649),
.B(n_4532),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4599),
.Y(n_4713)
);

AND2x4_ASAP7_75t_L g4714 ( 
.A(n_4595),
.B(n_4541),
.Y(n_4714)
);

INVx1_ASAP7_75t_SL g4715 ( 
.A(n_4576),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4593),
.Y(n_4716)
);

AND2x2_ASAP7_75t_L g4717 ( 
.A(n_4582),
.B(n_4566),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4598),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4624),
.Y(n_4719)
);

INVx2_ASAP7_75t_L g4720 ( 
.A(n_4643),
.Y(n_4720)
);

INVxp33_ASAP7_75t_L g4721 ( 
.A(n_4623),
.Y(n_4721)
);

INVx2_ASAP7_75t_SL g4722 ( 
.A(n_4609),
.Y(n_4722)
);

OA222x2_ASAP7_75t_L g4723 ( 
.A1(n_4605),
.A2(n_4568),
.B1(n_4445),
.B2(n_4490),
.C1(n_4570),
.C2(n_514),
.Y(n_4723)
);

INVx2_ASAP7_75t_SL g4724 ( 
.A(n_4628),
.Y(n_4724)
);

AOI22xp5_ASAP7_75t_L g4725 ( 
.A1(n_4663),
.A2(n_516),
.B1(n_512),
.B2(n_513),
.Y(n_4725)
);

INVx2_ASAP7_75t_SL g4726 ( 
.A(n_4682),
.Y(n_4726)
);

AND2x4_ASAP7_75t_L g4727 ( 
.A(n_4668),
.B(n_4666),
.Y(n_4727)
);

OAI33xp33_ASAP7_75t_L g4728 ( 
.A1(n_4669),
.A2(n_4672),
.A3(n_4675),
.B1(n_4610),
.B2(n_4665),
.B3(n_4673),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4681),
.Y(n_4729)
);

AND2x2_ASAP7_75t_L g4730 ( 
.A(n_4679),
.B(n_4650),
.Y(n_4730)
);

INVxp67_ASAP7_75t_L g4731 ( 
.A(n_4693),
.Y(n_4731)
);

AND2x2_ASAP7_75t_L g4732 ( 
.A(n_4700),
.B(n_4589),
.Y(n_4732)
);

INVxp67_ASAP7_75t_L g4733 ( 
.A(n_4671),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4689),
.B(n_4653),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_L g4735 ( 
.A(n_4684),
.B(n_4583),
.Y(n_4735)
);

OR2x2_ASAP7_75t_L g4736 ( 
.A(n_4686),
.B(n_4585),
.Y(n_4736)
);

NAND2xp5_ASAP7_75t_L g4737 ( 
.A(n_4699),
.B(n_4618),
.Y(n_4737)
);

OAI211xp5_ASAP7_75t_L g4738 ( 
.A1(n_4670),
.A2(n_4660),
.B(n_4645),
.C(n_4619),
.Y(n_4738)
);

NOR2xp67_ASAP7_75t_SL g4739 ( 
.A(n_4697),
.B(n_4657),
.Y(n_4739)
);

OR2x2_ASAP7_75t_L g4740 ( 
.A(n_4724),
.B(n_4694),
.Y(n_4740)
);

AND2x2_ASAP7_75t_L g4741 ( 
.A(n_4706),
.B(n_4662),
.Y(n_4741)
);

OR2x2_ASAP7_75t_L g4742 ( 
.A(n_4715),
.B(n_4614),
.Y(n_4742)
);

NAND2xp5_ASAP7_75t_L g4743 ( 
.A(n_4680),
.B(n_4592),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4709),
.B(n_4627),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4685),
.Y(n_4745)
);

OR2x2_ASAP7_75t_L g4746 ( 
.A(n_4674),
.B(n_4620),
.Y(n_4746)
);

OR2x2_ASAP7_75t_SL g4747 ( 
.A(n_4716),
.B(n_4630),
.Y(n_4747)
);

BUFx2_ASAP7_75t_L g4748 ( 
.A(n_4722),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4719),
.Y(n_4749)
);

OR2x2_ASAP7_75t_L g4750 ( 
.A(n_4720),
.B(n_4646),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_4711),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4695),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4714),
.B(n_4629),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_4688),
.B(n_4572),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4696),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4691),
.B(n_4632),
.Y(n_4756)
);

OR2x2_ASAP7_75t_L g4757 ( 
.A(n_4678),
.B(n_4637),
.Y(n_4757)
);

INVx3_ASAP7_75t_L g4758 ( 
.A(n_4698),
.Y(n_4758)
);

AND2x2_ASAP7_75t_L g4759 ( 
.A(n_4712),
.B(n_4639),
.Y(n_4759)
);

AND2x2_ASAP7_75t_L g4760 ( 
.A(n_4683),
.B(n_4648),
.Y(n_4760)
);

INVx3_ASAP7_75t_L g4761 ( 
.A(n_4705),
.Y(n_4761)
);

OR2x4_ASAP7_75t_L g4762 ( 
.A(n_4677),
.B(n_4607),
.Y(n_4762)
);

AND2x2_ASAP7_75t_L g4763 ( 
.A(n_4717),
.B(n_4640),
.Y(n_4763)
);

OR2x2_ASAP7_75t_L g4764 ( 
.A(n_4692),
.B(n_4644),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4676),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4713),
.B(n_4721),
.Y(n_4766)
);

AND2x4_ASAP7_75t_L g4767 ( 
.A(n_4701),
.B(n_4575),
.Y(n_4767)
);

AND2x2_ASAP7_75t_L g4768 ( 
.A(n_4723),
.B(n_4652),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4690),
.Y(n_4769)
);

INVxp67_ASAP7_75t_L g4770 ( 
.A(n_4702),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4710),
.B(n_513),
.Y(n_4771)
);

AND2x2_ASAP7_75t_L g4772 ( 
.A(n_4708),
.B(n_517),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4727),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4758),
.B(n_4707),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4732),
.B(n_4703),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4748),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_L g4777 ( 
.A(n_4726),
.B(n_4704),
.Y(n_4777)
);

INVx1_ASAP7_75t_SL g4778 ( 
.A(n_4736),
.Y(n_4778)
);

OAI31xp33_ASAP7_75t_L g4779 ( 
.A1(n_4738),
.A2(n_4718),
.A3(n_4667),
.B(n_4687),
.Y(n_4779)
);

NAND2xp5_ASAP7_75t_L g4780 ( 
.A(n_4768),
.B(n_4725),
.Y(n_4780)
);

HB1xp67_ASAP7_75t_L g4781 ( 
.A(n_4740),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4730),
.Y(n_4782)
);

INVx2_ASAP7_75t_L g4783 ( 
.A(n_4734),
.Y(n_4783)
);

NAND3xp33_ASAP7_75t_L g4784 ( 
.A(n_4754),
.B(n_517),
.C(n_518),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4759),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4753),
.B(n_518),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4744),
.B(n_519),
.Y(n_4787)
);

AND2x2_ASAP7_75t_L g4788 ( 
.A(n_4741),
.B(n_519),
.Y(n_4788)
);

OR2x2_ASAP7_75t_L g4789 ( 
.A(n_4747),
.B(n_520),
.Y(n_4789)
);

AOI22xp5_ASAP7_75t_L g4790 ( 
.A1(n_4731),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.Y(n_4790)
);

AND2x2_ASAP7_75t_L g4791 ( 
.A(n_4733),
.B(n_521),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4771),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4772),
.Y(n_4793)
);

AND2x2_ASAP7_75t_L g4794 ( 
.A(n_4760),
.B(n_523),
.Y(n_4794)
);

AND2x2_ASAP7_75t_L g4795 ( 
.A(n_4766),
.B(n_4763),
.Y(n_4795)
);

NAND3xp33_ASAP7_75t_L g4796 ( 
.A(n_4735),
.B(n_523),
.C(n_524),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4739),
.B(n_525),
.Y(n_4797)
);

NOR3xp33_ASAP7_75t_SL g4798 ( 
.A(n_4728),
.B(n_525),
.C(n_526),
.Y(n_4798)
);

NAND4xp25_ASAP7_75t_L g4799 ( 
.A(n_4746),
.B(n_528),
.C(n_526),
.D(n_527),
.Y(n_4799)
);

NAND3xp33_ASAP7_75t_L g4800 ( 
.A(n_4767),
.B(n_527),
.C(n_528),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4761),
.B(n_529),
.Y(n_4801)
);

AOI22xp33_ASAP7_75t_L g4802 ( 
.A1(n_4743),
.A2(n_4729),
.B1(n_4764),
.B2(n_4742),
.Y(n_4802)
);

OR2x2_ASAP7_75t_L g4803 ( 
.A(n_4737),
.B(n_529),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4745),
.B(n_530),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4756),
.Y(n_4805)
);

INVxp67_ASAP7_75t_L g4806 ( 
.A(n_4750),
.Y(n_4806)
);

XNOR2x2_ASAP7_75t_L g4807 ( 
.A(n_4757),
.B(n_530),
.Y(n_4807)
);

AND2x2_ASAP7_75t_L g4808 ( 
.A(n_4749),
.B(n_4751),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4752),
.B(n_4755),
.Y(n_4809)
);

NOR2xp67_ASAP7_75t_SL g4810 ( 
.A(n_4765),
.B(n_531),
.Y(n_4810)
);

INVx1_ASAP7_75t_SL g4811 ( 
.A(n_4769),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_SL g4812 ( 
.A(n_4770),
.B(n_532),
.Y(n_4812)
);

OAI22xp33_ASAP7_75t_L g4813 ( 
.A1(n_4762),
.A2(n_535),
.B1(n_533),
.B2(n_534),
.Y(n_4813)
);

AOI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4731),
.A2(n_537),
.B1(n_533),
.B2(n_536),
.Y(n_4814)
);

AOI211x1_ASAP7_75t_L g4815 ( 
.A1(n_4738),
.A2(n_538),
.B(n_536),
.C(n_537),
.Y(n_4815)
);

OR2x2_ASAP7_75t_L g4816 ( 
.A(n_4747),
.B(n_539),
.Y(n_4816)
);

NOR3xp33_ASAP7_75t_SL g4817 ( 
.A(n_4728),
.B(n_539),
.C(n_540),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_SL g4818 ( 
.A(n_4727),
.B(n_540),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_L g4819 ( 
.A(n_4727),
.B(n_541),
.Y(n_4819)
);

NOR2xp33_ASAP7_75t_L g4820 ( 
.A(n_4731),
.B(n_542),
.Y(n_4820)
);

NOR2xp33_ASAP7_75t_L g4821 ( 
.A(n_4731),
.B(n_542),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4781),
.Y(n_4822)
);

NOR2x1_ASAP7_75t_L g4823 ( 
.A(n_4799),
.B(n_543),
.Y(n_4823)
);

AOI221xp5_ASAP7_75t_L g4824 ( 
.A1(n_4813),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.C(n_546),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_L g4825 ( 
.A(n_4773),
.B(n_544),
.Y(n_4825)
);

NOR2x1_ASAP7_75t_L g4826 ( 
.A(n_4800),
.B(n_545),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4776),
.Y(n_4827)
);

OR2x2_ASAP7_75t_L g4828 ( 
.A(n_4778),
.B(n_547),
.Y(n_4828)
);

OAI311xp33_ASAP7_75t_L g4829 ( 
.A1(n_4775),
.A2(n_549),
.A3(n_547),
.B1(n_548),
.C1(n_550),
.Y(n_4829)
);

INVx1_ASAP7_75t_SL g4830 ( 
.A(n_4789),
.Y(n_4830)
);

AND2x2_ASAP7_75t_L g4831 ( 
.A(n_4795),
.B(n_551),
.Y(n_4831)
);

AND2x4_ASAP7_75t_L g4832 ( 
.A(n_4786),
.B(n_4783),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4788),
.Y(n_4833)
);

AND2x2_ASAP7_75t_L g4834 ( 
.A(n_4782),
.B(n_552),
.Y(n_4834)
);

OAI221xp5_ASAP7_75t_SL g4835 ( 
.A1(n_4779),
.A2(n_554),
.B1(n_552),
.B2(n_553),
.C(n_555),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_SL g4836 ( 
.A(n_4798),
.B(n_553),
.Y(n_4836)
);

AND2x2_ASAP7_75t_L g4837 ( 
.A(n_4774),
.B(n_556),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4787),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4819),
.Y(n_4839)
);

AND2x2_ASAP7_75t_L g4840 ( 
.A(n_4785),
.B(n_556),
.Y(n_4840)
);

AND2x4_ASAP7_75t_L g4841 ( 
.A(n_4805),
.B(n_557),
.Y(n_4841)
);

OAI221xp5_ASAP7_75t_L g4842 ( 
.A1(n_4817),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.C(n_560),
.Y(n_4842)
);

AND2x2_ASAP7_75t_L g4843 ( 
.A(n_4794),
.B(n_559),
.Y(n_4843)
);

AOI31xp33_ASAP7_75t_L g4844 ( 
.A1(n_4802),
.A2(n_4806),
.A3(n_4777),
.B(n_4780),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4791),
.Y(n_4845)
);

NAND2xp5_ASAP7_75t_L g4846 ( 
.A(n_4815),
.B(n_560),
.Y(n_4846)
);

OAI21xp5_ASAP7_75t_L g4847 ( 
.A1(n_4796),
.A2(n_561),
.B(n_562),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4816),
.Y(n_4848)
);

NOR2xp33_ASAP7_75t_L g4849 ( 
.A(n_4818),
.B(n_562),
.Y(n_4849)
);

INVx1_ASAP7_75t_SL g4850 ( 
.A(n_4807),
.Y(n_4850)
);

OAI32xp33_ASAP7_75t_L g4851 ( 
.A1(n_4811),
.A2(n_565),
.A3(n_567),
.B1(n_564),
.B2(n_566),
.Y(n_4851)
);

NAND2xp5_ASAP7_75t_L g4852 ( 
.A(n_4810),
.B(n_563),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4792),
.B(n_564),
.Y(n_4853)
);

AOI31xp33_ASAP7_75t_L g4854 ( 
.A1(n_4793),
.A2(n_568),
.A3(n_566),
.B(n_567),
.Y(n_4854)
);

AND2x4_ASAP7_75t_SL g4855 ( 
.A(n_4808),
.B(n_569),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4797),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4803),
.Y(n_4857)
);

NAND4xp25_ASAP7_75t_SL g4858 ( 
.A(n_4784),
.B(n_572),
.C(n_570),
.D(n_571),
.Y(n_4858)
);

OAI222xp33_ASAP7_75t_L g4859 ( 
.A1(n_4809),
.A2(n_573),
.B1(n_577),
.B2(n_570),
.C1(n_571),
.C2(n_576),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4801),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4820),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4821),
.Y(n_4862)
);

OAI21xp33_ASAP7_75t_L g4863 ( 
.A1(n_4804),
.A2(n_573),
.B(n_577),
.Y(n_4863)
);

OAI21xp5_ASAP7_75t_SL g4864 ( 
.A1(n_4790),
.A2(n_579),
.B(n_580),
.Y(n_4864)
);

OAI21xp33_ASAP7_75t_L g4865 ( 
.A1(n_4814),
.A2(n_579),
.B(n_580),
.Y(n_4865)
);

OAI21xp5_ASAP7_75t_L g4866 ( 
.A1(n_4812),
.A2(n_581),
.B(n_583),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4773),
.B(n_584),
.Y(n_4867)
);

XOR2xp5_ASAP7_75t_L g4868 ( 
.A(n_4773),
.B(n_584),
.Y(n_4868)
);

AOI221x1_ASAP7_75t_SL g4869 ( 
.A1(n_4813),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.C(n_588),
.Y(n_4869)
);

AND2x4_ASAP7_75t_L g4870 ( 
.A(n_4781),
.B(n_587),
.Y(n_4870)
);

OAI22xp33_ASAP7_75t_SL g4871 ( 
.A1(n_4775),
.A2(n_591),
.B1(n_589),
.B2(n_590),
.Y(n_4871)
);

AOI221x1_ASAP7_75t_L g4872 ( 
.A1(n_4776),
.A2(n_593),
.B1(n_589),
.B2(n_592),
.C(n_594),
.Y(n_4872)
);

AOI21xp33_ASAP7_75t_SL g4873 ( 
.A1(n_4813),
.A2(n_597),
.B(n_596),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4781),
.Y(n_4874)
);

OAI21xp5_ASAP7_75t_L g4875 ( 
.A1(n_4813),
.A2(n_592),
.B(n_597),
.Y(n_4875)
);

CKINVDCx16_ASAP7_75t_R g4876 ( 
.A(n_4781),
.Y(n_4876)
);

NOR4xp25_ASAP7_75t_L g4877 ( 
.A(n_4813),
.B(n_600),
.C(n_598),
.D(n_599),
.Y(n_4877)
);

AND2x2_ASAP7_75t_L g4878 ( 
.A(n_4773),
.B(n_598),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4781),
.Y(n_4879)
);

AOI321xp33_ASAP7_75t_L g4880 ( 
.A1(n_4835),
.A2(n_601),
.A3(n_603),
.B1(n_599),
.B2(n_600),
.C(n_602),
.Y(n_4880)
);

NOR2xp33_ASAP7_75t_L g4881 ( 
.A(n_4876),
.B(n_601),
.Y(n_4881)
);

OAI21xp33_ASAP7_75t_L g4882 ( 
.A1(n_4844),
.A2(n_610),
.B(n_602),
.Y(n_4882)
);

AND2x2_ASAP7_75t_L g4883 ( 
.A(n_4837),
.B(n_603),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_L g4884 ( 
.A(n_4850),
.B(n_604),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_L g4885 ( 
.A(n_4832),
.B(n_604),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4832),
.B(n_605),
.Y(n_4886)
);

NOR2xp33_ASAP7_75t_L g4887 ( 
.A(n_4842),
.B(n_606),
.Y(n_4887)
);

NOR2xp33_ASAP7_75t_L g4888 ( 
.A(n_4836),
.B(n_606),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4868),
.Y(n_4889)
);

INVxp67_ASAP7_75t_L g4890 ( 
.A(n_4831),
.Y(n_4890)
);

AND2x2_ASAP7_75t_L g4891 ( 
.A(n_4878),
.B(n_607),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4855),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_4870),
.B(n_607),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4870),
.B(n_608),
.Y(n_4894)
);

NOR2xp33_ASAP7_75t_SL g4895 ( 
.A(n_4822),
.B(n_608),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_L g4896 ( 
.A(n_4869),
.B(n_609),
.Y(n_4896)
);

INVxp67_ASAP7_75t_SL g4897 ( 
.A(n_4874),
.Y(n_4897)
);

AO22x2_ASAP7_75t_L g4898 ( 
.A1(n_4872),
.A2(n_612),
.B1(n_610),
.B2(n_611),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4879),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4828),
.Y(n_4900)
);

OAI21xp5_ASAP7_75t_L g4901 ( 
.A1(n_4823),
.A2(n_612),
.B(n_613),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4843),
.Y(n_4902)
);

NAND2xp5_ASAP7_75t_L g4903 ( 
.A(n_4877),
.B(n_615),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4834),
.Y(n_4904)
);

O2A1O1Ixp33_ASAP7_75t_L g4905 ( 
.A1(n_4829),
.A2(n_624),
.B(n_633),
.C(n_615),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4840),
.Y(n_4906)
);

NOR2xp33_ASAP7_75t_L g4907 ( 
.A(n_4830),
.B(n_616),
.Y(n_4907)
);

XOR2xp5_ASAP7_75t_L g4908 ( 
.A(n_4833),
.B(n_616),
.Y(n_4908)
);

INVx1_ASAP7_75t_L g4909 ( 
.A(n_4852),
.Y(n_4909)
);

AND2x4_ASAP7_75t_L g4910 ( 
.A(n_4838),
.B(n_617),
.Y(n_4910)
);

AND2x4_ASAP7_75t_L g4911 ( 
.A(n_4827),
.B(n_617),
.Y(n_4911)
);

INVxp33_ASAP7_75t_L g4912 ( 
.A(n_4826),
.Y(n_4912)
);

NAND2xp5_ASAP7_75t_L g4913 ( 
.A(n_4848),
.B(n_618),
.Y(n_4913)
);

AND2x2_ASAP7_75t_L g4914 ( 
.A(n_4845),
.B(n_619),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4841),
.Y(n_4915)
);

OAI33xp33_ASAP7_75t_L g4916 ( 
.A1(n_4856),
.A2(n_622),
.A3(n_624),
.B1(n_619),
.B2(n_621),
.B3(n_623),
.Y(n_4916)
);

INVx2_ASAP7_75t_L g4917 ( 
.A(n_4857),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_L g4918 ( 
.A(n_4873),
.B(n_621),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4825),
.Y(n_4919)
);

OR2x2_ASAP7_75t_L g4920 ( 
.A(n_4846),
.B(n_622),
.Y(n_4920)
);

INVx2_ASAP7_75t_L g4921 ( 
.A(n_4839),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4867),
.Y(n_4922)
);

AND2x2_ASAP7_75t_L g4923 ( 
.A(n_4875),
.B(n_625),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4849),
.B(n_626),
.Y(n_4924)
);

AND2x2_ASAP7_75t_L g4925 ( 
.A(n_4847),
.B(n_627),
.Y(n_4925)
);

OAI22xp5_ASAP7_75t_L g4926 ( 
.A1(n_4861),
.A2(n_629),
.B1(n_627),
.B2(n_628),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4854),
.Y(n_4927)
);

BUFx2_ASAP7_75t_L g4928 ( 
.A(n_4866),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4853),
.Y(n_4929)
);

NAND2x1p5_ASAP7_75t_L g4930 ( 
.A(n_4862),
.B(n_629),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4871),
.B(n_631),
.Y(n_4931)
);

AOI221xp5_ASAP7_75t_L g4932 ( 
.A1(n_4851),
.A2(n_634),
.B1(n_637),
.B2(n_632),
.C(n_635),
.Y(n_4932)
);

XNOR2x2_ASAP7_75t_L g4933 ( 
.A(n_4824),
.B(n_631),
.Y(n_4933)
);

AND2x2_ASAP7_75t_L g4934 ( 
.A(n_4860),
.B(n_632),
.Y(n_4934)
);

OR2x2_ASAP7_75t_L g4935 ( 
.A(n_4858),
.B(n_635),
.Y(n_4935)
);

NAND3xp33_ASAP7_75t_SL g4936 ( 
.A(n_4864),
.B(n_4865),
.C(n_4863),
.Y(n_4936)
);

HB1xp67_ASAP7_75t_L g4937 ( 
.A(n_4859),
.Y(n_4937)
);

HB1xp67_ASAP7_75t_L g4938 ( 
.A(n_4876),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4876),
.Y(n_4939)
);

AND2x2_ASAP7_75t_L g4940 ( 
.A(n_4876),
.B(n_637),
.Y(n_4940)
);

AOI21xp5_ASAP7_75t_L g4941 ( 
.A1(n_4836),
.A2(n_638),
.B(n_639),
.Y(n_4941)
);

OAI22xp5_ASAP7_75t_L g4942 ( 
.A1(n_4876),
.A2(n_641),
.B1(n_639),
.B2(n_640),
.Y(n_4942)
);

AND2x2_ASAP7_75t_L g4943 ( 
.A(n_4876),
.B(n_640),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4876),
.B(n_641),
.Y(n_4944)
);

AOI221xp5_ASAP7_75t_L g4945 ( 
.A1(n_4835),
.A2(n_644),
.B1(n_646),
.B2(n_643),
.C(n_645),
.Y(n_4945)
);

AND2x2_ASAP7_75t_L g4946 ( 
.A(n_4876),
.B(n_642),
.Y(n_4946)
);

INVx2_ASAP7_75t_L g4947 ( 
.A(n_4876),
.Y(n_4947)
);

AOI21xp33_ASAP7_75t_L g4948 ( 
.A1(n_4850),
.A2(n_646),
.B(n_644),
.Y(n_4948)
);

NOR2xp33_ASAP7_75t_L g4949 ( 
.A(n_4876),
.B(n_642),
.Y(n_4949)
);

NAND3xp33_ASAP7_75t_L g4950 ( 
.A(n_4835),
.B(n_647),
.C(n_648),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_4876),
.B(n_648),
.Y(n_4951)
);

NOR2xp33_ASAP7_75t_L g4952 ( 
.A(n_4876),
.B(n_649),
.Y(n_4952)
);

INVx1_ASAP7_75t_L g4953 ( 
.A(n_4876),
.Y(n_4953)
);

OAI22xp33_ASAP7_75t_L g4954 ( 
.A1(n_4876),
.A2(n_651),
.B1(n_649),
.B2(n_650),
.Y(n_4954)
);

OR2x2_ASAP7_75t_L g4955 ( 
.A(n_4876),
.B(n_651),
.Y(n_4955)
);

OAI211xp5_ASAP7_75t_L g4956 ( 
.A1(n_4850),
.A2(n_654),
.B(n_652),
.C(n_653),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4876),
.Y(n_4957)
);

INVx2_ASAP7_75t_L g4958 ( 
.A(n_4876),
.Y(n_4958)
);

OR2x2_ASAP7_75t_L g4959 ( 
.A(n_4876),
.B(n_653),
.Y(n_4959)
);

AND2x2_ASAP7_75t_L g4960 ( 
.A(n_4876),
.B(n_655),
.Y(n_4960)
);

XOR2x2_ASAP7_75t_L g4961 ( 
.A(n_4836),
.B(n_655),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4876),
.Y(n_4962)
);

BUFx6f_ASAP7_75t_L g4963 ( 
.A(n_4870),
.Y(n_4963)
);

NAND2xp5_ASAP7_75t_L g4964 ( 
.A(n_4876),
.B(n_657),
.Y(n_4964)
);

O2A1O1Ixp5_ASAP7_75t_L g4965 ( 
.A1(n_4835),
.A2(n_659),
.B(n_657),
.C(n_658),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4876),
.Y(n_4966)
);

NAND3xp33_ASAP7_75t_L g4967 ( 
.A(n_4835),
.B(n_658),
.C(n_660),
.Y(n_4967)
);

AND2x2_ASAP7_75t_L g4968 ( 
.A(n_4876),
.B(n_660),
.Y(n_4968)
);

INVx1_ASAP7_75t_SL g4969 ( 
.A(n_4876),
.Y(n_4969)
);

INVx1_ASAP7_75t_SL g4970 ( 
.A(n_4876),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4876),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4938),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_4969),
.B(n_661),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4940),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4943),
.Y(n_4975)
);

NAND2xp5_ASAP7_75t_L g4976 ( 
.A(n_4970),
.B(n_662),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4946),
.B(n_662),
.Y(n_4977)
);

INVx1_ASAP7_75t_L g4978 ( 
.A(n_4960),
.Y(n_4978)
);

NOR2x1_ASAP7_75t_L g4979 ( 
.A(n_4939),
.B(n_663),
.Y(n_4979)
);

AOI22xp5_ASAP7_75t_L g4980 ( 
.A1(n_4953),
.A2(n_665),
.B1(n_663),
.B2(n_664),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_L g4981 ( 
.A(n_4968),
.B(n_665),
.Y(n_4981)
);

INVx5_ASAP7_75t_L g4982 ( 
.A(n_4963),
.Y(n_4982)
);

AO21x1_ASAP7_75t_L g4983 ( 
.A1(n_4881),
.A2(n_4952),
.B(n_4949),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_SL g4984 ( 
.A(n_4963),
.B(n_666),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4955),
.Y(n_4985)
);

XNOR2xp5_ASAP7_75t_L g4986 ( 
.A(n_4961),
.B(n_4908),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_SL g4987 ( 
.A(n_4947),
.B(n_667),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4957),
.B(n_668),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4962),
.B(n_668),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4966),
.B(n_4971),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4959),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4958),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4944),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_4951),
.Y(n_4994)
);

INVxp33_ASAP7_75t_SL g4995 ( 
.A(n_4937),
.Y(n_4995)
);

AND2x2_ASAP7_75t_L g4996 ( 
.A(n_4927),
.B(n_4892),
.Y(n_4996)
);

OAI21xp5_ASAP7_75t_L g4997 ( 
.A1(n_4965),
.A2(n_669),
.B(n_670),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4964),
.Y(n_4998)
);

OR2x2_ASAP7_75t_L g4999 ( 
.A(n_4884),
.B(n_670),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4885),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4886),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4883),
.Y(n_5002)
);

AND2x2_ASAP7_75t_L g5003 ( 
.A(n_4915),
.B(n_671),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4902),
.B(n_671),
.Y(n_5004)
);

AND2x2_ASAP7_75t_L g5005 ( 
.A(n_4890),
.B(n_672),
.Y(n_5005)
);

AND2x2_ASAP7_75t_L g5006 ( 
.A(n_4904),
.B(n_672),
.Y(n_5006)
);

INVx2_ASAP7_75t_L g5007 ( 
.A(n_4930),
.Y(n_5007)
);

NAND2xp5_ASAP7_75t_L g5008 ( 
.A(n_4898),
.B(n_673),
.Y(n_5008)
);

NOR3xp33_ASAP7_75t_SL g5009 ( 
.A(n_4882),
.B(n_673),
.C(n_674),
.Y(n_5009)
);

OR2x2_ASAP7_75t_L g5010 ( 
.A(n_4903),
.B(n_4896),
.Y(n_5010)
);

INVx2_ASAP7_75t_L g5011 ( 
.A(n_4891),
.Y(n_5011)
);

INVx2_ASAP7_75t_L g5012 ( 
.A(n_4910),
.Y(n_5012)
);

CKINVDCx5p33_ASAP7_75t_R g5013 ( 
.A(n_4889),
.Y(n_5013)
);

NAND4xp25_ASAP7_75t_SL g5014 ( 
.A(n_4905),
.B(n_677),
.C(n_675),
.D(n_676),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_L g5015 ( 
.A(n_4898),
.B(n_678),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4897),
.B(n_678),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4935),
.Y(n_5017)
);

AOI22xp5_ASAP7_75t_L g5018 ( 
.A1(n_4887),
.A2(n_681),
.B1(n_679),
.B2(n_680),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4893),
.Y(n_5019)
);

INVx1_ASAP7_75t_L g5020 ( 
.A(n_4894),
.Y(n_5020)
);

AND4x1_ASAP7_75t_L g5021 ( 
.A(n_4895),
.B(n_4888),
.C(n_4907),
.D(n_4901),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4914),
.Y(n_5022)
);

INVxp67_ASAP7_75t_SL g5023 ( 
.A(n_4931),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4911),
.Y(n_5024)
);

AND2x2_ASAP7_75t_L g5025 ( 
.A(n_4906),
.B(n_681),
.Y(n_5025)
);

NAND2xp5_ASAP7_75t_L g5026 ( 
.A(n_4954),
.B(n_683),
.Y(n_5026)
);

AOI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_4941),
.A2(n_683),
.B(n_684),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4918),
.Y(n_5028)
);

OR2x2_ASAP7_75t_L g5029 ( 
.A(n_4920),
.B(n_684),
.Y(n_5029)
);

NOR3xp33_ASAP7_75t_SL g5030 ( 
.A(n_4936),
.B(n_685),
.C(n_686),
.Y(n_5030)
);

NAND2xp33_ASAP7_75t_SL g5031 ( 
.A(n_4912),
.B(n_687),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_SL g5032 ( 
.A(n_4880),
.B(n_687),
.Y(n_5032)
);

INVx2_ASAP7_75t_SL g5033 ( 
.A(n_4917),
.Y(n_5033)
);

INVx1_ASAP7_75t_L g5034 ( 
.A(n_4923),
.Y(n_5034)
);

AOI21xp5_ASAP7_75t_L g5035 ( 
.A1(n_4913),
.A2(n_689),
.B(n_690),
.Y(n_5035)
);

NOR2xp33_ASAP7_75t_R g5036 ( 
.A(n_4900),
.B(n_689),
.Y(n_5036)
);

NOR2xp33_ASAP7_75t_R g5037 ( 
.A(n_4899),
.B(n_691),
.Y(n_5037)
);

INVxp67_ASAP7_75t_L g5038 ( 
.A(n_4925),
.Y(n_5038)
);

HB1xp67_ASAP7_75t_L g5039 ( 
.A(n_4942),
.Y(n_5039)
);

OR2x2_ASAP7_75t_L g5040 ( 
.A(n_4950),
.B(n_691),
.Y(n_5040)
);

INVxp67_ASAP7_75t_L g5041 ( 
.A(n_4928),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_4945),
.B(n_692),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_4934),
.Y(n_5043)
);

INVxp67_ASAP7_75t_L g5044 ( 
.A(n_4916),
.Y(n_5044)
);

NAND2x1_ASAP7_75t_L g5045 ( 
.A(n_4921),
.B(n_692),
.Y(n_5045)
);

AND2x2_ASAP7_75t_L g5046 ( 
.A(n_4909),
.B(n_693),
.Y(n_5046)
);

INVx1_ASAP7_75t_SL g5047 ( 
.A(n_4933),
.Y(n_5047)
);

NAND3xp33_ASAP7_75t_L g5048 ( 
.A(n_4956),
.B(n_693),
.C(n_694),
.Y(n_5048)
);

AND2x2_ASAP7_75t_SL g5049 ( 
.A(n_4932),
.B(n_694),
.Y(n_5049)
);

OAI221xp5_ASAP7_75t_SL g5050 ( 
.A1(n_4919),
.A2(n_698),
.B1(n_696),
.B2(n_697),
.C(n_699),
.Y(n_5050)
);

NOR2x1_ASAP7_75t_L g5051 ( 
.A(n_4967),
.B(n_696),
.Y(n_5051)
);

AND2x2_ASAP7_75t_L g5052 ( 
.A(n_4922),
.B(n_4948),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4924),
.Y(n_5053)
);

INVx2_ASAP7_75t_L g5054 ( 
.A(n_4929),
.Y(n_5054)
);

NOR3xp33_ASAP7_75t_SL g5055 ( 
.A(n_4926),
.B(n_697),
.C(n_698),
.Y(n_5055)
);

INVx1_ASAP7_75t_SL g5056 ( 
.A(n_4969),
.Y(n_5056)
);

AOI21xp5_ASAP7_75t_L g5057 ( 
.A1(n_4938),
.A2(n_699),
.B(n_701),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4938),
.Y(n_5058)
);

NAND2xp33_ASAP7_75t_L g5059 ( 
.A(n_4938),
.B(n_701),
.Y(n_5059)
);

INVxp33_ASAP7_75t_L g5060 ( 
.A(n_4938),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4938),
.Y(n_5061)
);

AOI21xp5_ASAP7_75t_L g5062 ( 
.A1(n_5060),
.A2(n_702),
.B(n_703),
.Y(n_5062)
);

NOR3xp33_ASAP7_75t_L g5063 ( 
.A(n_4990),
.B(n_705),
.C(n_704),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_4982),
.B(n_703),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4982),
.Y(n_5065)
);

AO22x1_ASAP7_75t_L g5066 ( 
.A1(n_4982),
.A2(n_706),
.B1(n_704),
.B2(n_705),
.Y(n_5066)
);

AOI21xp5_ASAP7_75t_L g5067 ( 
.A1(n_5059),
.A2(n_706),
.B(n_709),
.Y(n_5067)
);

AOI22xp5_ASAP7_75t_L g5068 ( 
.A1(n_4995),
.A2(n_5056),
.B1(n_5058),
.B2(n_4972),
.Y(n_5068)
);

NOR2x1_ASAP7_75t_L g5069 ( 
.A(n_4979),
.B(n_709),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_5061),
.B(n_5047),
.Y(n_5070)
);

AND2x2_ASAP7_75t_L g5071 ( 
.A(n_4996),
.B(n_710),
.Y(n_5071)
);

NOR3x1_ASAP7_75t_L g5072 ( 
.A(n_5048),
.B(n_710),
.C(n_711),
.Y(n_5072)
);

NAND2xp5_ASAP7_75t_L g5073 ( 
.A(n_5003),
.B(n_712),
.Y(n_5073)
);

AOI211xp5_ASAP7_75t_L g5074 ( 
.A1(n_5014),
.A2(n_716),
.B(n_712),
.C(n_714),
.Y(n_5074)
);

OAI21xp5_ASAP7_75t_L g5075 ( 
.A1(n_5041),
.A2(n_718),
.B(n_717),
.Y(n_5075)
);

OAI21xp33_ASAP7_75t_L g5076 ( 
.A1(n_4992),
.A2(n_716),
.B(n_717),
.Y(n_5076)
);

OAI211xp5_ASAP7_75t_SL g5077 ( 
.A1(n_5044),
.A2(n_720),
.B(n_718),
.C(n_719),
.Y(n_5077)
);

AOI21xp5_ASAP7_75t_L g5078 ( 
.A1(n_5031),
.A2(n_719),
.B(n_721),
.Y(n_5078)
);

AOI21xp5_ASAP7_75t_L g5079 ( 
.A1(n_5032),
.A2(n_4987),
.B(n_5008),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_5004),
.B(n_721),
.Y(n_5080)
);

NAND2xp5_ASAP7_75t_L g5081 ( 
.A(n_4974),
.B(n_722),
.Y(n_5081)
);

NAND3xp33_ASAP7_75t_L g5082 ( 
.A(n_5030),
.B(n_722),
.C(n_723),
.Y(n_5082)
);

AO22x1_ASAP7_75t_L g5083 ( 
.A1(n_4997),
.A2(n_5051),
.B1(n_5015),
.B2(n_5007),
.Y(n_5083)
);

AOI22xp5_ASAP7_75t_L g5084 ( 
.A1(n_5013),
.A2(n_725),
.B1(n_723),
.B2(n_724),
.Y(n_5084)
);

NAND3xp33_ASAP7_75t_L g5085 ( 
.A(n_5055),
.B(n_724),
.C(n_726),
.Y(n_5085)
);

AOI21xp5_ASAP7_75t_L g5086 ( 
.A1(n_4973),
.A2(n_726),
.B(n_727),
.Y(n_5086)
);

AO22x2_ASAP7_75t_L g5087 ( 
.A1(n_4975),
.A2(n_729),
.B1(n_727),
.B2(n_728),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_5045),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_4976),
.Y(n_5089)
);

AOI221xp5_ASAP7_75t_L g5090 ( 
.A1(n_5033),
.A2(n_730),
.B1(n_728),
.B2(n_729),
.C(n_731),
.Y(n_5090)
);

AOI21xp5_ASAP7_75t_L g5091 ( 
.A1(n_4984),
.A2(n_731),
.B(n_732),
.Y(n_5091)
);

AOI211xp5_ASAP7_75t_L g5092 ( 
.A1(n_4983),
.A2(n_734),
.B(n_732),
.C(n_733),
.Y(n_5092)
);

AOI22xp5_ASAP7_75t_L g5093 ( 
.A1(n_4978),
.A2(n_736),
.B1(n_734),
.B2(n_735),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_4977),
.Y(n_5094)
);

INVx1_ASAP7_75t_L g5095 ( 
.A(n_4981),
.Y(n_5095)
);

NOR3x1_ASAP7_75t_L g5096 ( 
.A(n_5042),
.B(n_737),
.C(n_738),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_5006),
.Y(n_5097)
);

INVx1_ASAP7_75t_L g5098 ( 
.A(n_5025),
.Y(n_5098)
);

AOI31xp33_ASAP7_75t_L g5099 ( 
.A1(n_4986),
.A2(n_5039),
.A3(n_4985),
.B(n_4991),
.Y(n_5099)
);

AOI21xp5_ASAP7_75t_L g5100 ( 
.A1(n_5057),
.A2(n_738),
.B(n_739),
.Y(n_5100)
);

NAND4xp25_ASAP7_75t_L g5101 ( 
.A(n_5017),
.B(n_5010),
.C(n_5002),
.D(n_5034),
.Y(n_5101)
);

INVx2_ASAP7_75t_L g5102 ( 
.A(n_5029),
.Y(n_5102)
);

NOR2xp33_ASAP7_75t_L g5103 ( 
.A(n_5012),
.B(n_739),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_5005),
.Y(n_5104)
);

OAI21xp5_ASAP7_75t_L g5105 ( 
.A1(n_5027),
.A2(n_743),
.B(n_742),
.Y(n_5105)
);

AOI22xp5_ASAP7_75t_L g5106 ( 
.A1(n_5049),
.A2(n_743),
.B1(n_741),
.B2(n_742),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_5016),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_4999),
.Y(n_5108)
);

AOI22xp33_ASAP7_75t_L g5109 ( 
.A1(n_5011),
.A2(n_5024),
.B1(n_5022),
.B2(n_5043),
.Y(n_5109)
);

NAND2x1_ASAP7_75t_L g5110 ( 
.A(n_5009),
.B(n_741),
.Y(n_5110)
);

NOR3xp33_ASAP7_75t_L g5111 ( 
.A(n_4988),
.B(n_746),
.C(n_745),
.Y(n_5111)
);

NAND4xp75_ASAP7_75t_L g5112 ( 
.A(n_5052),
.B(n_747),
.C(n_744),
.D(n_746),
.Y(n_5112)
);

NOR4xp25_ASAP7_75t_L g5113 ( 
.A(n_5038),
.B(n_748),
.C(n_744),
.D(n_747),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_SL g5114 ( 
.A(n_5036),
.B(n_748),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4989),
.Y(n_5115)
);

NAND2xp5_ASAP7_75t_L g5116 ( 
.A(n_5046),
.B(n_749),
.Y(n_5116)
);

NAND3xp33_ASAP7_75t_L g5117 ( 
.A(n_5021),
.B(n_749),
.C(n_750),
.Y(n_5117)
);

AND2x2_ASAP7_75t_L g5118 ( 
.A(n_5023),
.B(n_750),
.Y(n_5118)
);

OAI22xp5_ASAP7_75t_L g5119 ( 
.A1(n_5018),
.A2(n_753),
.B1(n_751),
.B2(n_752),
.Y(n_5119)
);

OAI222xp33_ASAP7_75t_L g5120 ( 
.A1(n_4993),
.A2(n_755),
.B1(n_757),
.B2(n_752),
.C1(n_754),
.C2(n_756),
.Y(n_5120)
);

AOI221xp5_ASAP7_75t_L g5121 ( 
.A1(n_4994),
.A2(n_759),
.B1(n_754),
.B2(n_755),
.C(n_761),
.Y(n_5121)
);

OAI22xp5_ASAP7_75t_L g5122 ( 
.A1(n_5040),
.A2(n_5026),
.B1(n_5054),
.B2(n_4998),
.Y(n_5122)
);

AND2x2_ASAP7_75t_L g5123 ( 
.A(n_5028),
.B(n_759),
.Y(n_5123)
);

AO22x1_ASAP7_75t_L g5124 ( 
.A1(n_5000),
.A2(n_763),
.B1(n_761),
.B2(n_762),
.Y(n_5124)
);

INVx1_ASAP7_75t_L g5125 ( 
.A(n_4980),
.Y(n_5125)
);

AO22x2_ASAP7_75t_L g5126 ( 
.A1(n_5035),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.Y(n_5126)
);

AOI21xp5_ASAP7_75t_L g5127 ( 
.A1(n_5001),
.A2(n_764),
.B(n_765),
.Y(n_5127)
);

XNOR2x1_ASAP7_75t_SL g5128 ( 
.A(n_5019),
.B(n_5020),
.Y(n_5128)
);

NOR2x1_ASAP7_75t_L g5129 ( 
.A(n_5053),
.B(n_765),
.Y(n_5129)
);

AO22x2_ASAP7_75t_L g5130 ( 
.A1(n_5037),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.Y(n_5130)
);

INVx2_ASAP7_75t_L g5131 ( 
.A(n_5050),
.Y(n_5131)
);

INVx1_ASAP7_75t_L g5132 ( 
.A(n_4982),
.Y(n_5132)
);

OA22x2_ASAP7_75t_L g5133 ( 
.A1(n_5056),
.A2(n_769),
.B1(n_766),
.B2(n_768),
.Y(n_5133)
);

NOR2x1_ASAP7_75t_L g5134 ( 
.A(n_4979),
.B(n_769),
.Y(n_5134)
);

AOI21xp5_ASAP7_75t_L g5135 ( 
.A1(n_5060),
.A2(n_770),
.B(n_771),
.Y(n_5135)
);

AND2x4_ASAP7_75t_L g5136 ( 
.A(n_4982),
.B(n_770),
.Y(n_5136)
);

AOI21xp5_ASAP7_75t_L g5137 ( 
.A1(n_5060),
.A2(n_771),
.B(n_772),
.Y(n_5137)
);

NOR3xp33_ASAP7_75t_L g5138 ( 
.A(n_4990),
.B(n_774),
.C(n_773),
.Y(n_5138)
);

OAI21xp5_ASAP7_75t_L g5139 ( 
.A1(n_5060),
.A2(n_776),
.B(n_774),
.Y(n_5139)
);

OAI22xp33_ASAP7_75t_L g5140 ( 
.A1(n_5060),
.A2(n_778),
.B1(n_772),
.B2(n_777),
.Y(n_5140)
);

NAND3xp33_ASAP7_75t_L g5141 ( 
.A(n_4982),
.B(n_777),
.C(n_778),
.Y(n_5141)
);

AOI31xp33_ASAP7_75t_L g5142 ( 
.A1(n_5060),
.A2(n_788),
.A3(n_797),
.B(n_779),
.Y(n_5142)
);

AOI211x1_ASAP7_75t_SL g5143 ( 
.A1(n_4997),
.A2(n_782),
.B(n_780),
.C(n_781),
.Y(n_5143)
);

AO22x2_ASAP7_75t_L g5144 ( 
.A1(n_5047),
.A2(n_785),
.B1(n_782),
.B2(n_783),
.Y(n_5144)
);

NOR3xp33_ASAP7_75t_SL g5145 ( 
.A(n_5013),
.B(n_783),
.C(n_786),
.Y(n_5145)
);

OAI21xp33_ASAP7_75t_L g5146 ( 
.A1(n_5060),
.A2(n_786),
.B(n_787),
.Y(n_5146)
);

XNOR2x1_ASAP7_75t_SL g5147 ( 
.A(n_5033),
.B(n_789),
.Y(n_5147)
);

NOR3xp33_ASAP7_75t_L g5148 ( 
.A(n_4990),
.B(n_791),
.C(n_790),
.Y(n_5148)
);

OAI211xp5_ASAP7_75t_L g5149 ( 
.A1(n_4997),
.A2(n_792),
.B(n_789),
.C(n_791),
.Y(n_5149)
);

AOI21xp5_ASAP7_75t_L g5150 ( 
.A1(n_5065),
.A2(n_792),
.B(n_794),
.Y(n_5150)
);

HB1xp67_ASAP7_75t_L g5151 ( 
.A(n_5147),
.Y(n_5151)
);

AOI22xp5_ASAP7_75t_L g5152 ( 
.A1(n_5068),
.A2(n_796),
.B1(n_794),
.B2(n_795),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_5130),
.Y(n_5153)
);

AND2x2_ASAP7_75t_L g5154 ( 
.A(n_5071),
.B(n_795),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_5130),
.Y(n_5155)
);

INVxp67_ASAP7_75t_L g5156 ( 
.A(n_5069),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_L g5157 ( 
.A(n_5066),
.B(n_797),
.Y(n_5157)
);

INVxp67_ASAP7_75t_L g5158 ( 
.A(n_5134),
.Y(n_5158)
);

NOR2x1_ASAP7_75t_L g5159 ( 
.A(n_5141),
.B(n_798),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_5144),
.Y(n_5160)
);

NOR3xp33_ASAP7_75t_L g5161 ( 
.A(n_5099),
.B(n_798),
.C(n_799),
.Y(n_5161)
);

AOI221x1_ASAP7_75t_L g5162 ( 
.A1(n_5144),
.A2(n_801),
.B1(n_799),
.B2(n_800),
.C(n_802),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_5133),
.Y(n_5163)
);

OAI21xp5_ASAP7_75t_L g5164 ( 
.A1(n_5082),
.A2(n_802),
.B(n_803),
.Y(n_5164)
);

AOI22xp33_ASAP7_75t_L g5165 ( 
.A1(n_5131),
.A2(n_805),
.B1(n_803),
.B2(n_804),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_5064),
.Y(n_5166)
);

AND2x4_ASAP7_75t_L g5167 ( 
.A(n_5088),
.B(n_804),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_5136),
.Y(n_5168)
);

AOI22xp5_ASAP7_75t_L g5169 ( 
.A1(n_5070),
.A2(n_807),
.B1(n_805),
.B2(n_806),
.Y(n_5169)
);

NOR2xp33_ASAP7_75t_L g5170 ( 
.A(n_5077),
.B(n_808),
.Y(n_5170)
);

AOI22xp5_ASAP7_75t_L g5171 ( 
.A1(n_5125),
.A2(n_812),
.B1(n_808),
.B2(n_809),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_5126),
.Y(n_5172)
);

INVxp67_ASAP7_75t_SL g5173 ( 
.A(n_5129),
.Y(n_5173)
);

NAND2x1p5_ASAP7_75t_L g5174 ( 
.A(n_5114),
.B(n_812),
.Y(n_5174)
);

AOI211xp5_ASAP7_75t_L g5175 ( 
.A1(n_5149),
.A2(n_814),
.B(n_809),
.C(n_813),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_5124),
.B(n_813),
.Y(n_5176)
);

XNOR2xp5_ASAP7_75t_L g5177 ( 
.A(n_5128),
.B(n_814),
.Y(n_5177)
);

OAI21xp5_ASAP7_75t_L g5178 ( 
.A1(n_5085),
.A2(n_815),
.B(n_816),
.Y(n_5178)
);

CKINVDCx5p33_ASAP7_75t_R g5179 ( 
.A(n_5145),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_5126),
.Y(n_5180)
);

INVx2_ASAP7_75t_L g5181 ( 
.A(n_5087),
.Y(n_5181)
);

NAND3xp33_ASAP7_75t_SL g5182 ( 
.A(n_5074),
.B(n_5143),
.C(n_5078),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_5087),
.Y(n_5183)
);

NOR2xp33_ASAP7_75t_L g5184 ( 
.A(n_5146),
.B(n_817),
.Y(n_5184)
);

NAND2xp5_ASAP7_75t_L g5185 ( 
.A(n_5113),
.B(n_5142),
.Y(n_5185)
);

AOI22xp33_ASAP7_75t_L g5186 ( 
.A1(n_5102),
.A2(n_819),
.B1(n_817),
.B2(n_818),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_5132),
.Y(n_5187)
);

INVxp67_ASAP7_75t_L g5188 ( 
.A(n_5103),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_5118),
.Y(n_5189)
);

NOR2xp33_ASAP7_75t_L g5190 ( 
.A(n_5076),
.B(n_818),
.Y(n_5190)
);

OAI322xp33_ASAP7_75t_L g5191 ( 
.A1(n_5110),
.A2(n_825),
.A3(n_824),
.B1(n_822),
.B2(n_820),
.C1(n_821),
.C2(n_823),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_5083),
.B(n_820),
.Y(n_5192)
);

HB1xp67_ASAP7_75t_L g5193 ( 
.A(n_5112),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_5073),
.Y(n_5194)
);

OA22x2_ASAP7_75t_L g5195 ( 
.A1(n_5106),
.A2(n_823),
.B1(n_821),
.B2(n_822),
.Y(n_5195)
);

A2O1A1Ixp33_ASAP7_75t_L g5196 ( 
.A1(n_5062),
.A2(n_826),
.B(n_824),
.C(n_825),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_5080),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_5123),
.Y(n_5198)
);

NAND3xp33_ASAP7_75t_SL g5199 ( 
.A(n_5092),
.B(n_826),
.C(n_828),
.Y(n_5199)
);

OAI22xp5_ASAP7_75t_L g5200 ( 
.A1(n_5109),
.A2(n_830),
.B1(n_828),
.B2(n_829),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_5116),
.Y(n_5201)
);

NAND2xp5_ASAP7_75t_L g5202 ( 
.A(n_5140),
.B(n_830),
.Y(n_5202)
);

AOI21xp33_ASAP7_75t_SL g5203 ( 
.A1(n_5063),
.A2(n_831),
.B(n_832),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_5081),
.Y(n_5204)
);

OA22x2_ASAP7_75t_SL g5205 ( 
.A1(n_5097),
.A2(n_834),
.B1(n_831),
.B2(n_833),
.Y(n_5205)
);

AND2x2_ASAP7_75t_L g5206 ( 
.A(n_5098),
.B(n_834),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_5096),
.Y(n_5207)
);

AOI21xp33_ASAP7_75t_L g5208 ( 
.A1(n_5122),
.A2(n_835),
.B(n_836),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_5117),
.Y(n_5209)
);

NOR2x1_ASAP7_75t_L g5210 ( 
.A(n_5120),
.B(n_835),
.Y(n_5210)
);

AOI211xp5_ASAP7_75t_L g5211 ( 
.A1(n_5101),
.A2(n_5105),
.B(n_5079),
.C(n_5100),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5104),
.Y(n_5212)
);

NAND3xp33_ASAP7_75t_L g5213 ( 
.A(n_5138),
.B(n_836),
.C(n_837),
.Y(n_5213)
);

NAND2xp5_ASAP7_75t_L g5214 ( 
.A(n_5067),
.B(n_839),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_5072),
.Y(n_5215)
);

NAND3xp33_ASAP7_75t_L g5216 ( 
.A(n_5148),
.B(n_840),
.C(n_841),
.Y(n_5216)
);

INVx2_ASAP7_75t_L g5217 ( 
.A(n_5108),
.Y(n_5217)
);

AND2x2_ASAP7_75t_L g5218 ( 
.A(n_5139),
.B(n_840),
.Y(n_5218)
);

INVx1_ASAP7_75t_SL g5219 ( 
.A(n_5135),
.Y(n_5219)
);

NOR3xp33_ASAP7_75t_L g5220 ( 
.A(n_5089),
.B(n_842),
.C(n_843),
.Y(n_5220)
);

NAND3xp33_ASAP7_75t_L g5221 ( 
.A(n_5111),
.B(n_842),
.C(n_843),
.Y(n_5221)
);

XNOR2xp5_ASAP7_75t_L g5222 ( 
.A(n_5084),
.B(n_844),
.Y(n_5222)
);

XNOR2xp5_ASAP7_75t_L g5223 ( 
.A(n_5119),
.B(n_844),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_5137),
.B(n_5127),
.Y(n_5224)
);

NOR2x1_ASAP7_75t_L g5225 ( 
.A(n_5075),
.B(n_845),
.Y(n_5225)
);

INVx2_ASAP7_75t_L g5226 ( 
.A(n_5094),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_5177),
.Y(n_5227)
);

INVx2_ASAP7_75t_L g5228 ( 
.A(n_5205),
.Y(n_5228)
);

INVx2_ASAP7_75t_L g5229 ( 
.A(n_5167),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_5151),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_5160),
.B(n_5153),
.Y(n_5231)
);

AOI31xp33_ASAP7_75t_L g5232 ( 
.A1(n_5174),
.A2(n_5086),
.A3(n_5107),
.B(n_5095),
.Y(n_5232)
);

NAND2xp5_ASAP7_75t_SL g5233 ( 
.A(n_5172),
.B(n_5091),
.Y(n_5233)
);

INVxp67_ASAP7_75t_L g5234 ( 
.A(n_5157),
.Y(n_5234)
);

INVx2_ASAP7_75t_L g5235 ( 
.A(n_5167),
.Y(n_5235)
);

AOI22xp5_ASAP7_75t_L g5236 ( 
.A1(n_5161),
.A2(n_5115),
.B1(n_5090),
.B2(n_5121),
.Y(n_5236)
);

AOI22xp5_ASAP7_75t_L g5237 ( 
.A1(n_5179),
.A2(n_5093),
.B1(n_847),
.B2(n_845),
.Y(n_5237)
);

NOR2x1_ASAP7_75t_L g5238 ( 
.A(n_5180),
.B(n_846),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5154),
.Y(n_5239)
);

NAND2xp5_ASAP7_75t_SL g5240 ( 
.A(n_5156),
.B(n_846),
.Y(n_5240)
);

NAND2xp5_ASAP7_75t_L g5241 ( 
.A(n_5155),
.B(n_848),
.Y(n_5241)
);

AOI22xp5_ASAP7_75t_L g5242 ( 
.A1(n_5163),
.A2(n_851),
.B1(n_848),
.B2(n_849),
.Y(n_5242)
);

NAND2xp5_ASAP7_75t_L g5243 ( 
.A(n_5183),
.B(n_849),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_5176),
.Y(n_5244)
);

NAND2xp5_ASAP7_75t_L g5245 ( 
.A(n_5181),
.B(n_851),
.Y(n_5245)
);

INVx1_ASAP7_75t_L g5246 ( 
.A(n_5206),
.Y(n_5246)
);

NOR2xp33_ASAP7_75t_SL g5247 ( 
.A(n_5210),
.B(n_5158),
.Y(n_5247)
);

AOI221xp5_ASAP7_75t_L g5248 ( 
.A1(n_5203),
.A2(n_854),
.B1(n_852),
.B2(n_853),
.C(n_856),
.Y(n_5248)
);

NOR2xp33_ASAP7_75t_L g5249 ( 
.A(n_5191),
.B(n_852),
.Y(n_5249)
);

AO22x2_ASAP7_75t_L g5250 ( 
.A1(n_5162),
.A2(n_856),
.B1(n_853),
.B2(n_854),
.Y(n_5250)
);

OAI22xp5_ASAP7_75t_SL g5251 ( 
.A1(n_5185),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.Y(n_5251)
);

AOI22xp5_ASAP7_75t_L g5252 ( 
.A1(n_5170),
.A2(n_860),
.B1(n_858),
.B2(n_859),
.Y(n_5252)
);

NAND2xp33_ASAP7_75t_L g5253 ( 
.A(n_5220),
.B(n_860),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_5195),
.Y(n_5254)
);

NOR2x1_ASAP7_75t_L g5255 ( 
.A(n_5168),
.B(n_861),
.Y(n_5255)
);

AOI22xp5_ASAP7_75t_L g5256 ( 
.A1(n_5182),
.A2(n_864),
.B1(n_862),
.B2(n_863),
.Y(n_5256)
);

OAI31xp33_ASAP7_75t_SL g5257 ( 
.A1(n_5173),
.A2(n_5225),
.A3(n_5159),
.B(n_5199),
.Y(n_5257)
);

AOI22xp5_ASAP7_75t_L g5258 ( 
.A1(n_5215),
.A2(n_866),
.B1(n_862),
.B2(n_864),
.Y(n_5258)
);

AOI221xp5_ASAP7_75t_L g5259 ( 
.A1(n_5187),
.A2(n_868),
.B1(n_866),
.B2(n_867),
.C(n_869),
.Y(n_5259)
);

INVxp67_ASAP7_75t_SL g5260 ( 
.A(n_5192),
.Y(n_5260)
);

AOI22xp5_ASAP7_75t_L g5261 ( 
.A1(n_5212),
.A2(n_5209),
.B1(n_5217),
.B2(n_5189),
.Y(n_5261)
);

NAND2xp5_ASAP7_75t_SL g5262 ( 
.A(n_5175),
.B(n_867),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_5193),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_5202),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_5214),
.Y(n_5265)
);

NAND2xp5_ASAP7_75t_L g5266 ( 
.A(n_5150),
.B(n_869),
.Y(n_5266)
);

AOI22xp5_ASAP7_75t_L g5267 ( 
.A1(n_5207),
.A2(n_872),
.B1(n_870),
.B2(n_871),
.Y(n_5267)
);

AOI22xp5_ASAP7_75t_L g5268 ( 
.A1(n_5184),
.A2(n_873),
.B1(n_870),
.B2(n_871),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_5223),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_5218),
.Y(n_5270)
);

AOI221xp5_ASAP7_75t_L g5271 ( 
.A1(n_5208),
.A2(n_876),
.B1(n_873),
.B2(n_874),
.C(n_877),
.Y(n_5271)
);

NOR2xp33_ASAP7_75t_L g5272 ( 
.A(n_5198),
.B(n_874),
.Y(n_5272)
);

NOR4xp25_ASAP7_75t_L g5273 ( 
.A(n_5219),
.B(n_880),
.C(n_878),
.D(n_879),
.Y(n_5273)
);

AOI22xp5_ASAP7_75t_L g5274 ( 
.A1(n_5190),
.A2(n_883),
.B1(n_878),
.B2(n_882),
.Y(n_5274)
);

INVx1_ASAP7_75t_L g5275 ( 
.A(n_5152),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_5222),
.Y(n_5276)
);

AOI22xp5_ASAP7_75t_L g5277 ( 
.A1(n_5226),
.A2(n_886),
.B1(n_882),
.B2(n_884),
.Y(n_5277)
);

AOI221xp5_ASAP7_75t_L g5278 ( 
.A1(n_5164),
.A2(n_887),
.B1(n_884),
.B2(n_886),
.C(n_888),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5169),
.Y(n_5279)
);

NOR4xp25_ASAP7_75t_L g5280 ( 
.A(n_5224),
.B(n_890),
.C(n_888),
.D(n_889),
.Y(n_5280)
);

AOI221xp5_ASAP7_75t_L g5281 ( 
.A1(n_5178),
.A2(n_892),
.B1(n_889),
.B2(n_890),
.C(n_893),
.Y(n_5281)
);

AND2x2_ASAP7_75t_L g5282 ( 
.A(n_5165),
.B(n_892),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_5250),
.Y(n_5283)
);

AOI22xp33_ASAP7_75t_SL g5284 ( 
.A1(n_5247),
.A2(n_5166),
.B1(n_5197),
.B2(n_5194),
.Y(n_5284)
);

NAND2xp5_ASAP7_75t_L g5285 ( 
.A(n_5280),
.B(n_5200),
.Y(n_5285)
);

INVx1_ASAP7_75t_L g5286 ( 
.A(n_5250),
.Y(n_5286)
);

AOI322xp5_ASAP7_75t_L g5287 ( 
.A1(n_5230),
.A2(n_5188),
.A3(n_5204),
.B1(n_5201),
.B2(n_5196),
.C1(n_5186),
.C2(n_5171),
.Y(n_5287)
);

OAI22xp5_ASAP7_75t_L g5288 ( 
.A1(n_5256),
.A2(n_5213),
.B1(n_5216),
.B2(n_5221),
.Y(n_5288)
);

INVx1_ASAP7_75t_SL g5289 ( 
.A(n_5255),
.Y(n_5289)
);

NOR2xp33_ASAP7_75t_R g5290 ( 
.A(n_5254),
.B(n_5211),
.Y(n_5290)
);

AOI21xp33_ASAP7_75t_L g5291 ( 
.A1(n_5231),
.A2(n_893),
.B(n_894),
.Y(n_5291)
);

NOR2xp33_ASAP7_75t_R g5292 ( 
.A(n_5227),
.B(n_894),
.Y(n_5292)
);

AOI21xp5_ASAP7_75t_L g5293 ( 
.A1(n_5233),
.A2(n_895),
.B(n_896),
.Y(n_5293)
);

OR2x2_ASAP7_75t_L g5294 ( 
.A(n_5273),
.B(n_897),
.Y(n_5294)
);

HB1xp67_ASAP7_75t_L g5295 ( 
.A(n_5238),
.Y(n_5295)
);

INVx1_ASAP7_75t_SL g5296 ( 
.A(n_5229),
.Y(n_5296)
);

NOR2x1_ASAP7_75t_L g5297 ( 
.A(n_5235),
.B(n_5228),
.Y(n_5297)
);

AOI211xp5_ASAP7_75t_L g5298 ( 
.A1(n_5249),
.A2(n_900),
.B(n_897),
.C(n_898),
.Y(n_5298)
);

AOI322xp5_ASAP7_75t_L g5299 ( 
.A1(n_5263),
.A2(n_904),
.A3(n_903),
.B1(n_901),
.B2(n_898),
.C1(n_900),
.C2(n_902),
.Y(n_5299)
);

OAI22xp33_ASAP7_75t_L g5300 ( 
.A1(n_5261),
.A2(n_904),
.B1(n_901),
.B2(n_903),
.Y(n_5300)
);

BUFx2_ASAP7_75t_L g5301 ( 
.A(n_5251),
.Y(n_5301)
);

NOR2xp33_ASAP7_75t_L g5302 ( 
.A(n_5239),
.B(n_905),
.Y(n_5302)
);

AOI21xp5_ASAP7_75t_L g5303 ( 
.A1(n_5257),
.A2(n_905),
.B(n_906),
.Y(n_5303)
);

NAND2xp5_ASAP7_75t_L g5304 ( 
.A(n_5272),
.B(n_907),
.Y(n_5304)
);

NAND4xp25_ASAP7_75t_SL g5305 ( 
.A(n_5236),
.B(n_910),
.C(n_908),
.D(n_909),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_5242),
.B(n_908),
.Y(n_5306)
);

AND2x2_ASAP7_75t_SL g5307 ( 
.A(n_5253),
.B(n_909),
.Y(n_5307)
);

AND2x2_ASAP7_75t_L g5308 ( 
.A(n_5282),
.B(n_911),
.Y(n_5308)
);

INVx2_ASAP7_75t_SL g5309 ( 
.A(n_5240),
.Y(n_5309)
);

NOR2x1_ASAP7_75t_L g5310 ( 
.A(n_5243),
.B(n_911),
.Y(n_5310)
);

OAI211xp5_ASAP7_75t_SL g5311 ( 
.A1(n_5234),
.A2(n_914),
.B(n_912),
.C(n_913),
.Y(n_5311)
);

AOI22xp5_ASAP7_75t_L g5312 ( 
.A1(n_5246),
.A2(n_914),
.B1(n_912),
.B2(n_913),
.Y(n_5312)
);

AND2x2_ASAP7_75t_L g5313 ( 
.A(n_5260),
.B(n_915),
.Y(n_5313)
);

NAND4xp25_ASAP7_75t_L g5314 ( 
.A(n_5275),
.B(n_918),
.C(n_915),
.D(n_916),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_5258),
.B(n_916),
.Y(n_5315)
);

OAI221xp5_ASAP7_75t_L g5316 ( 
.A1(n_5241),
.A2(n_921),
.B1(n_918),
.B2(n_919),
.C(n_922),
.Y(n_5316)
);

BUFx6f_ASAP7_75t_L g5317 ( 
.A(n_5245),
.Y(n_5317)
);

OAI22xp5_ASAP7_75t_SL g5318 ( 
.A1(n_5307),
.A2(n_5252),
.B1(n_5266),
.B2(n_5244),
.Y(n_5318)
);

AND2x4_ASAP7_75t_L g5319 ( 
.A(n_5297),
.B(n_5270),
.Y(n_5319)
);

NOR2xp33_ASAP7_75t_L g5320 ( 
.A(n_5296),
.B(n_5232),
.Y(n_5320)
);

NAND4xp75_ASAP7_75t_L g5321 ( 
.A(n_5310),
.B(n_5276),
.C(n_5269),
.D(n_5264),
.Y(n_5321)
);

INVx2_ASAP7_75t_L g5322 ( 
.A(n_5294),
.Y(n_5322)
);

INVx1_ASAP7_75t_L g5323 ( 
.A(n_5295),
.Y(n_5323)
);

AND2x2_ASAP7_75t_L g5324 ( 
.A(n_5308),
.B(n_5279),
.Y(n_5324)
);

INVx2_ASAP7_75t_L g5325 ( 
.A(n_5313),
.Y(n_5325)
);

INVx1_ASAP7_75t_L g5326 ( 
.A(n_5283),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_5286),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_L g5328 ( 
.A(n_5302),
.B(n_5248),
.Y(n_5328)
);

NAND4xp75_ASAP7_75t_L g5329 ( 
.A(n_5303),
.B(n_5265),
.C(n_5262),
.D(n_5271),
.Y(n_5329)
);

AND2x2_ASAP7_75t_L g5330 ( 
.A(n_5301),
.B(n_5237),
.Y(n_5330)
);

AOI22xp5_ASAP7_75t_L g5331 ( 
.A1(n_5309),
.A2(n_5281),
.B1(n_5278),
.B2(n_5274),
.Y(n_5331)
);

AOI211x1_ASAP7_75t_L g5332 ( 
.A1(n_5293),
.A2(n_5268),
.B(n_5259),
.C(n_5267),
.Y(n_5332)
);

OR2x2_ASAP7_75t_L g5333 ( 
.A(n_5289),
.B(n_5277),
.Y(n_5333)
);

NOR2x1_ASAP7_75t_L g5334 ( 
.A(n_5314),
.B(n_919),
.Y(n_5334)
);

INVxp67_ASAP7_75t_L g5335 ( 
.A(n_5305),
.Y(n_5335)
);

OAI211xp5_ASAP7_75t_SL g5336 ( 
.A1(n_5326),
.A2(n_5287),
.B(n_5284),
.C(n_5298),
.Y(n_5336)
);

OAI221xp5_ASAP7_75t_L g5337 ( 
.A1(n_5327),
.A2(n_5285),
.B1(n_5306),
.B2(n_5315),
.C(n_5288),
.Y(n_5337)
);

AND2x4_ASAP7_75t_L g5338 ( 
.A(n_5319),
.B(n_5317),
.Y(n_5338)
);

OAI22xp5_ASAP7_75t_L g5339 ( 
.A1(n_5323),
.A2(n_5304),
.B1(n_5317),
.B2(n_5300),
.Y(n_5339)
);

INVx2_ASAP7_75t_L g5340 ( 
.A(n_5325),
.Y(n_5340)
);

AOI211xp5_ASAP7_75t_L g5341 ( 
.A1(n_5320),
.A2(n_5291),
.B(n_5311),
.C(n_5290),
.Y(n_5341)
);

OAI22xp5_ASAP7_75t_SL g5342 ( 
.A1(n_5318),
.A2(n_5316),
.B1(n_5317),
.B2(n_5312),
.Y(n_5342)
);

AOI211xp5_ASAP7_75t_L g5343 ( 
.A1(n_5335),
.A2(n_5292),
.B(n_5299),
.C(n_923),
.Y(n_5343)
);

NOR3xp33_ASAP7_75t_L g5344 ( 
.A(n_5321),
.B(n_921),
.C(n_922),
.Y(n_5344)
);

OAI22xp5_ASAP7_75t_L g5345 ( 
.A1(n_5331),
.A2(n_925),
.B1(n_923),
.B2(n_924),
.Y(n_5345)
);

NAND3xp33_ASAP7_75t_L g5346 ( 
.A(n_5334),
.B(n_5330),
.C(n_5324),
.Y(n_5346)
);

OAI211xp5_ASAP7_75t_SL g5347 ( 
.A1(n_5333),
.A2(n_928),
.B(n_925),
.C(n_927),
.Y(n_5347)
);

NAND3xp33_ASAP7_75t_L g5348 ( 
.A(n_5344),
.B(n_5322),
.C(n_5332),
.Y(n_5348)
);

INVx4_ASAP7_75t_L g5349 ( 
.A(n_5338),
.Y(n_5349)
);

OAI21xp5_ASAP7_75t_L g5350 ( 
.A1(n_5346),
.A2(n_5329),
.B(n_5328),
.Y(n_5350)
);

NOR3xp33_ASAP7_75t_SL g5351 ( 
.A(n_5336),
.B(n_927),
.C(n_928),
.Y(n_5351)
);

OR2x2_ASAP7_75t_L g5352 ( 
.A(n_5340),
.B(n_929),
.Y(n_5352)
);

XNOR2x1_ASAP7_75t_SL g5353 ( 
.A(n_5341),
.B(n_929),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5342),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_5347),
.Y(n_5355)
);

INVx1_ASAP7_75t_SL g5356 ( 
.A(n_5352),
.Y(n_5356)
);

BUFx2_ASAP7_75t_L g5357 ( 
.A(n_5349),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_5353),
.Y(n_5358)
);

NAND2xp5_ASAP7_75t_L g5359 ( 
.A(n_5351),
.B(n_5343),
.Y(n_5359)
);

OR3x2_ASAP7_75t_L g5360 ( 
.A(n_5354),
.B(n_5337),
.C(n_5339),
.Y(n_5360)
);

AOI22x1_ASAP7_75t_L g5361 ( 
.A1(n_5357),
.A2(n_5350),
.B1(n_5355),
.B2(n_5348),
.Y(n_5361)
);

OAI22xp5_ASAP7_75t_L g5362 ( 
.A1(n_5360),
.A2(n_5345),
.B1(n_932),
.B2(n_930),
.Y(n_5362)
);

OAI221xp5_ASAP7_75t_L g5363 ( 
.A1(n_5361),
.A2(n_5358),
.B1(n_5359),
.B2(n_5356),
.C(n_933),
.Y(n_5363)
);

OA21x2_ASAP7_75t_L g5364 ( 
.A1(n_5363),
.A2(n_5362),
.B(n_931),
.Y(n_5364)
);

HB1xp67_ASAP7_75t_L g5365 ( 
.A(n_5364),
.Y(n_5365)
);

OAI21x1_ASAP7_75t_L g5366 ( 
.A1(n_5365),
.A2(n_931),
.B(n_932),
.Y(n_5366)
);

OAI22xp33_ASAP7_75t_L g5367 ( 
.A1(n_5366),
.A2(n_935),
.B1(n_933),
.B2(n_934),
.Y(n_5367)
);

NAND2xp5_ASAP7_75t_L g5368 ( 
.A(n_5367),
.B(n_934),
.Y(n_5368)
);

INVx1_ASAP7_75t_L g5369 ( 
.A(n_5368),
.Y(n_5369)
);

AOI22xp33_ASAP7_75t_SL g5370 ( 
.A1(n_5368),
.A2(n_937),
.B1(n_935),
.B2(n_936),
.Y(n_5370)
);

NAND2xp5_ASAP7_75t_L g5371 ( 
.A(n_5370),
.B(n_936),
.Y(n_5371)
);

OA21x2_ASAP7_75t_L g5372 ( 
.A1(n_5369),
.A2(n_937),
.B(n_938),
.Y(n_5372)
);

AOI21xp5_ASAP7_75t_L g5373 ( 
.A1(n_5371),
.A2(n_938),
.B(n_939),
.Y(n_5373)
);

AOI211xp5_ASAP7_75t_L g5374 ( 
.A1(n_5373),
.A2(n_5372),
.B(n_940),
.C(n_939),
.Y(n_5374)
);


endmodule