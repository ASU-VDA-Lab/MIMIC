module fake_jpeg_2166_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_SL g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx8_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_14),
.B(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_19),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_15),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_17),
.A2(n_10),
.B1(n_13),
.B2(n_18),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_6),
.B1(n_7),
.B2(n_12),
.Y(n_18)
);

OAI21x1_ASAP7_75t_R g25 ( 
.A1(n_18),
.A2(n_23),
.B(n_24),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_7),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_10),
.B1(n_7),
.B2(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_25),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_18),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_31),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_18),
.Y(n_33)
);

INVxp33_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_13),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_26),
.B1(n_29),
.B2(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_35),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_43),
.B1(n_42),
.B2(n_36),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_42),
.Y(n_46)
);


endmodule