module fake_jpeg_3036_n_182 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_182);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_0),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_56),
.B1(n_46),
.B2(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_80),
.B1(n_49),
.B2(n_53),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_55),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_45),
.B1(n_61),
.B2(n_56),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_45),
.B1(n_61),
.B2(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_47),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_100),
.B1(n_75),
.B2(n_40),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_95),
.Y(n_109)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_3),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_53),
.B1(n_51),
.B2(n_57),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_97),
.A2(n_77),
.B1(n_84),
.B2(n_83),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_5),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_101)
);

OR2x2_ASAP7_75t_SL g110 ( 
.A(n_101),
.B(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_110),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_74),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_74),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_77),
.B(n_4),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_111),
.B(n_114),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_75),
.B1(n_43),
.B2(n_42),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_75),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_28),
.Y(n_139)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_125),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_118),
.A2(n_90),
.B1(n_94),
.B2(n_92),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_98),
.B1(n_7),
.B2(n_8),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_102),
.B1(n_120),
.B2(n_107),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_39),
.C(n_38),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_131),
.C(n_138),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_36),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_6),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_31),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_17),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_29),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_26),
.B1(n_22),
.B2(n_21),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_140),
.A2(n_111),
.B1(n_107),
.B2(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_150),
.Y(n_160)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_152),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_114),
.B1(n_10),
.B2(n_11),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_149),
.B1(n_155),
.B2(n_131),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_149)
);

AOI21x1_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_13),
.B(n_14),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_13),
.C(n_14),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_155)
);

OAI322xp33_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_18),
.A3(n_19),
.B1(n_20),
.B2(n_130),
.C1(n_154),
.C2(n_152),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_164),
.B1(n_157),
.B2(n_163),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_141),
.C(n_153),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_140),
.B1(n_137),
.B2(n_138),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_141),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_162),
.B(n_146),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_169),
.B1(n_162),
.B2(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_166),
.B(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_153),
.Y(n_174)
);

AOI31xp67_ASAP7_75t_SL g176 ( 
.A1(n_174),
.A2(n_175),
.A3(n_167),
.B(n_160),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_158),
.C(n_164),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_173),
.C(n_151),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_159),
.C(n_19),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g180 ( 
.A(n_179),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_18),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_20),
.Y(n_182)
);


endmodule