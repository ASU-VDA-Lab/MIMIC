module real_aes_8476_n_254 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_254);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_254;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_693;
wire n_496;
wire n_281;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_756;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_740;
wire n_371;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_668;
wire n_797;
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_0), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_1), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_2), .A2(n_201), .B1(n_399), .B2(n_489), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_3), .A2(n_17), .B1(n_431), .B2(n_432), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_4), .A2(n_164), .B1(n_472), .B2(n_475), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_5), .A2(n_220), .B1(n_501), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_6), .A2(n_55), .B1(n_463), .B2(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g494 ( .A(n_7), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_8), .A2(n_410), .B1(n_445), .B2(n_446), .Y(n_409) );
INVx1_ASAP7_75t_L g445 ( .A(n_8), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_9), .A2(n_226), .B1(n_303), .B2(n_535), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_10), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_11), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g616 ( .A(n_12), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_13), .A2(n_123), .B1(n_438), .B2(n_698), .Y(n_790) );
OA22x2_ASAP7_75t_L g586 ( .A1(n_14), .A2(n_587), .B1(n_588), .B2(n_617), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_14), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_15), .A2(n_140), .B1(n_566), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_16), .A2(n_97), .B1(n_475), .B2(n_535), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_18), .A2(n_22), .B1(n_326), .B2(n_393), .C(n_396), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_19), .A2(n_60), .B1(n_442), .B2(n_444), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_20), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_21), .B(n_667), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_23), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_24), .A2(n_72), .B1(n_326), .B2(n_329), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_25), .A2(n_187), .B1(n_471), .B2(n_474), .Y(n_470) );
INVx1_ASAP7_75t_L g652 ( .A(n_26), .Y(n_652) );
AO22x2_ASAP7_75t_L g278 ( .A1(n_27), .A2(n_78), .B1(n_279), .B2(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g738 ( .A(n_27), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_28), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_29), .A2(n_142), .B1(n_443), .B2(n_623), .Y(n_622) );
AOI222xp33_ASAP7_75t_L g541 ( .A1(n_30), .A2(n_95), .B1(n_115), .B2(n_369), .C1(n_454), .C2(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_31), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_32), .A2(n_223), .B1(n_350), .B2(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g719 ( .A(n_33), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_34), .A2(n_85), .B1(n_236), .B2(n_297), .C1(n_309), .C2(n_633), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_35), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_36), .A2(n_174), .B1(n_309), .B2(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g614 ( .A(n_37), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_38), .A2(n_49), .B1(n_484), .B2(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_39), .A2(n_199), .B1(n_348), .B2(n_487), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_40), .A2(n_149), .B1(n_329), .B2(n_524), .Y(n_523) );
AO22x2_ASAP7_75t_L g282 ( .A1(n_41), .A2(n_82), .B1(n_279), .B2(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g739 ( .A(n_41), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_42), .A2(n_119), .B1(n_440), .B2(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g607 ( .A(n_43), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_44), .A2(n_252), .B1(n_381), .B2(n_384), .C(n_385), .Y(n_380) );
INVx1_ASAP7_75t_L g599 ( .A(n_45), .Y(n_599) );
INVx1_ASAP7_75t_L g606 ( .A(n_46), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_47), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_48), .A2(n_134), .B1(n_442), .B2(n_444), .Y(n_441) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_50), .A2(n_132), .B1(n_399), .B2(n_431), .Y(n_679) );
INVx1_ASAP7_75t_L g355 ( .A(n_51), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_52), .B(n_667), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_53), .Y(n_803) );
AOI22xp5_ASAP7_75t_SL g639 ( .A1(n_54), .A2(n_242), .B1(n_597), .B2(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g397 ( .A(n_56), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_57), .A2(n_108), .B1(n_438), .B2(n_440), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_58), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_59), .A2(n_202), .B1(n_333), .B2(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_61), .A2(n_81), .B1(n_342), .B2(n_435), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_62), .A2(n_244), .B1(n_309), .B2(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_63), .B(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_64), .A2(n_238), .B1(n_471), .B2(n_649), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_65), .Y(n_361) );
OA22x2_ASAP7_75t_L g660 ( .A1(n_66), .A2(n_661), .B1(n_662), .B2(n_682), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_66), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_67), .B(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_68), .A2(n_153), .B1(n_480), .B2(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g582 ( .A(n_69), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_70), .A2(n_175), .B1(n_326), .B2(n_381), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_71), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_73), .A2(n_148), .B1(n_342), .B2(n_346), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_74), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_75), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g477 ( .A1(n_76), .A2(n_107), .B1(n_383), .B2(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_77), .A2(n_245), .B1(n_465), .B2(n_533), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_79), .A2(n_131), .B1(n_333), .B2(n_336), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_80), .A2(n_83), .B1(n_475), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_84), .A2(n_241), .B1(n_383), .B2(n_507), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_86), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_87), .A2(n_196), .B1(n_381), .B2(n_489), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g669 ( .A1(n_88), .A2(n_214), .B1(n_633), .B2(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g262 ( .A(n_89), .Y(n_262) );
AOI211xp5_ASAP7_75t_L g254 ( .A1(n_90), .A2(n_255), .B(n_264), .C(n_740), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_91), .A2(n_118), .B1(n_538), .B2(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_92), .B(n_467), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_93), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_93), .A2(n_782), .B1(n_787), .B2(n_812), .Y(n_786) );
INVx1_ASAP7_75t_L g260 ( .A(n_94), .Y(n_260) );
INVx1_ASAP7_75t_L g655 ( .A(n_96), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_98), .A2(n_136), .B1(n_346), .B2(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_99), .A2(n_163), .B1(n_344), .B2(n_439), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_100), .A2(n_109), .B1(n_487), .B2(n_630), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_101), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_102), .Y(n_273) );
INVx1_ASAP7_75t_L g721 ( .A(n_103), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_104), .B(n_423), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_105), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_106), .A2(n_158), .B1(n_303), .B2(n_309), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_110), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_111), .A2(n_211), .B1(n_540), .B2(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g715 ( .A(n_112), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_113), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_114), .A2(n_169), .B1(n_594), .B2(n_597), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_116), .A2(n_203), .B1(n_754), .B2(n_756), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_117), .Y(n_377) );
INVx1_ASAP7_75t_L g591 ( .A(n_120), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_121), .A2(n_124), .B1(n_326), .B2(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g717 ( .A(n_122), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_125), .A2(n_160), .B1(n_689), .B2(n_690), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_126), .B(n_578), .Y(n_577) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_127), .A2(n_172), .B1(n_178), .B2(n_298), .C1(n_303), .C2(n_423), .Y(n_722) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_128), .A2(n_165), .B1(n_205), .B2(n_298), .C1(n_372), .C2(n_496), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_129), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_130), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_133), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_135), .A2(n_742), .B1(n_772), .B2(n_773), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_135), .Y(n_772) );
AOI22xp33_ASAP7_75t_SL g488 ( .A1(n_137), .A2(n_176), .B1(n_403), .B2(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g263 ( .A(n_138), .Y(n_263) );
AO22x1_ASAP7_75t_L g357 ( .A1(n_139), .A2(n_358), .B1(n_404), .B2(n_405), .Y(n_357) );
INVx1_ASAP7_75t_L g404 ( .A(n_139), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_141), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_143), .A2(n_253), .B1(n_496), .B2(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_144), .A2(n_151), .B1(n_432), .B2(n_681), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_145), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_146), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_147), .A2(n_237), .B1(n_526), .B2(n_527), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_150), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_152), .A2(n_231), .B1(n_474), .B2(n_670), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_154), .A2(n_248), .B1(n_597), .B2(n_677), .Y(n_676) );
AND2x6_ASAP7_75t_L g259 ( .A(n_155), .B(n_260), .Y(n_259) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_155), .Y(n_732) );
AO22x2_ASAP7_75t_L g288 ( .A1(n_156), .A2(n_218), .B1(n_279), .B2(n_283), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_157), .A2(n_243), .B1(n_690), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g457 ( .A1(n_159), .A2(n_192), .B1(n_423), .B2(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_161), .B(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_162), .A2(n_217), .B1(n_350), .B2(n_352), .Y(n_349) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_166), .A2(n_250), .B1(n_484), .B2(n_485), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_167), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_168), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_170), .A2(n_247), .B1(n_395), .B2(n_524), .Y(n_696) );
INVx1_ASAP7_75t_L g709 ( .A(n_171), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_173), .Y(n_544) );
INVx1_ASAP7_75t_L g723 ( .A(n_177), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_179), .B(n_372), .Y(n_371) );
AO22x2_ASAP7_75t_L g286 ( .A1(n_180), .A2(n_228), .B1(n_279), .B2(n_280), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_181), .A2(n_213), .B1(n_444), .B2(n_754), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_182), .Y(n_571) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_183), .A2(n_233), .B1(n_352), .B2(n_395), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_184), .Y(n_425) );
XOR2x2_ASAP7_75t_L g684 ( .A(n_185), .B(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_186), .A2(n_190), .B1(n_333), .B2(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g401 ( .A(n_188), .Y(n_401) );
INVx1_ASAP7_75t_L g613 ( .A(n_189), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_191), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_193), .A2(n_235), .B1(n_633), .B2(n_670), .Y(n_712) );
INVx1_ASAP7_75t_L g317 ( .A(n_194), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_195), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_197), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_198), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_200), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_204), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_206), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_207), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_208), .B(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_209), .Y(n_747) );
INVx1_ASAP7_75t_L g592 ( .A(n_210), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_212), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_215), .Y(n_580) );
XOR2x2_ASAP7_75t_L g449 ( .A(n_216), .B(n_450), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_218), .B(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_219), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_221), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_222), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_224), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_225), .A2(n_234), .B1(n_435), .B2(n_698), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_227), .Y(n_386) );
INVx1_ASAP7_75t_L g735 ( .A(n_228), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_229), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_230), .A2(n_249), .B1(n_463), .B2(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g456 ( .A(n_232), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_239), .Y(n_413) );
INVx1_ASAP7_75t_L g279 ( .A(n_240), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_240), .Y(n_281) );
INVx1_ASAP7_75t_L g600 ( .A(n_246), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_251), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_256), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_257), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_260), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_261), .A2(n_730), .B(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_658), .B1(n_725), .B2(n_726), .C(n_727), .Y(n_264) );
INVx1_ASAP7_75t_L g725 ( .A(n_265), .Y(n_725) );
OAI22xp5_ASAP7_75t_SL g265 ( .A1(n_266), .A2(n_267), .B1(n_515), .B2(n_516), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
XOR2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_407), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_356), .B1(n_357), .B2(n_406), .Y(n_268) );
INVx2_ASAP7_75t_SL g406 ( .A(n_269), .Y(n_406) );
XOR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_355), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_323), .Y(n_270) );
NOR3xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_294), .C(n_312), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_289), .B2(n_290), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_274), .A2(n_290), .B1(n_580), .B2(n_581), .Y(n_579) );
BUFx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g363 ( .A(n_275), .Y(n_363) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_275), .Y(n_414) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_284), .Y(n_275) );
INVx2_ASAP7_75t_L g345 ( .A(n_276), .Y(n_345) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_282), .Y(n_276) );
AND2x2_ASAP7_75t_L g293 ( .A(n_277), .B(n_282), .Y(n_293) );
AND2x2_ASAP7_75t_L g328 ( .A(n_277), .B(n_307), .Y(n_328) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g299 ( .A(n_278), .B(n_282), .Y(n_299) );
AND2x2_ASAP7_75t_L g308 ( .A(n_278), .B(n_288), .Y(n_308) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g283 ( .A(n_281), .Y(n_283) );
INVx2_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
INVx1_ASAP7_75t_L g338 ( .A(n_282), .Y(n_338) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_285), .B(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g351 ( .A(n_285), .B(n_328), .Y(n_351) );
AND2x6_ASAP7_75t_L g465 ( .A(n_285), .B(n_293), .Y(n_465) );
AND2x4_ASAP7_75t_L g469 ( .A(n_285), .B(n_345), .Y(n_469) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g301 ( .A(n_286), .Y(n_301) );
INVx1_ASAP7_75t_L g306 ( .A(n_286), .Y(n_306) );
INVx1_ASAP7_75t_L g322 ( .A(n_286), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_286), .B(n_288), .Y(n_339) );
AND2x2_ASAP7_75t_L g300 ( .A(n_287), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g331 ( .A(n_288), .B(n_322), .Y(n_331) );
OAI221xp5_ASAP7_75t_L g604 ( .A1(n_290), .A2(n_605), .B1(n_606), .B2(n_607), .C(n_608), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_290), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_SL g365 ( .A(n_291), .Y(n_365) );
INVx2_ASAP7_75t_L g811 ( .A(n_291), .Y(n_811) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g531 ( .A(n_292), .Y(n_531) );
AND2x2_ASAP7_75t_L g335 ( .A(n_293), .B(n_331), .Y(n_335) );
AND2x4_ASAP7_75t_L g348 ( .A(n_293), .B(n_300), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_293), .B(n_331), .Y(n_388) );
OAI21xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_302), .Y(n_294) );
OAI221xp5_ASAP7_75t_L g366 ( .A1(n_296), .A2(n_367), .B1(n_368), .B2(n_370), .C(n_371), .Y(n_366) );
OAI21xp5_ASAP7_75t_SL g493 ( .A1(n_296), .A2(n_494), .B(n_495), .Y(n_493) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_296), .A2(n_665), .B(n_666), .Y(n_664) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_298), .Y(n_418) );
INVx4_ASAP7_75t_L g455 ( .A(n_298), .Y(n_455) );
INVx2_ASAP7_75t_SL g763 ( .A(n_298), .Y(n_763) );
AND2x6_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g319 ( .A(n_299), .Y(n_319) );
AND2x4_ASAP7_75t_L g475 ( .A(n_299), .B(n_321), .Y(n_475) );
AND2x2_ASAP7_75t_L g327 ( .A(n_300), .B(n_328), .Y(n_327) );
AND2x6_ASAP7_75t_L g344 ( .A(n_300), .B(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_303), .Y(n_369) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_304), .Y(n_460) );
BUFx4f_ASAP7_75t_SL g496 ( .A(n_304), .Y(n_496) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_304), .Y(n_578) );
BUFx2_ASAP7_75t_L g654 ( .A(n_304), .Y(n_654) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g311 ( .A(n_306), .Y(n_311) );
INVx1_ASAP7_75t_L g316 ( .A(n_307), .Y(n_316) );
AND2x4_ASAP7_75t_L g310 ( .A(n_308), .B(n_311), .Y(n_310) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_308), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g472 ( .A(n_308), .B(n_473), .Y(n_472) );
BUFx4f_ASAP7_75t_SL g372 ( .A(n_309), .Y(n_372) );
INVx2_ASAP7_75t_L g543 ( .A(n_309), .Y(n_543) );
BUFx12f_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_310), .Y(n_423) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_310), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_317), .B2(n_318), .Y(n_312) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx4_ASAP7_75t_L g376 ( .A(n_315), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_315), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_315), .A2(n_378), .B1(n_802), .B2(n_803), .Y(n_801) );
AND2x2_ASAP7_75t_L g507 ( .A(n_316), .B(n_354), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g379 ( .A(n_318), .Y(n_379) );
BUFx2_ASAP7_75t_L g427 ( .A(n_318), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_318), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
OR2x6_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_340), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_332), .Y(n_324) );
BUFx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_327), .Y(n_439) );
INVx2_ASAP7_75t_L g513 ( .A(n_327), .Y(n_513) );
BUFx2_ASAP7_75t_SL g538 ( .A(n_327), .Y(n_538) );
AND2x2_ASAP7_75t_L g330 ( .A(n_328), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g353 ( .A(n_328), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_328), .B(n_331), .Y(n_561) );
BUFx3_ASAP7_75t_L g431 ( .A(n_329), .Y(n_431) );
BUFx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx3_ASAP7_75t_L g395 ( .A(n_330), .Y(n_395) );
BUFx3_ASAP7_75t_L g487 ( .A(n_330), .Y(n_487) );
BUFx3_ASAP7_75t_L g603 ( .A(n_330), .Y(n_603) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_333), .Y(n_677) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx5_ASAP7_75t_L g443 ( .A(n_334), .Y(n_443) );
INVx3_ASAP7_75t_L g526 ( .A(n_334), .Y(n_526) );
INVx4_ASAP7_75t_L g596 ( .A(n_334), .Y(n_596) );
BUFx3_ASAP7_75t_L g707 ( .A(n_334), .Y(n_707) );
INVx1_ASAP7_75t_L g755 ( .A(n_334), .Y(n_755) );
INVx8_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx4f_ASAP7_75t_SL g391 ( .A(n_336), .Y(n_391) );
BUFx2_ASAP7_75t_L g444 ( .A(n_336), .Y(n_444) );
BUFx2_ASAP7_75t_L g527 ( .A(n_336), .Y(n_527) );
BUFx2_ASAP7_75t_L g597 ( .A(n_336), .Y(n_597) );
BUFx2_ASAP7_75t_L g690 ( .A(n_336), .Y(n_690) );
INVx6_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g554 ( .A(n_337), .Y(n_554) );
INVx1_ASAP7_75t_SL g756 ( .A(n_337), .Y(n_756) );
OR2x6_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g473 ( .A(n_338), .Y(n_473) );
INVx1_ASAP7_75t_L g354 ( .A(n_339), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_349), .Y(n_340) );
INVx4_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_SL g480 ( .A(n_343), .Y(n_480) );
INVx2_ASAP7_75t_L g643 ( .A(n_343), .Y(n_643) );
INVx1_ASAP7_75t_L g698 ( .A(n_343), .Y(n_698) );
INVx11_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx11_ASAP7_75t_L g400 ( .A(n_344), .Y(n_400) );
INVx1_ASAP7_75t_L g557 ( .A(n_346), .Y(n_557) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g403 ( .A(n_347), .Y(n_403) );
INVx2_ASAP7_75t_L g435 ( .A(n_347), .Y(n_435) );
INVx6_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx3_ASAP7_75t_L g540 ( .A(n_348), .Y(n_540) );
BUFx3_ASAP7_75t_L g623 ( .A(n_348), .Y(n_623) );
BUFx2_ASAP7_75t_L g675 ( .A(n_350), .Y(n_675) );
BUFx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_351), .Y(n_383) );
BUFx3_ASAP7_75t_L g440 ( .A(n_351), .Y(n_440) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx3_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
BUFx3_ASAP7_75t_L g433 ( .A(n_353), .Y(n_433) );
BUFx2_ASAP7_75t_SL g489 ( .A(n_353), .Y(n_489) );
BUFx3_ASAP7_75t_L g524 ( .A(n_353), .Y(n_524) );
BUFx2_ASAP7_75t_SL g566 ( .A(n_353), .Y(n_566) );
BUFx3_ASAP7_75t_L g630 ( .A(n_353), .Y(n_630) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g405 ( .A(n_358), .Y(n_405) );
AND3x1_ASAP7_75t_L g358 ( .A(n_359), .B(n_380), .C(n_392), .Y(n_358) );
NOR3xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_366), .C(n_373), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B1(n_364), .B2(n_365), .Y(n_360) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g605 ( .A(n_363), .Y(n_605) );
INVx2_ASAP7_75t_L g760 ( .A(n_363), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_365), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_412) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_SL g420 ( .A(n_369), .Y(n_420) );
INVx1_ASAP7_75t_L g615 ( .A(n_372), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_377), .B2(n_378), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_375), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx3_ASAP7_75t_SL g570 ( .A(n_376), .Y(n_570) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g771 ( .A(n_379), .Y(n_771) );
INVx4_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_382), .A2(n_563), .B1(n_564), .B2(n_565), .Y(n_562) );
OAI221xp5_ASAP7_75t_SL g589 ( .A1(n_382), .A2(n_590), .B1(n_591), .B2(n_592), .C(n_593), .Y(n_589) );
INVx3_ASAP7_75t_L g704 ( .A(n_382), .Y(n_704) );
INVx4_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_389), .B2(n_390), .Y(n_385) );
BUFx2_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B1(n_401), .B2(n_402), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx4_ASAP7_75t_L g510 ( .A(n_400), .Y(n_510) );
INVx3_ASAP7_75t_L g552 ( .A(n_400), .Y(n_552) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_400), .A2(n_402), .B1(n_599), .B2(n_600), .C(n_601), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_402), .A2(n_793), .B1(n_794), .B2(n_795), .Y(n_792) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_447), .B2(n_448), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g446 ( .A(n_410), .Y(n_446) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_428), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_416), .C(n_424), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_414), .A2(n_809), .B1(n_810), .B2(n_811), .Y(n_808) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_420), .B2(n_421), .C(n_422), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g804 ( .A1(n_420), .A2(n_453), .B1(n_805), .B2(n_806), .C(n_807), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_436), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_434), .Y(n_429) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_441), .Y(n_436) );
BUFx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_439), .Y(n_484) );
INVx3_ASAP7_75t_L g590 ( .A(n_439), .Y(n_590) );
INVx1_ASAP7_75t_L g798 ( .A(n_440), .Y(n_798) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_443), .Y(n_689) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
XNOR2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_490), .Y(n_448) );
NAND3x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_476), .C(n_482), .Y(n_450) );
NOR2x1_ASAP7_75t_SL g451 ( .A(n_452), .B(n_461), .Y(n_451) );
OAI21xp5_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_456), .B(n_457), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx4_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_455), .A2(n_573), .B1(n_574), .B2(n_576), .C(n_577), .Y(n_572) );
OAI222xp33_ASAP7_75t_L g611 ( .A1(n_455), .A2(n_612), .B1(n_613), .B2(n_614), .C1(n_615), .C2(n_616), .Y(n_611) );
BUFx2_ASAP7_75t_L g651 ( .A(n_455), .Y(n_651) );
INVx1_ASAP7_75t_L g612 ( .A(n_458), .Y(n_612) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx4_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_466), .C(n_470), .Y(n_461) );
INVx1_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g672 ( .A(n_464), .Y(n_672) );
INVx1_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
BUFx4f_ASAP7_75t_L g499 ( .A(n_465), .Y(n_499) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g501 ( .A(n_468), .Y(n_501) );
INVx5_ASAP7_75t_L g533 ( .A(n_468), .Y(n_533) );
INVx2_ASAP7_75t_L g647 ( .A(n_468), .Y(n_647) );
INVx4_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g535 ( .A(n_472), .Y(n_535) );
INVx1_ASAP7_75t_L g610 ( .A(n_472), .Y(n_610) );
BUFx2_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
BUFx3_ASAP7_75t_L g633 ( .A(n_475), .Y(n_633) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_475), .Y(n_649) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_488), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
XOR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_514), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_492), .B(n_503), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_497), .Y(n_492) );
INVx1_ASAP7_75t_L g765 ( .A(n_496), .Y(n_765) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .C(n_502), .Y(n_497) );
BUFx2_ASAP7_75t_L g711 ( .A(n_501), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_508), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g681 ( .A(n_513), .Y(n_681) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B1(n_583), .B2(n_584), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g518 ( .A1(n_519), .A2(n_520), .B1(n_545), .B2(n_546), .Y(n_518) );
INVx3_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
XOR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_544), .Y(n_520) );
NAND4xp75_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .C(n_536), .D(n_541), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVxp67_ASAP7_75t_L g716 ( .A(n_524), .Y(n_716) );
OA211x2_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_532), .C(n_534), .Y(n_528) );
OA211x2_ASAP7_75t_L g708 ( .A1(n_530), .A2(n_709), .B(n_710), .C(n_712), .Y(n_708) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_533), .Y(n_693) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
INVx1_ASAP7_75t_L g750 ( .A(n_540), .Y(n_750) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
XOR2xp5_ASAP7_75t_SL g547 ( .A(n_548), .B(n_582), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_567), .Y(n_548) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_555), .C(n_562), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
INVx1_ASAP7_75t_L g720 ( .A(n_552), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_557), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_559), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_714) );
OAI221xp5_ASAP7_75t_SL g749 ( .A1(n_559), .A2(n_750), .B1(n_751), .B2(n_752), .C(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g795 ( .A(n_560), .Y(n_795) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
NOR3xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .C(n_579), .Y(n_567) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g667 ( .A(n_575), .Y(n_667) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_618), .B1(n_656), .B2(n_657), .Y(n_585) );
INVx1_ASAP7_75t_L g656 ( .A(n_586), .Y(n_656) );
INVx1_ASAP7_75t_L g617 ( .A(n_588), .Y(n_617) );
OR4x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_598), .C(n_604), .D(n_611), .Y(n_588) );
OAI221xp5_ASAP7_75t_SL g744 ( .A1(n_590), .A2(n_745), .B1(n_746), .B2(n_747), .C(n_748), .Y(n_744) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_596), .Y(n_640) );
BUFx4f_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g670 ( .A(n_610), .Y(n_670) );
INVx1_ASAP7_75t_L g657 ( .A(n_618), .Y(n_657) );
XNOR2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_635), .Y(n_618) );
XOR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_634), .Y(n_619) );
NAND4xp75_ASAP7_75t_L g620 ( .A(n_621), .B(n_625), .C(n_628), .D(n_632), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_SL g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
XOR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_655), .Y(n_635) );
NOR4xp75_ASAP7_75t_L g636 ( .A(n_637), .B(n_641), .C(n_645), .D(n_650), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NAND2x1_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_646), .B(n_648), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B(n_653), .Y(n_650) );
CKINVDCx16_ASAP7_75t_R g726 ( .A(n_658), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_683), .B2(n_724), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g682 ( .A(n_662), .Y(n_682) );
NAND3x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_673), .C(n_678), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_668), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g746 ( .A(n_675), .Y(n_746) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g724 ( .A(n_683), .Y(n_724) );
XOR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_700), .Y(n_683) );
NAND4xp75_ASAP7_75t_L g685 ( .A(n_686), .B(n_691), .C(n_695), .D(n_699), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
AND2x2_ASAP7_75t_SL g691 ( .A(n_692), .B(n_694), .Y(n_691) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
XOR2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_723), .Y(n_700) );
NAND4xp75_ASAP7_75t_L g701 ( .A(n_702), .B(n_708), .C(n_713), .D(n_722), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
INVx3_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_718), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_716), .A2(n_797), .B1(n_798), .B2(n_799), .Y(n_796) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
NOR2x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_733), .Y(n_728) );
OR2x2_ASAP7_75t_SL g815 ( .A(n_729), .B(n_734), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_731), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_731), .B(n_778), .Y(n_781) );
CKINVDCx16_ASAP7_75t_R g778 ( .A(n_732), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
OAI322xp33_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_774), .A3(n_775), .B1(n_779), .B2(n_782), .C1(n_783), .C2(n_813), .Y(n_740) );
INVx2_ASAP7_75t_L g773 ( .A(n_742), .Y(n_773) );
AND2x2_ASAP7_75t_SL g742 ( .A(n_743), .B(n_757), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_749), .Y(n_743) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NOR3xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_762), .C(n_768), .Y(n_757) );
OAI221xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B1(n_765), .B2(n_766), .C(n_767), .Y(n_762) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
CKINVDCx16_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g812 ( .A(n_787), .Y(n_812) );
AND2x2_ASAP7_75t_SL g787 ( .A(n_788), .B(n_800), .Y(n_787) );
NOR3xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_792), .C(n_796), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
NOR3xp33_ASAP7_75t_SL g800 ( .A(n_801), .B(n_804), .C(n_808), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
endmodule