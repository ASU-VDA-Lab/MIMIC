module fake_jpeg_15269_n_389 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_389);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_389;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_45),
.Y(n_69)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_60),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_15),
.B(n_0),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_62),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_24),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_68),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_20),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_71),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_72),
.B(n_84),
.Y(n_141)
);

BUFx12f_ASAP7_75t_SL g73 ( 
.A(n_49),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_73),
.A2(n_85),
.B1(n_109),
.B2(n_32),
.Y(n_149)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_74),
.B(n_89),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_16),
.B1(n_21),
.B2(n_17),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_76),
.A2(n_86),
.B(n_110),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_54),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_83),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_20),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_43),
.A2(n_25),
.B1(n_37),
.B2(n_20),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_16),
.B1(n_21),
.B2(n_25),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_45),
.Y(n_89)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_16),
.B1(n_25),
.B2(n_37),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_93),
.A2(n_106),
.B1(n_29),
.B2(n_26),
.Y(n_163)
);

CKINVDCx6p67_ASAP7_75t_R g94 ( 
.A(n_59),
.Y(n_94)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_19),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_108),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_27),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_38),
.A2(n_16),
.B1(n_28),
.B2(n_34),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_52),
.B(n_36),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_27),
.B1(n_18),
.B2(n_23),
.Y(n_110)
);

AND2x4_ASAP7_75t_SL g111 ( 
.A(n_52),
.B(n_0),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_111),
.A2(n_29),
.B(n_26),
.C(n_3),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_44),
.A2(n_35),
.B1(n_34),
.B2(n_30),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_22),
.B1(n_35),
.B2(n_34),
.Y(n_121)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_64),
.Y(n_148)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_15),
.C(n_32),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_15),
.C(n_32),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_121),
.A2(n_123),
.B1(n_138),
.B2(n_164),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_19),
.B1(n_35),
.B2(n_22),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_126),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_69),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_133),
.Y(n_177)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_132),
.A2(n_168),
.B1(n_79),
.B2(n_95),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_158),
.C(n_61),
.Y(n_174)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_19),
.B1(n_22),
.B2(n_30),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_72),
.B(n_30),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_139),
.B(n_147),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_144),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_151),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_96),
.B(n_29),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_163),
.B1(n_79),
.B2(n_90),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_18),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_152),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_23),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_77),
.B(n_23),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_160),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_78),
.B(n_63),
.C(n_62),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_83),
.Y(n_159)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_91),
.B(n_18),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_165),
.B(n_4),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_78),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_106),
.A2(n_1),
.B(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_75),
.B(n_39),
.Y(n_166)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_166),
.B(n_5),
.CI(n_7),
.CON(n_213),
.SN(n_213)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_104),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_1),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_170),
.B1(n_117),
.B2(n_103),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_80),
.B(n_3),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_174),
.B(n_180),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_82),
.B1(n_95),
.B2(n_118),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_179),
.A2(n_190),
.B1(n_192),
.B2(n_196),
.Y(n_236)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_40),
.A3(n_39),
.B1(n_80),
.B2(n_70),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_195),
.Y(n_218)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_188),
.B(n_191),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_186),
.B(n_189),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_129),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_102),
.B1(n_74),
.B2(n_103),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_90),
.B1(n_107),
.B2(n_87),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_160),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_137),
.A2(n_107),
.B1(n_39),
.B2(n_6),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_149),
.A2(n_116),
.B1(n_5),
.B2(n_6),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_202),
.B1(n_152),
.B2(n_154),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_153),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_122),
.B(n_4),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_162),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_153),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_212),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_170),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_116),
.C(n_104),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_145),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_150),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_169),
.B1(n_170),
.B2(n_134),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_135),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_141),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_124),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_214),
.A2(n_140),
.B1(n_132),
.B2(n_124),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_215),
.B(n_223),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_224),
.B1(n_228),
.B2(n_234),
.Y(n_259)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_220),
.A2(n_232),
.B1(n_248),
.B2(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_225),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_150),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_239),
.Y(n_265)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_131),
.B1(n_169),
.B2(n_133),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_175),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_229),
.B(n_233),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_237),
.C(n_206),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_178),
.B(n_194),
.CI(n_174),
.CON(n_231),
.SN(n_231)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_213),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_182),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_235),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_178),
.B(n_163),
.Y(n_237)
);

AO21x2_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_196),
.B(n_180),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_208),
.B1(n_197),
.B2(n_187),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_144),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_193),
.B(n_130),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_243),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_181),
.A2(n_142),
.B(n_128),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_244),
.A2(n_205),
.B(n_140),
.Y(n_281)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_245),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_193),
.B(n_121),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_254),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_173),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_181),
.A2(n_167),
.B1(n_140),
.B2(n_135),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_249),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_203),
.A2(n_136),
.B1(n_157),
.B2(n_156),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_179),
.B1(n_190),
.B2(n_161),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_267),
.C(n_268),
.Y(n_288)
);

AO21x1_ASAP7_75t_L g304 ( 
.A1(n_257),
.A2(n_284),
.B(n_244),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_258),
.A2(n_253),
.B1(n_224),
.B2(n_218),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_263),
.A2(n_225),
.B1(n_221),
.B2(n_216),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_188),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_264),
.B(n_270),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_226),
.A2(n_185),
.B(n_186),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_266),
.A2(n_275),
.B(n_281),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_177),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_231),
.C(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_189),
.Y(n_272)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_238),
.A2(n_212),
.B1(n_187),
.B2(n_198),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_273),
.A2(n_282),
.B1(n_283),
.B2(n_249),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_201),
.B(n_176),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_199),
.C(n_173),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_279),
.C(n_274),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_205),
.C(n_202),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_238),
.A2(n_171),
.B1(n_127),
.B2(n_200),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_238),
.A2(n_236),
.B1(n_253),
.B2(n_219),
.Y(n_283)
);

OR2x6_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_223),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_222),
.B(n_171),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_289),
.A2(n_281),
.B1(n_279),
.B2(n_257),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_290),
.A2(n_292),
.B1(n_293),
.B2(n_295),
.Y(n_316)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_291),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_264),
.A2(n_235),
.B1(n_243),
.B2(n_215),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_269),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_299),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_259),
.A2(n_254),
.B1(n_241),
.B2(n_240),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_304),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_256),
.A2(n_251),
.B(n_220),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_297),
.A2(n_313),
.B(n_287),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_256),
.B1(n_282),
.B2(n_283),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_298),
.A2(n_300),
.B1(n_308),
.B2(n_309),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_232),
.B1(n_216),
.B2(n_245),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_247),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_306),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_227),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_261),
.B(n_8),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_307),
.Y(n_332)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_273),
.B(n_260),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_265),
.B(n_9),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_310),
.A2(n_312),
.B(n_305),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_10),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_312),
.B(n_286),
.Y(n_317)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_255),
.B(n_268),
.C(n_267),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_10),
.C(n_275),
.Y(n_315)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_298),
.A2(n_284),
.B1(n_258),
.B2(n_277),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_319),
.A2(n_324),
.B1(n_327),
.B2(n_334),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_270),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_325),
.Y(n_343)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_300),
.A2(n_284),
.B(n_285),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_323),
.A2(n_331),
.B(n_333),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_278),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_299),
.A2(n_280),
.B1(n_287),
.B2(n_302),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_311),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_325),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_303),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_297),
.A2(n_295),
.B(n_293),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_292),
.A2(n_301),
.B1(n_302),
.B2(n_290),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_301),
.A2(n_303),
.B1(n_304),
.B2(n_296),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_315),
.Y(n_338)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_338),
.B(n_344),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_291),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_340),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_336),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_288),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_351),
.C(n_353),
.Y(n_359)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_320),
.B(n_331),
.C(n_330),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_321),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_335),
.C(n_324),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_348),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_347),
.A2(n_323),
.B(n_317),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_334),
.Y(n_348)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_347),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_328),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_349),
.B(n_329),
.Y(n_354)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_354),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_316),
.B1(n_326),
.B2(n_319),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_363),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_322),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_353),
.C(n_351),
.Y(n_368)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_342),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_349),
.B(n_326),
.Y(n_364)
);

INVx6_ASAP7_75t_L g370 ( 
.A(n_364),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_365),
.A2(n_366),
.B(n_341),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_368),
.B(n_371),
.C(n_359),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_357),
.A2(n_345),
.B(n_350),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_369),
.A2(n_362),
.B(n_360),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_343),
.Y(n_371)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_372),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_369),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_374),
.B(n_373),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_378),
.C(n_368),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_376),
.B(n_372),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_356),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_380),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_381),
.B(n_371),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_382),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_384),
.A2(n_379),
.B(n_377),
.Y(n_385)
);

AOI221xp5_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_374),
.B1(n_370),
.B2(n_355),
.C(n_344),
.Y(n_386)
);

AO21x1_ASAP7_75t_L g387 ( 
.A1(n_386),
.A2(n_355),
.B(n_370),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_387),
.B(n_359),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_343),
.Y(n_389)
);


endmodule