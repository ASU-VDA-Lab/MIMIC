module fake_netlist_6_4479_n_1080 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1080);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1080;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_1058;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_982;
wire n_831;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_60),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_179),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_117),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_90),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_26),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_165),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_25),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_32),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_91),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_129),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_13),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_17),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_76),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_71),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_62),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_135),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_46),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_82),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_182),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_105),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_126),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_33),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_160),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_12),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_153),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_35),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_61),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_136),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_1),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_13),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_87),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_198),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_12),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_168),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_47),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_204),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_45),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_42),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_67),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_20),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_15),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_164),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_132),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_30),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_103),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_173),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_15),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_156),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_172),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_121),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_66),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_152),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_122),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_207),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_109),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_97),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_202),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_190),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_88),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_199),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_10),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_218),
.Y(n_281)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_229),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_254),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_218),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_209),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_220),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_251),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_214),
.B(n_0),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_221),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_223),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_225),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_241),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_247),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_235),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_248),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_259),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_210),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_258),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_226),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_211),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_208),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_215),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_244),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_226),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_244),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_226),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_226),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_237),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_237),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_216),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_242),
.Y(n_325)
);

BUFx2_ASAP7_75t_SL g326 ( 
.A(n_257),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_237),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_212),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_217),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_217),
.Y(n_330)
);

BUFx8_ASAP7_75t_SL g331 ( 
.A(n_287),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_290),
.B(n_252),
.Y(n_332)
);

OA21x2_ASAP7_75t_L g333 ( 
.A1(n_308),
.A2(n_219),
.B(n_213),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_282),
.B(n_252),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_308),
.A2(n_279),
.B(n_228),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_284),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

OAI21x1_ASAP7_75t_L g340 ( 
.A1(n_319),
.A2(n_279),
.B(n_230),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_282),
.A2(n_263),
.B1(n_264),
.B2(n_238),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_289),
.B(n_295),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

CKINVDCx11_ASAP7_75t_R g346 ( 
.A(n_287),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_323),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_305),
.B(n_222),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_281),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_231),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_297),
.A2(n_256),
.B1(n_274),
.B2(n_273),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_294),
.B(n_232),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_297),
.A2(n_298),
.B1(n_302),
.B2(n_301),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_311),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_329),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_293),
.A2(n_278),
.B1(n_272),
.B2(n_271),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_296),
.A2(n_270),
.B1(n_269),
.B2(n_267),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_285),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_286),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_283),
.A2(n_303),
.B1(n_302),
.B2(n_298),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_299),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_301),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_304),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_291),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_310),
.B(n_233),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_311),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_330),
.A2(n_265),
.B1(n_262),
.B2(n_261),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_309),
.B(n_234),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_291),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_300),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_306),
.B(n_307),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_288),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_312),
.B(n_236),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_313),
.B(n_255),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_315),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_292),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_309),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_328),
.B(n_239),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_314),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_325),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_324),
.B(n_243),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_334),
.B(n_384),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

NAND2xp33_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_349),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_384),
.B(n_245),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_344),
.B(n_246),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_350),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_339),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_344),
.B(n_249),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_341),
.Y(n_399)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_337),
.Y(n_400)
);

INVxp33_ASAP7_75t_SL g401 ( 
.A(n_342),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_347),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_352),
.B(n_253),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_339),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_352),
.B(n_0),
.Y(n_405)
);

NOR2x1p5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_1),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_344),
.B(n_2),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_364),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_344),
.B(n_31),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_364),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

NAND3xp33_ASAP7_75t_L g415 ( 
.A(n_342),
.B(n_2),
.C(n_3),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_372),
.B(n_34),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_337),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_337),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_337),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_381),
.B(n_3),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_383),
.B(n_4),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_375),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_331),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_343),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_345),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_353),
.B(n_36),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_345),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_361),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_380),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_360),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_362),
.B(n_37),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_349),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_368),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_383),
.B(n_5),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_SL g444 ( 
.A(n_368),
.B(n_332),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_353),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_359),
.B(n_6),
.Y(n_446)
);

INVx8_ASAP7_75t_L g447 ( 
.A(n_353),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_360),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_341),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_380),
.Y(n_450)
);

OAI22xp33_ASAP7_75t_L g451 ( 
.A1(n_357),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_353),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_341),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_377),
.B(n_38),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_360),
.Y(n_456)
);

OAI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_351),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_348),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_358),
.B(n_10),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_371),
.B(n_11),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_360),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_402),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_402),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_389),
.B(n_382),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_392),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_418),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_418),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_395),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_392),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_410),
.A2(n_333),
.B(n_340),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_421),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_435),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_442),
.B(n_354),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_433),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_409),
.B(n_354),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_438),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_406),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_426),
.B(n_369),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_398),
.B(n_366),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_391),
.B(n_363),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_409),
.B(n_377),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_426),
.B(n_385),
.Y(n_489)
);

XNOR2x2_ASAP7_75t_L g490 ( 
.A(n_415),
.B(n_355),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_453),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_393),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_461),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_391),
.B(n_377),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_403),
.B(n_388),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_441),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_396),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_412),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_401),
.B(n_385),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_393),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_394),
.B(n_388),
.Y(n_501)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_407),
.B(n_377),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_424),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_427),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_444),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_427),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_428),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_422),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_444),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_413),
.B(n_378),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_428),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_430),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_401),
.B(n_355),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_445),
.B(n_386),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_445),
.B(n_452),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_430),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_413),
.B(n_386),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_460),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_R g522 ( 
.A(n_410),
.B(n_365),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_432),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_446),
.B(n_356),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_434),
.Y(n_525)
);

XNOR2x1_ASAP7_75t_L g526 ( 
.A(n_439),
.B(n_387),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_429),
.B(n_387),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_459),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_452),
.B(n_378),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_434),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_423),
.B(n_378),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_SL g532 ( 
.A(n_443),
.B(n_365),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_SL g533 ( 
.A(n_455),
.B(n_378),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_416),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_437),
.B(n_335),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_397),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_408),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_408),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_422),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_457),
.B(n_346),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_411),
.Y(n_541)
);

AND3x1_ASAP7_75t_L g542 ( 
.A(n_487),
.B(n_379),
.C(n_451),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_476),
.B(n_447),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_475),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g545 ( 
.A1(n_487),
.A2(n_447),
.B1(n_340),
.B2(n_437),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_469),
.B(n_447),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_503),
.A2(n_333),
.B1(n_447),
.B2(n_411),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_494),
.B(n_417),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_494),
.A2(n_333),
.B1(n_462),
.B2(n_456),
.Y(n_549)
);

NOR2x1p5_ASAP7_75t_L g550 ( 
.A(n_524),
.B(n_379),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_503),
.A2(n_490),
.B1(n_510),
.B2(n_463),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_510),
.B(n_502),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_469),
.B(n_333),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_477),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_519),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_390),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_465),
.B(n_390),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_517),
.A2(n_414),
.B(n_417),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_480),
.B(n_419),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_478),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_464),
.B(n_390),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_480),
.B(n_419),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_474),
.B(n_379),
.C(n_370),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_480),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_486),
.B(n_362),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_481),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_467),
.B(n_431),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_482),
.B(n_420),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_479),
.Y(n_569)
);

AND2x6_ASAP7_75t_SL g570 ( 
.A(n_495),
.B(n_11),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_482),
.B(n_420),
.Y(n_571)
);

NAND3xp33_ASAP7_75t_L g572 ( 
.A(n_486),
.B(n_516),
.C(n_496),
.Y(n_572)
);

A2O1A1Ixp33_ASAP7_75t_L g573 ( 
.A1(n_531),
.A2(n_335),
.B(n_462),
.C(n_456),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_484),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_482),
.B(n_436),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_496),
.A2(n_440),
.B1(n_436),
.B2(n_448),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_529),
.B(n_440),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_468),
.B(n_431),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_535),
.B(n_448),
.Y(n_579)
);

O2A1O1Ixp5_ASAP7_75t_L g580 ( 
.A1(n_471),
.A2(n_454),
.B(n_404),
.C(n_414),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_497),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_507),
.B(n_370),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_472),
.B(n_454),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_521),
.B(n_454),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_481),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_488),
.B(n_373),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_523),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_485),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_473),
.B(n_404),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_491),
.B(n_414),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_535),
.B(n_399),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_537),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_538),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_525),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_530),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_533),
.A2(n_373),
.B1(n_367),
.B2(n_399),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_466),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_493),
.B(n_399),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_511),
.B(n_367),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_SL g600 ( 
.A(n_582),
.B(n_528),
.C(n_501),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_544),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_555),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_581),
.B(n_488),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_553),
.A2(n_471),
.B(n_541),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_551),
.B(n_504),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_565),
.B(n_512),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_554),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_552),
.B(n_539),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_564),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_566),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_SL g611 ( 
.A(n_572),
.B(n_522),
.C(n_532),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_R g612 ( 
.A(n_599),
.B(n_498),
.Y(n_612)
);

AND2x4_ASAP7_75t_SL g613 ( 
.A(n_543),
.B(n_512),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_551),
.B(n_505),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_560),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_564),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_552),
.B(n_515),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_L g618 ( 
.A(n_546),
.B(n_527),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_550),
.A2(n_526),
.B1(n_499),
.B2(n_506),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_553),
.B(n_508),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_556),
.B(n_542),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_569),
.A2(n_513),
.B1(n_509),
.B2(n_514),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_557),
.B(n_518),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_R g624 ( 
.A(n_585),
.B(n_574),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_588),
.B(n_470),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_586),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_570),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_587),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_589),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_586),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_592),
.B(n_492),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_584),
.B(n_540),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_593),
.Y(n_633)
);

O2A1O1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_573),
.A2(n_536),
.B(n_520),
.C(n_500),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_584),
.B(n_483),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_594),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_595),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_543),
.B(n_489),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_543),
.B(n_399),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_586),
.B(n_367),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_597),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_575),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_561),
.Y(n_643)
);

NOR3xp33_ASAP7_75t_SL g644 ( 
.A(n_563),
.B(n_14),
.C(n_16),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_575),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_R g646 ( 
.A(n_598),
.B(n_39),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_583),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_559),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_567),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_R g650 ( 
.A(n_578),
.B(n_40),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_577),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_620),
.A2(n_548),
.B(n_604),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_611),
.A2(n_545),
.B(n_547),
.C(n_549),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_639),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_634),
.A2(n_580),
.B(n_548),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_602),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_603),
.B(n_559),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_600),
.A2(n_547),
.B1(n_576),
.B2(n_590),
.Y(n_658)
);

BUFx12f_ASAP7_75t_L g659 ( 
.A(n_602),
.Y(n_659)
);

CKINVDCx8_ASAP7_75t_R g660 ( 
.A(n_602),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_610),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_617),
.B(n_596),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_634),
.A2(n_558),
.B(n_579),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_604),
.A2(n_579),
.B(n_568),
.Y(n_664)
);

AOI221xp5_ASAP7_75t_SL g665 ( 
.A1(n_618),
.A2(n_596),
.B1(n_562),
.B2(n_571),
.C(n_568),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_608),
.B(n_591),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_625),
.Y(n_667)
);

AND2x6_ASAP7_75t_L g668 ( 
.A(n_651),
.B(n_591),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_601),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_606),
.B(n_562),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_621),
.A2(n_400),
.B(n_399),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_625),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_624),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_605),
.A2(n_400),
.B(n_449),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_607),
.Y(n_675)
);

AOI21xp33_ASAP7_75t_L g676 ( 
.A1(n_635),
.A2(n_14),
.B(n_16),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_631),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_603),
.B(n_449),
.Y(n_678)
);

A2O1A1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_611),
.A2(n_458),
.B(n_449),
.C(n_348),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_639),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_631),
.Y(n_681)
);

NAND2x1p5_ASAP7_75t_L g682 ( 
.A(n_609),
.B(n_449),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_615),
.Y(n_683)
);

NAND2x1_ASAP7_75t_L g684 ( 
.A(n_639),
.B(n_449),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_623),
.A2(n_458),
.B(n_400),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_612),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_605),
.A2(n_400),
.B(n_458),
.Y(n_687)
);

NAND2x1p5_ASAP7_75t_L g688 ( 
.A(n_609),
.B(n_458),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_633),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_620),
.A2(n_458),
.B(n_400),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_614),
.A2(n_348),
.B(n_43),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_622),
.A2(n_348),
.B(n_44),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_629),
.B(n_17),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_613),
.B(n_41),
.Y(n_694)
);

AO31x2_ASAP7_75t_L g695 ( 
.A1(n_614),
.A2(n_18),
.A3(n_19),
.B(n_20),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_626),
.B(n_48),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_609),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_643),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_600),
.A2(n_348),
.B1(n_19),
.B2(n_21),
.Y(n_699)
);

AO221x2_ASAP7_75t_L g700 ( 
.A1(n_644),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.C(n_23),
.Y(n_700)
);

NAND2x1p5_ASAP7_75t_L g701 ( 
.A(n_616),
.B(n_49),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_649),
.B(n_22),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_636),
.Y(n_703)
);

AOI21x1_ASAP7_75t_L g704 ( 
.A1(n_637),
.A2(n_118),
.B(n_205),
.Y(n_704)
);

BUFx12f_ASAP7_75t_L g705 ( 
.A(n_638),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_686),
.B(n_619),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_661),
.Y(n_707)
);

OAI21xp33_ASAP7_75t_L g708 ( 
.A1(n_699),
.A2(n_644),
.B(n_632),
.Y(n_708)
);

O2A1O1Ixp5_ASAP7_75t_L g709 ( 
.A1(n_691),
.A2(n_628),
.B(n_640),
.C(n_641),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_669),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_653),
.A2(n_642),
.B(n_647),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_652),
.A2(n_648),
.B(n_645),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_675),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_674),
.A2(n_648),
.B(n_645),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_687),
.A2(n_648),
.B(n_645),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_SL g716 ( 
.A1(n_679),
.A2(n_630),
.B(n_641),
.C(n_650),
.Y(n_716)
);

O2A1O1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_676),
.A2(n_638),
.B(n_640),
.C(n_627),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_656),
.Y(n_718)
);

BUFx10_ASAP7_75t_L g719 ( 
.A(n_696),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_663),
.A2(n_638),
.B(n_616),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_671),
.A2(n_616),
.B(n_646),
.Y(n_721)
);

OAI22x1_ASAP7_75t_L g722 ( 
.A1(n_666),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_SL g723 ( 
.A(n_660),
.B(n_24),
.Y(n_723)
);

BUFx12f_ASAP7_75t_L g724 ( 
.A(n_659),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_667),
.A2(n_206),
.B(n_119),
.Y(n_725)
);

NAND3x1_ASAP7_75t_L g726 ( 
.A(n_693),
.B(n_26),
.C(n_27),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_SL g727 ( 
.A1(n_694),
.A2(n_120),
.B(n_197),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_662),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_685),
.A2(n_116),
.B(n_196),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_696),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_658),
.A2(n_28),
.B(n_29),
.C(n_50),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_667),
.B(n_51),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_672),
.B(n_203),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_672),
.B(n_52),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_673),
.Y(n_735)
);

AO32x2_ASAP7_75t_L g736 ( 
.A1(n_654),
.A2(n_53),
.A3(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_736)
);

CKINVDCx16_ASAP7_75t_R g737 ( 
.A(n_705),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_658),
.A2(n_57),
.B(n_58),
.Y(n_738)
);

OAI21xp5_ASAP7_75t_L g739 ( 
.A1(n_665),
.A2(n_59),
.B(n_63),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_700),
.B(n_64),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_677),
.A2(n_65),
.B(n_68),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_698),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_677),
.A2(n_69),
.B(n_70),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_681),
.A2(n_72),
.B(n_73),
.Y(n_744)
);

AO21x1_ASAP7_75t_L g745 ( 
.A1(n_702),
.A2(n_74),
.B(n_75),
.Y(n_745)
);

AOI221x1_ASAP7_75t_L g746 ( 
.A1(n_690),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.C(n_80),
.Y(n_746)
);

AOI221x1_ASAP7_75t_L g747 ( 
.A1(n_681),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.C(n_85),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_683),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_689),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_700),
.B(n_86),
.C(n_89),
.Y(n_750)
);

AOI31xp67_ASAP7_75t_L g751 ( 
.A1(n_657),
.A2(n_92),
.A3(n_93),
.B(n_94),
.Y(n_751)
);

AOI21x1_ASAP7_75t_L g752 ( 
.A1(n_704),
.A2(n_95),
.B(n_96),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_698),
.B(n_194),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_655),
.A2(n_98),
.B(n_99),
.Y(n_754)
);

AO31x2_ASAP7_75t_L g755 ( 
.A1(n_703),
.A2(n_100),
.A3(n_101),
.B(n_102),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_694),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_680),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_703),
.Y(n_758)
);

BUFx10_ASAP7_75t_L g759 ( 
.A(n_697),
.Y(n_759)
);

AO32x2_ASAP7_75t_L g760 ( 
.A1(n_654),
.A2(n_108),
.A3(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_692),
.A2(n_113),
.B(n_114),
.C(n_115),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_664),
.A2(n_123),
.B(n_125),
.Y(n_762)
);

AO22x2_ASAP7_75t_L g763 ( 
.A1(n_657),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_670),
.Y(n_764)
);

AO31x2_ASAP7_75t_L g765 ( 
.A1(n_668),
.A2(n_131),
.A3(n_133),
.B(n_134),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_682),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_684),
.A2(n_137),
.B(n_139),
.Y(n_767)
);

INVx3_ASAP7_75t_SL g768 ( 
.A(n_737),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_763),
.A2(n_680),
.B1(n_701),
.B2(n_668),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_758),
.Y(n_770)
);

INVx4_ASAP7_75t_SL g771 ( 
.A(n_724),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_708),
.A2(n_680),
.B1(n_678),
.B2(n_688),
.Y(n_772)
);

INVx6_ASAP7_75t_L g773 ( 
.A(n_719),
.Y(n_773)
);

INVx6_ASAP7_75t_L g774 ( 
.A(n_719),
.Y(n_774)
);

INVx5_ASAP7_75t_L g775 ( 
.A(n_759),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_738),
.A2(n_668),
.B(n_678),
.Y(n_776)
);

BUFx4f_ASAP7_75t_L g777 ( 
.A(n_756),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_742),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_764),
.B(n_668),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_735),
.Y(n_780)
);

INVx6_ASAP7_75t_L g781 ( 
.A(n_730),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_710),
.Y(n_782)
);

BUFx5_ASAP7_75t_L g783 ( 
.A(n_730),
.Y(n_783)
);

INVx6_ASAP7_75t_L g784 ( 
.A(n_759),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_709),
.A2(n_695),
.B(n_141),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_713),
.Y(n_786)
);

CKINVDCx11_ASAP7_75t_R g787 ( 
.A(n_748),
.Y(n_787)
);

BUFx8_ASAP7_75t_L g788 ( 
.A(n_740),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_706),
.A2(n_695),
.B1(n_142),
.B2(n_143),
.Y(n_789)
);

AOI21xp33_ASAP7_75t_L g790 ( 
.A1(n_717),
.A2(n_695),
.B(n_144),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_750),
.A2(n_140),
.B1(n_145),
.B2(n_146),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_763),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_749),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_707),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_718),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_SL g796 ( 
.A1(n_728),
.A2(n_150),
.B1(n_151),
.B2(n_154),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_766),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_731),
.A2(n_155),
.B1(n_157),
.B2(n_159),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_739),
.A2(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_753),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_711),
.B(n_167),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_732),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_755),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_767),
.Y(n_804)
);

CKINVDCx11_ASAP7_75t_R g805 ( 
.A(n_757),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_733),
.Y(n_806)
);

BUFx8_ASAP7_75t_L g807 ( 
.A(n_736),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_755),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_722),
.A2(n_169),
.B1(n_171),
.B2(n_175),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_720),
.Y(n_810)
);

BUFx8_ASAP7_75t_L g811 ( 
.A(n_736),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_723),
.A2(n_176),
.B1(n_178),
.B2(n_180),
.Y(n_812)
);

INVx6_ASAP7_75t_L g813 ( 
.A(n_727),
.Y(n_813)
);

INVx6_ASAP7_75t_L g814 ( 
.A(n_726),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_745),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_734),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_765),
.Y(n_817)
);

CKINVDCx6p67_ASAP7_75t_R g818 ( 
.A(n_736),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_762),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_725),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_820)
);

OAI22xp33_ASAP7_75t_L g821 ( 
.A1(n_747),
.A2(n_746),
.B1(n_744),
.B2(n_743),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_765),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_765),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_712),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_741),
.A2(n_714),
.B1(n_715),
.B2(n_721),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_770),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_807),
.Y(n_827)
);

OA21x2_ASAP7_75t_L g828 ( 
.A1(n_785),
.A2(n_729),
.B(n_754),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_818),
.B(n_760),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_810),
.B(n_760),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_824),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_811),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_778),
.B(n_761),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_803),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_808),
.Y(n_835)
);

BUFx12f_ASAP7_75t_L g836 ( 
.A(n_787),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_782),
.Y(n_837)
);

AO21x2_ASAP7_75t_L g838 ( 
.A1(n_821),
.A2(n_752),
.B(n_716),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_804),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_794),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_817),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_798),
.A2(n_751),
.B(n_760),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_822),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_823),
.B(n_802),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_804),
.Y(n_845)
);

AO21x2_ASAP7_75t_L g846 ( 
.A1(n_790),
.A2(n_776),
.B(n_789),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_773),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_816),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_779),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_769),
.B(n_800),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_793),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_786),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_786),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_783),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_783),
.Y(n_855)
);

OAI21xp33_ASAP7_75t_SL g856 ( 
.A1(n_792),
.A2(n_815),
.B(n_819),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_783),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_783),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_795),
.B(n_806),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_773),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_774),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_797),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_801),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_825),
.Y(n_864)
);

OAI21x1_ASAP7_75t_L g865 ( 
.A1(n_772),
.A2(n_820),
.B(n_791),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_774),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_775),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_781),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_814),
.B(n_809),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_775),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_781),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_826),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_868),
.B(n_768),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_837),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_829),
.B(n_780),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_856),
.A2(n_814),
.B1(n_788),
.B2(n_813),
.Y(n_876)
);

OA21x2_ASAP7_75t_L g877 ( 
.A1(n_842),
.A2(n_812),
.B(n_799),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_843),
.B(n_771),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_851),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_849),
.B(n_813),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_826),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_829),
.B(n_771),
.Y(n_882)
);

AO21x2_ASAP7_75t_L g883 ( 
.A1(n_842),
.A2(n_805),
.B(n_796),
.Y(n_883)
);

AND2x4_ASAP7_75t_SL g884 ( 
.A(n_866),
.B(n_777),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_837),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_843),
.Y(n_886)
);

INVxp67_ASAP7_75t_SL g887 ( 
.A(n_851),
.Y(n_887)
);

OR2x6_ASAP7_75t_L g888 ( 
.A(n_829),
.B(n_784),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_836),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_849),
.B(n_784),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_834),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_834),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_868),
.B(n_859),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_848),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_843),
.B(n_855),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_862),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_848),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_839),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_844),
.B(n_835),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_839),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_859),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_835),
.Y(n_902)
);

BUFx2_ASAP7_75t_SL g903 ( 
.A(n_847),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_835),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_895),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_876),
.A2(n_827),
.B1(n_832),
.B2(n_869),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_902),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_872),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_902),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_888),
.B(n_832),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_893),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_904),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_888),
.B(n_827),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_895),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_904),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_888),
.B(n_827),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_901),
.B(n_840),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_891),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_888),
.B(n_850),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_889),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_891),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_874),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_875),
.B(n_850),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_892),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_895),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_875),
.B(n_850),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_899),
.B(n_840),
.Y(n_927)
);

INVxp33_ASAP7_75t_L g928 ( 
.A(n_906),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_919),
.B(n_923),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_920),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_919),
.B(n_882),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_923),
.B(n_882),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_926),
.B(n_878),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_926),
.B(n_878),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_905),
.B(n_878),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_918),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_920),
.Y(n_937)
);

NOR2xp67_ASAP7_75t_L g938 ( 
.A(n_905),
.B(n_836),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_910),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_905),
.B(n_886),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_914),
.B(n_886),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_927),
.B(n_899),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_918),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_SL g944 ( 
.A(n_913),
.B(n_836),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_931),
.B(n_910),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_936),
.B(n_908),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_936),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_937),
.B(n_911),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_930),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_931),
.B(n_913),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_943),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_930),
.Y(n_952)
);

NAND2xp33_ASAP7_75t_SL g953 ( 
.A(n_928),
.B(n_916),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_938),
.B(n_916),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_929),
.B(n_914),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_943),
.B(n_921),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_929),
.B(n_921),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_947),
.Y(n_958)
);

NOR2xp67_ASAP7_75t_L g959 ( 
.A(n_949),
.B(n_939),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_950),
.B(n_938),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_953),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_951),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_948),
.B(n_939),
.Y(n_963)
);

OAI21xp33_ASAP7_75t_SL g964 ( 
.A1(n_945),
.A2(n_932),
.B(n_933),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_949),
.B(n_957),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_957),
.B(n_942),
.Y(n_966)
);

OAI22xp33_ASAP7_75t_L g967 ( 
.A1(n_961),
.A2(n_959),
.B1(n_944),
.B2(n_952),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_965),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_965),
.B(n_937),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_963),
.B(n_932),
.Y(n_970)
);

AO221x2_ASAP7_75t_L g971 ( 
.A1(n_964),
.A2(n_856),
.B1(n_889),
.B2(n_890),
.C(n_917),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_SL g972 ( 
.A(n_960),
.B(n_954),
.Y(n_972)
);

OAI22xp33_ASAP7_75t_L g973 ( 
.A1(n_966),
.A2(n_877),
.B1(n_954),
.B2(n_942),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_972),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_969),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_968),
.B(n_958),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_970),
.B(n_962),
.Y(n_977)
);

AOI31xp33_ASAP7_75t_L g978 ( 
.A1(n_967),
.A2(n_867),
.A3(n_870),
.B(n_873),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_971),
.B(n_955),
.Y(n_979)
);

NOR2x1_ASAP7_75t_L g980 ( 
.A(n_973),
.B(n_956),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_972),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_969),
.B(n_946),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_968),
.B(n_933),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_975),
.B(n_934),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_974),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_977),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_981),
.A2(n_935),
.B1(n_934),
.B2(n_946),
.Y(n_987)
);

NAND2xp33_ASAP7_75t_L g988 ( 
.A(n_980),
.B(n_870),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_978),
.A2(n_935),
.B1(n_956),
.B2(n_867),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_979),
.A2(n_883),
.B1(n_877),
.B2(n_846),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_976),
.A2(n_869),
.B(n_865),
.C(n_884),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_988),
.A2(n_983),
.B1(n_883),
.B2(n_982),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_985),
.B(n_927),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_SL g994 ( 
.A1(n_990),
.A2(n_869),
.B(n_884),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_989),
.A2(n_883),
.B(n_847),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_986),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_984),
.B(n_941),
.Y(n_997)
);

OAI22xp33_ASAP7_75t_L g998 ( 
.A1(n_987),
.A2(n_877),
.B1(n_847),
.B2(n_880),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_994),
.A2(n_991),
.B1(n_871),
.B2(n_860),
.Y(n_999)
);

OAI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_993),
.A2(n_877),
.B1(n_860),
.B2(n_871),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_992),
.A2(n_846),
.B1(n_864),
.B2(n_833),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_995),
.A2(n_865),
.B(n_871),
.C(n_861),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_996),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_1003),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_999),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_1002),
.B(n_997),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_1000),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_1001),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_1003),
.Y(n_1009)
);

NAND4xp75_ASAP7_75t_L g1010 ( 
.A(n_1004),
.B(n_998),
.C(n_941),
.D(n_940),
.Y(n_1010)
);

NOR2x1_ASAP7_75t_L g1011 ( 
.A(n_1007),
.B(n_871),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1009),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_L g1013 ( 
.A(n_1005),
.B(n_860),
.C(n_861),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1008),
.A2(n_861),
.B1(n_860),
.B2(n_866),
.Y(n_1014)
);

NOR3xp33_ASAP7_75t_SL g1015 ( 
.A(n_1006),
.B(n_864),
.C(n_852),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1012),
.B(n_1009),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_L g1017 ( 
.A(n_1011),
.B(n_1013),
.C(n_1014),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_1015),
.A2(n_866),
.B(n_861),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_SL g1019 ( 
.A(n_1010),
.B(n_903),
.Y(n_1019)
);

NAND4xp25_ASAP7_75t_SL g1020 ( 
.A(n_1017),
.B(n_940),
.C(n_852),
.D(n_862),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1016),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_SL g1022 ( 
.A(n_1018),
.B(n_887),
.C(n_924),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1019),
.B(n_924),
.Y(n_1023)
);

NOR2x1_ASAP7_75t_L g1024 ( 
.A(n_1016),
.B(n_903),
.Y(n_1024)
);

NAND4xp25_ASAP7_75t_L g1025 ( 
.A(n_1017),
.B(n_833),
.C(n_862),
.D(n_853),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_1016),
.B(n_853),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1016),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1021),
.A2(n_846),
.B(n_863),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1027),
.Y(n_1029)
);

AO22x2_ASAP7_75t_L g1030 ( 
.A1(n_1023),
.A2(n_925),
.B1(n_914),
.B2(n_853),
.Y(n_1030)
);

AND3x2_ASAP7_75t_L g1031 ( 
.A(n_1026),
.B(n_879),
.C(n_896),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1024),
.Y(n_1032)
);

NOR2xp67_ASAP7_75t_SL g1033 ( 
.A(n_1025),
.B(n_1020),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1022),
.B(n_925),
.Y(n_1034)
);

AND4x1_ASAP7_75t_L g1035 ( 
.A(n_1021),
.B(n_844),
.C(n_881),
.D(n_872),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_1026),
.Y(n_1036)
);

XNOR2xp5_ASAP7_75t_L g1037 ( 
.A(n_1021),
.B(n_865),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_1032),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1033),
.B(n_925),
.Y(n_1039)
);

AND3x4_ASAP7_75t_L g1040 ( 
.A(n_1035),
.B(n_858),
.C(n_857),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_L g1041 ( 
.A(n_1029),
.B(n_898),
.Y(n_1041)
);

NAND4xp25_ASAP7_75t_L g1042 ( 
.A(n_1036),
.B(n_898),
.C(n_900),
.D(n_863),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1034),
.A2(n_898),
.B1(n_900),
.B2(n_912),
.Y(n_1043)
);

NAND3x1_ASAP7_75t_SL g1044 ( 
.A(n_1031),
.B(n_830),
.C(n_844),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_1037),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_1028),
.B(n_900),
.Y(n_1046)
);

AND4x1_ASAP7_75t_L g1047 ( 
.A(n_1030),
.B(n_881),
.C(n_915),
.D(n_912),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1032),
.B(n_915),
.Y(n_1048)
);

AND3x4_ASAP7_75t_L g1049 ( 
.A(n_1032),
.B(n_855),
.C(n_858),
.Y(n_1049)
);

AND3x4_ASAP7_75t_L g1050 ( 
.A(n_1032),
.B(n_855),
.C(n_858),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_1038),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_1049),
.Y(n_1052)
);

XNOR2x1_ASAP7_75t_L g1053 ( 
.A(n_1045),
.B(n_863),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_1050),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1041),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_1039),
.A2(n_909),
.B1(n_907),
.B2(n_846),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1048),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1040),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1051),
.A2(n_1058),
.B1(n_1052),
.B2(n_1054),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1055),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_1057),
.A2(n_1043),
.B1(n_1046),
.B2(n_1044),
.Y(n_1061)
);

OAI22x1_ASAP7_75t_L g1062 ( 
.A1(n_1053),
.A2(n_1047),
.B1(n_1042),
.B2(n_857),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1056),
.A2(n_909),
.B1(n_907),
.B2(n_922),
.Y(n_1063)
);

AO22x1_ASAP7_75t_L g1064 ( 
.A1(n_1051),
.A2(n_857),
.B1(n_854),
.B2(n_845),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1051),
.A2(n_922),
.B1(n_854),
.B2(n_845),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1060),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1062),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1059),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1068),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1069),
.B(n_1066),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1070),
.A2(n_1067),
.B1(n_1061),
.B2(n_1065),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1071),
.A2(n_1063),
.B1(n_1064),
.B2(n_854),
.Y(n_1072)
);

OAI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1071),
.A2(n_839),
.B1(n_845),
.B2(n_892),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1072),
.A2(n_1073),
.B(n_838),
.Y(n_1074)
);

OA21x2_ASAP7_75t_L g1075 ( 
.A1(n_1072),
.A2(n_848),
.B(n_897),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1074),
.A2(n_828),
.B(n_831),
.Y(n_1076)
);

AO21x2_ASAP7_75t_L g1077 ( 
.A1(n_1075),
.A2(n_838),
.B(n_885),
.Y(n_1077)
);

AOI221xp5_ASAP7_75t_L g1078 ( 
.A1(n_1076),
.A2(n_1077),
.B1(n_839),
.B2(n_841),
.C(n_894),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1076),
.A2(n_839),
.B1(n_838),
.B2(n_841),
.Y(n_1079)
);

AOI211xp5_ASAP7_75t_L g1080 ( 
.A1(n_1078),
.A2(n_1079),
.B(n_839),
.C(n_830),
.Y(n_1080)
);


endmodule