module fake_jpeg_4884_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_31),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx9p33_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_16),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_27),
.B1(n_25),
.B2(n_28),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_53),
.B1(n_16),
.B2(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_27),
.B1(n_25),
.B2(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_60),
.B1(n_63),
.B2(n_68),
.Y(n_97)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_27),
.B1(n_19),
.B2(n_28),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_64),
.B1(n_33),
.B2(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_19),
.B1(n_25),
.B2(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_24),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_19),
.B1(n_25),
.B2(n_30),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_34),
.A2(n_19),
.B1(n_24),
.B2(n_26),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_34),
.A2(n_19),
.B1(n_32),
.B2(n_16),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_90),
.B1(n_69),
.B2(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_40),
.B1(n_24),
.B2(n_33),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_43),
.B1(n_35),
.B2(n_40),
.Y(n_77)
);

AO22x1_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_66),
.B1(n_56),
.B2(n_55),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_88),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_43),
.B(n_17),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_91),
.B(n_26),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_40),
.C(n_37),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_47),
.B(n_33),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_37),
.C(n_36),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_96),
.Y(n_112)
);

AOI32xp33_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_36),
.A3(n_29),
.B1(n_22),
.B2(n_21),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_71),
.C(n_62),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_49),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

AO22x1_ASAP7_75t_SL g137 ( 
.A1(n_104),
.A2(n_118),
.B1(n_96),
.B2(n_74),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_116),
.B1(n_81),
.B2(n_78),
.Y(n_125)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_48),
.B1(n_58),
.B2(n_52),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_113),
.B1(n_117),
.B2(n_120),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_66),
.B1(n_60),
.B2(n_63),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_48),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_115),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_68),
.B1(n_59),
.B2(n_73),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_59),
.B1(n_67),
.B2(n_50),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_92),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_70),
.B1(n_33),
.B2(n_67),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_65),
.C(n_54),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_81),
.C(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_131),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_138),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_78),
.B1(n_85),
.B2(n_94),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_130),
.A2(n_133),
.B1(n_139),
.B2(n_144),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_86),
.B1(n_54),
.B2(n_79),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_79),
.B1(n_92),
.B2(n_82),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_104),
.B1(n_102),
.B2(n_33),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_82),
.B1(n_80),
.B2(n_74),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_26),
.B(n_32),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_142),
.B(n_118),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_32),
.B(n_23),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_74),
.C(n_29),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_110),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_117),
.B1(n_114),
.B2(n_99),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_146),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_32),
.C(n_22),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_120),
.Y(n_154)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_174),
.C(n_128),
.Y(n_187)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_156),
.B(n_159),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_161),
.B(n_168),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_124),
.B(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_100),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_144),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_104),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_109),
.B(n_98),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_169),
.A2(n_171),
.B(n_29),
.Y(n_207)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_177),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_122),
.B(n_104),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_136),
.B1(n_141),
.B2(n_149),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_107),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_107),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_145),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_182),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_168),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_186),
.A2(n_202),
.B1(n_156),
.B2(n_181),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_189),
.C(n_204),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_154),
.C(n_174),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_198),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_148),
.B1(n_153),
.B2(n_136),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_209),
.Y(n_211)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_157),
.B(n_143),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_199),
.A2(n_158),
.B(n_146),
.Y(n_228)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_208),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_153),
.B1(n_102),
.B2(n_135),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_134),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_132),
.C(n_127),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_176),
.C(n_169),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_161),
.B(n_176),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_162),
.A2(n_159),
.B1(n_164),
.B2(n_160),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_210),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_195),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_227),
.B(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_224),
.B(n_200),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_199),
.B(n_166),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_221),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_167),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_226),
.C(n_235),
.Y(n_244)
);

XOR2x2_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_168),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_189),
.C(n_187),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_206),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_197),
.A2(n_127),
.B1(n_134),
.B2(n_108),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_196),
.B1(n_197),
.B2(n_194),
.Y(n_243)
);

OAI22x1_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_108),
.B1(n_22),
.B2(n_21),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_236),
.B1(n_21),
.B2(n_20),
.Y(n_257)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_22),
.C(n_21),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_203),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_214),
.A2(n_191),
.B1(n_193),
.B2(n_188),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_255),
.B(n_256),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_188),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_193),
.C(n_183),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_20),
.C(n_17),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_229),
.B(n_183),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_191),
.B1(n_207),
.B2(n_194),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_258),
.B1(n_231),
.B2(n_235),
.Y(n_274)
);

FAx1_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_22),
.CI(n_21),
.CON(n_255),
.SN(n_255)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_228),
.A2(n_1),
.B(n_2),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_259),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_215),
.A2(n_20),
.B1(n_17),
.B2(n_3),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_216),
.B1(n_234),
.B2(n_211),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_260),
.A2(n_255),
.B1(n_258),
.B2(n_17),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_SL g262 ( 
.A(n_242),
.B(n_220),
.C(n_217),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_274),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_241),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_263),
.B(n_267),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_225),
.B(n_232),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_276),
.B1(n_260),
.B2(n_265),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_249),
.B(n_219),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_272),
.C(n_278),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_212),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_SL g269 ( 
.A(n_255),
.B(n_227),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_230),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_218),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_277),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_237),
.A2(n_226),
.B1(n_213),
.B2(n_20),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_20),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_250),
.C(n_244),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_279),
.A2(n_282),
.B(n_284),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_13),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_244),
.C(n_254),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_252),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_293),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_245),
.C(n_239),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_243),
.C(n_253),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_14),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_1),
.B(n_3),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_289),
.B1(n_270),
.B2(n_261),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_17),
.C(n_2),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_11),
.B(n_10),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_15),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_287),
.A2(n_269),
.B(n_274),
.C(n_270),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_302),
.B1(n_303),
.B2(n_306),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_268),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_298),
.B(n_300),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_294),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_291),
.A2(n_13),
.B(n_12),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_9),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_292),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_308),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_285),
.C(n_279),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_1),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_318),
.C(n_314),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_SL g312 ( 
.A(n_301),
.B(n_294),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_314),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_1),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_316),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_9),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_319),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_298),
.A2(n_297),
.B(n_304),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_3),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_324),
.Y(n_329)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_311),
.A2(n_303),
.B(n_4),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_3),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_5),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_4),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_5),
.C(n_6),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_SL g328 ( 
.A1(n_322),
.A2(n_323),
.B(n_321),
.C(n_8),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_328),
.A2(n_330),
.B(n_332),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_5),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_7),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_333),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_SL g336 ( 
.A(n_334),
.B(n_329),
.C(n_331),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_335),
.Y(n_337)
);

OAI221xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_322),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_7),
.Y(n_339)
);


endmodule