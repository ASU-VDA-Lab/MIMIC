module real_aes_11812_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_1612;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_602;
wire n_402;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1596;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1595;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_1584;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AO221x1_ASAP7_75t_L g1333 ( .A1(n_0), .A2(n_165), .B1(n_1258), .B2(n_1324), .C(n_1334), .Y(n_1333) );
CKINVDCx5p33_ASAP7_75t_R g1490 ( .A(n_1), .Y(n_1490) );
CKINVDCx5p33_ASAP7_75t_R g1581 ( .A(n_2), .Y(n_1581) );
AO22x2_ASAP7_75t_L g678 ( .A1(n_3), .A2(n_679), .B1(n_733), .B2(n_734), .Y(n_678) );
INVxp67_ASAP7_75t_L g733 ( .A(n_3), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_4), .A2(n_233), .B1(n_319), .B2(n_327), .Y(n_318) );
INVx1_ASAP7_75t_L g441 ( .A(n_4), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_5), .A2(n_247), .B1(n_723), .B2(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g857 ( .A(n_5), .Y(n_857) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_6), .Y(n_296) );
INVx1_ASAP7_75t_L g485 ( .A(n_6), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_6), .B(n_205), .Y(n_527) );
AND2x2_ASAP7_75t_L g531 ( .A(n_6), .B(n_323), .Y(n_531) );
OAI211xp5_ASAP7_75t_L g1470 ( .A1(n_7), .A2(n_1471), .B(n_1477), .C(n_1523), .Y(n_1470) );
AOI22xp5_ASAP7_75t_L g1278 ( .A1(n_8), .A2(n_126), .B1(n_1258), .B2(n_1262), .Y(n_1278) );
CKINVDCx5p33_ASAP7_75t_R g1507 ( .A(n_9), .Y(n_1507) );
OAI22xp33_ASAP7_75t_L g1588 ( .A1(n_10), .A2(n_188), .B1(n_569), .B2(n_578), .Y(n_1588) );
INVx1_ASAP7_75t_L g1605 ( .A(n_10), .Y(n_1605) );
INVx1_ASAP7_75t_L g628 ( .A(n_11), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_11), .A2(n_146), .B1(n_664), .B2(n_667), .Y(n_663) );
INVx1_ASAP7_75t_L g973 ( .A(n_12), .Y(n_973) );
OAI221xp5_ASAP7_75t_L g988 ( .A1(n_12), .A2(n_540), .B1(n_775), .B2(n_989), .C(n_992), .Y(n_988) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_13), .Y(n_359) );
INVx1_ASAP7_75t_L g811 ( .A(n_14), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_14), .A2(n_80), .B1(n_854), .B2(n_855), .Y(n_853) );
XNOR2x2_ASAP7_75t_L g488 ( .A(n_15), .B(n_489), .Y(n_488) );
AOI21xp33_ASAP7_75t_L g512 ( .A1(n_16), .A2(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g592 ( .A(n_16), .Y(n_592) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_17), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_17), .A2(n_257), .B1(n_648), .B2(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g999 ( .A(n_18), .Y(n_999) );
OAI22xp33_ASAP7_75t_L g1014 ( .A1(n_18), .A2(n_28), .B1(n_1015), .B2(n_1017), .Y(n_1014) );
XNOR2xp5_ASAP7_75t_L g867 ( .A(n_19), .B(n_868), .Y(n_867) );
AO22x2_ASAP7_75t_L g1020 ( .A1(n_20), .A2(n_1021), .B1(n_1022), .B2(n_1074), .Y(n_1020) );
INVxp67_ASAP7_75t_SL g1021 ( .A(n_20), .Y(n_1021) );
AO221x2_ASAP7_75t_L g1321 ( .A1(n_20), .A2(n_180), .B1(n_1322), .B2(n_1324), .C(n_1326), .Y(n_1321) );
OAI22xp5_ASAP7_75t_L g371 ( .A1(n_21), .A2(n_47), .B1(n_372), .B2(n_380), .Y(n_371) );
INVx1_ASAP7_75t_L g473 ( .A(n_21), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_22), .A2(n_217), .B1(n_757), .B2(n_824), .C(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g1157 ( .A(n_22), .Y(n_1157) );
INVx2_ASAP7_75t_L g366 ( .A(n_23), .Y(n_366) );
OR2x2_ASAP7_75t_L g591 ( .A(n_23), .B(n_576), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_24), .A2(n_169), .B1(n_529), .B2(n_535), .Y(n_528) );
INVx1_ASAP7_75t_L g567 ( .A(n_24), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_25), .Y(n_516) );
AOI22xp33_ASAP7_75t_SL g640 ( .A1(n_26), .A2(n_85), .B1(n_637), .B2(n_641), .Y(n_640) );
INVxp33_ASAP7_75t_L g674 ( .A(n_26), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_27), .A2(n_145), .B1(n_599), .B2(n_602), .Y(n_1091) );
INVx1_ASAP7_75t_L g1113 ( .A(n_27), .Y(n_1113) );
AOI221xp5_ASAP7_75t_L g1002 ( .A1(n_28), .A2(n_135), .B1(n_513), .B2(n_514), .C(n_624), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_29), .A2(n_108), .B1(n_823), .B2(n_824), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_29), .A2(n_108), .B1(n_839), .B2(n_841), .Y(n_838) );
OAI221xp5_ASAP7_75t_L g1492 ( .A1(n_30), .A2(n_219), .B1(n_1493), .B2(n_1497), .C(n_1499), .Y(n_1492) );
INVx1_ASAP7_75t_L g1548 ( .A(n_30), .Y(n_1548) );
BUFx2_ASAP7_75t_L g314 ( .A(n_31), .Y(n_314) );
BUFx2_ASAP7_75t_L g412 ( .A(n_31), .Y(n_412) );
INVx1_ASAP7_75t_L g483 ( .A(n_31), .Y(n_483) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_31), .B(n_527), .Y(n_1475) );
AOI22xp33_ASAP7_75t_SL g937 ( .A1(n_32), .A2(n_196), .B1(n_826), .B2(n_889), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_32), .A2(n_196), .B1(n_942), .B2(n_943), .Y(n_941) );
INVx1_ASAP7_75t_L g880 ( .A(n_33), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_33), .A2(n_195), .B1(n_637), .B2(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g621 ( .A(n_34), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_34), .A2(n_68), .B1(n_654), .B2(n_655), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_35), .A2(n_241), .B1(n_667), .B2(n_689), .C(n_690), .Y(n_688) );
INVx1_ASAP7_75t_L g700 ( .A(n_35), .Y(n_700) );
INVx1_ASAP7_75t_L g1586 ( .A(n_36), .Y(n_1586) );
OAI22xp5_ASAP7_75t_L g1592 ( .A1(n_36), .A2(n_77), .B1(n_529), .B2(n_535), .Y(n_1592) );
OAI22xp33_ASAP7_75t_L g931 ( .A1(n_37), .A2(n_65), .B1(n_297), .B2(n_619), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_37), .A2(n_177), .B1(n_947), .B2(n_948), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g1149 ( .A1(n_38), .A2(n_61), .B1(n_451), .B2(n_622), .C(n_1150), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_38), .A2(n_61), .B1(n_919), .B2(n_1176), .Y(n_1175) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_39), .A2(n_45), .B1(n_540), .B2(n_542), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g560 ( .A1(n_39), .A2(n_45), .B1(n_549), .B2(n_561), .C(n_563), .Y(n_560) );
OAI22xp33_ASAP7_75t_L g983 ( .A1(n_40), .A2(n_59), .B1(n_569), .B2(n_578), .Y(n_983) );
INVx1_ASAP7_75t_L g1007 ( .A(n_40), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_41), .A2(n_71), .B1(n_1059), .B2(n_1062), .Y(n_1061) );
INVxp67_ASAP7_75t_SL g1067 ( .A(n_41), .Y(n_1067) );
INVx1_ASAP7_75t_L g1216 ( .A(n_42), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g1238 ( .A1(n_42), .A2(n_63), .B1(n_1015), .B2(n_1017), .Y(n_1238) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_43), .A2(n_234), .B1(n_549), .B2(n_651), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g895 ( .A1(n_43), .A2(n_234), .B1(n_634), .B2(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g1602 ( .A(n_44), .Y(n_1602) );
OAI22xp33_ASAP7_75t_L g1608 ( .A1(n_44), .A2(n_232), .B1(n_602), .B2(n_1013), .Y(n_1608) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_46), .Y(n_495) );
INVx1_ASAP7_75t_L g351 ( .A(n_47), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_48), .A2(n_86), .B1(n_637), .B2(n_639), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_48), .A2(n_86), .B1(n_648), .B2(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g817 ( .A(n_49), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_49), .A2(n_258), .B1(n_831), .B2(n_834), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_50), .Y(n_420) );
INVx1_ASAP7_75t_L g1335 ( .A(n_51), .Y(n_1335) );
AOI222xp33_ASAP7_75t_L g1465 ( .A1(n_51), .A2(n_1466), .B1(n_1564), .B2(n_1568), .C1(n_1611), .C2(n_1613), .Y(n_1465) );
OAI22xp5_ASAP7_75t_L g1469 ( .A1(n_51), .A2(n_1335), .B1(n_1470), .B2(n_1563), .Y(n_1469) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_52), .A2(n_239), .B1(n_667), .B2(n_874), .Y(n_873) );
OAI22xp33_ASAP7_75t_L g906 ( .A1(n_52), .A2(n_239), .B1(n_627), .B2(n_907), .Y(n_906) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_53), .A2(n_78), .B1(n_451), .B2(n_517), .C(n_624), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_53), .A2(n_78), .B1(n_654), .B2(n_782), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_54), .A2(n_171), .B1(n_1117), .B2(n_1118), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_54), .A2(n_171), .B1(n_1129), .B2(n_1130), .Y(n_1128) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_55), .Y(n_498) );
INVx1_ASAP7_75t_L g1086 ( .A(n_56), .Y(n_1086) );
INVx1_ASAP7_75t_L g976 ( .A(n_57), .Y(n_976) );
OAI211xp5_ASAP7_75t_L g996 ( .A1(n_57), .A2(n_542), .B(n_997), .C(n_1003), .Y(n_996) );
INVx1_ASAP7_75t_L g1590 ( .A(n_58), .Y(n_1590) );
INVx1_ASAP7_75t_L g1004 ( .A(n_59), .Y(n_1004) );
AOI221xp5_ASAP7_75t_L g1603 ( .A1(n_60), .A2(n_232), .B1(n_513), .B2(n_514), .C(n_1486), .Y(n_1603) );
OAI22xp33_ASAP7_75t_L g1609 ( .A1(n_60), .A2(n_93), .B1(n_1015), .B2(n_1017), .Y(n_1609) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_62), .A2(n_98), .B1(n_634), .B2(n_643), .Y(n_642) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_62), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g1219 ( .A1(n_63), .A2(n_73), .B1(n_634), .B2(n_643), .C(n_1220), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_64), .A2(n_152), .B1(n_848), .B2(n_950), .Y(n_1198) );
INVx1_ASAP7_75t_L g1230 ( .A(n_64), .Y(n_1230) );
OAI22xp33_ASAP7_75t_L g926 ( .A1(n_65), .A2(n_230), .B1(n_372), .B2(n_380), .Y(n_926) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_66), .A2(n_121), .B1(n_624), .B2(n_1046), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_66), .A2(n_121), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_67), .Y(n_506) );
INVxp33_ASAP7_75t_L g616 ( .A(n_68), .Y(n_616) );
AO22x2_ASAP7_75t_L g801 ( .A1(n_69), .A2(n_802), .B1(n_862), .B2(n_863), .Y(n_801) );
INVxp67_ASAP7_75t_SL g862 ( .A(n_69), .Y(n_862) );
CKINVDCx16_ASAP7_75t_R g1135 ( .A(n_70), .Y(n_1135) );
INVxp33_ASAP7_75t_L g1073 ( .A(n_71), .Y(n_1073) );
OAI221xp5_ASAP7_75t_L g1095 ( .A1(n_72), .A2(n_540), .B1(n_775), .B2(n_1096), .C(n_1100), .Y(n_1095) );
AOI22xp33_ASAP7_75t_SL g1127 ( .A1(n_72), .A2(n_210), .B1(n_846), .B2(n_945), .Y(n_1127) );
OAI22xp5_ASAP7_75t_L g1237 ( .A1(n_73), .A2(n_203), .B1(n_602), .B2(n_1013), .Y(n_1237) );
INVx1_ASAP7_75t_L g1336 ( .A(n_74), .Y(n_1336) );
INVx1_ASAP7_75t_L g1488 ( .A(n_75), .Y(n_1488) );
AOI221xp5_ASAP7_75t_L g1555 ( .A1(n_75), .A2(n_140), .B1(n_1062), .B2(n_1556), .C(n_1558), .Y(n_1555) );
INVx1_ASAP7_75t_L g698 ( .A(n_76), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_76), .A2(n_215), .B1(n_594), .B2(n_723), .Y(n_732) );
INVx1_ASAP7_75t_L g1587 ( .A(n_77), .Y(n_1587) );
INVxp67_ASAP7_75t_SL g1031 ( .A(n_79), .Y(n_1031) );
AOI22xp33_ASAP7_75t_SL g1051 ( .A1(n_79), .A2(n_116), .B1(n_824), .B2(n_1046), .Y(n_1051) );
INVx1_ASAP7_75t_L g814 ( .A(n_80), .Y(n_814) );
INVx1_ASAP7_75t_L g1516 ( .A(n_81), .Y(n_1516) );
OAI22xp5_ASAP7_75t_L g1560 ( .A1(n_81), .A2(n_250), .B1(n_1561), .B2(n_1562), .Y(n_1560) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_82), .A2(n_225), .B1(n_637), .B2(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_82), .A2(n_225), .B1(n_648), .B2(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g1099 ( .A(n_83), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_83), .A2(n_212), .B1(n_1124), .B2(n_1125), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1144 ( .A1(n_84), .A2(n_128), .B1(n_761), .B2(n_765), .Y(n_1144) );
INVx1_ASAP7_75t_L g1169 ( .A(n_84), .Y(n_1169) );
INVxp67_ASAP7_75t_SL g675 ( .A(n_85), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_87), .A2(n_130), .B1(n_362), .B2(n_925), .Y(n_924) );
AOI22xp33_ASAP7_75t_SL g938 ( .A1(n_87), .A2(n_130), .B1(n_889), .B2(n_893), .Y(n_938) );
AO221x1_ASAP7_75t_L g1286 ( .A1(n_88), .A2(n_132), .B1(n_1258), .B2(n_1262), .C(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g923 ( .A(n_89), .Y(n_923) );
OAI222xp33_ASAP7_75t_L g929 ( .A1(n_89), .A2(n_177), .B1(n_189), .B2(n_511), .C1(n_855), .C2(n_930), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_90), .A2(n_122), .B1(n_848), .B2(n_950), .Y(n_1064) );
INVxp33_ASAP7_75t_SL g1070 ( .A(n_90), .Y(n_1070) );
INVx1_ASAP7_75t_L g1328 ( .A(n_91), .Y(n_1328) );
INVx1_ASAP7_75t_L g981 ( .A(n_92), .Y(n_981) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_92), .A2(n_154), .B1(n_529), .B2(n_535), .Y(n_987) );
INVx1_ASAP7_75t_L g1600 ( .A(n_93), .Y(n_1600) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_94), .A2(n_109), .B1(n_754), .B2(n_755), .C(n_757), .Y(n_753) );
INVx1_ASAP7_75t_L g787 ( .A(n_94), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_95), .Y(n_432) );
AO221x1_ASAP7_75t_L g1280 ( .A1(n_96), .A2(n_174), .B1(n_1258), .B2(n_1262), .C(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1283 ( .A(n_97), .Y(n_1283) );
INVxp33_ASAP7_75t_L g669 ( .A(n_98), .Y(n_669) );
INVx1_ASAP7_75t_L g410 ( .A(n_99), .Y(n_410) );
INVx1_ASAP7_75t_L g576 ( .A(n_99), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_100), .A2(n_166), .B1(n_549), .B2(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g912 ( .A(n_100), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_101), .A2(n_103), .B1(n_578), .B2(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1222 ( .A(n_101), .Y(n_1222) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_102), .A2(n_142), .B1(n_885), .B2(n_886), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_102), .A2(n_142), .B1(n_893), .B2(n_894), .Y(n_892) );
INVx1_ASAP7_75t_L g1223 ( .A(n_103), .Y(n_1223) );
INVx1_ASAP7_75t_L g1146 ( .A(n_104), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g1181 ( .A1(n_104), .A2(n_105), .B1(n_844), .B2(n_943), .Y(n_1181) );
INVx1_ASAP7_75t_L g1147 ( .A(n_105), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_106), .A2(n_240), .B1(n_893), .B2(n_1049), .Y(n_1139) );
INVx1_ASAP7_75t_L g1160 ( .A(n_106), .Y(n_1160) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_107), .Y(n_429) );
INVx1_ASAP7_75t_L g789 ( .A(n_109), .Y(n_789) );
XNOR2xp5_ASAP7_75t_L g958 ( .A(n_110), .B(n_959), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_111), .A2(n_226), .B1(n_1258), .B2(n_1262), .Y(n_1257) );
INVx1_ASAP7_75t_L g767 ( .A(n_112), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_112), .A2(n_249), .B1(n_556), .B2(n_724), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_113), .A2(n_223), .B1(n_751), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_113), .A2(n_223), .B1(n_556), .B2(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g871 ( .A(n_114), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_114), .A2(n_192), .B1(n_624), .B2(n_634), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_115), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g471 ( .A(n_115), .Y(n_471) );
INVxp33_ASAP7_75t_SL g1025 ( .A(n_116), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_117), .A2(n_275), .B1(n_634), .B2(n_635), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_117), .A2(n_275), .B1(n_391), .B2(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g1143 ( .A(n_118), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_118), .A2(n_266), .B1(n_1176), .B2(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1201 ( .A(n_119), .Y(n_1201) );
OAI221xp5_ASAP7_75t_L g1224 ( .A1(n_119), .A2(n_540), .B1(n_1225), .B2(n_1227), .C(n_1234), .Y(n_1224) );
INVx1_ASAP7_75t_L g1521 ( .A(n_120), .Y(n_1521) );
OAI211xp5_ASAP7_75t_SL g1524 ( .A1(n_120), .A2(n_1525), .B(n_1529), .C(n_1538), .Y(n_1524) );
INVxp67_ASAP7_75t_SL g1071 ( .A(n_122), .Y(n_1071) );
INVx1_ASAP7_75t_L g1289 ( .A(n_123), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_124), .A2(n_255), .B1(n_826), .B2(n_827), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_124), .A2(n_255), .B1(n_723), .B2(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g288 ( .A(n_125), .Y(n_288) );
OA22x2_ASAP7_75t_L g311 ( .A1(n_126), .A2(n_312), .B1(n_486), .B2(n_487), .Y(n_311) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_126), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g877 ( .A(n_127), .Y(n_877) );
INVx1_ASAP7_75t_L g1170 ( .A(n_128), .Y(n_1170) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_129), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g1273 ( .A1(n_131), .A2(n_206), .B1(n_1264), .B2(n_1267), .Y(n_1273) );
INVx1_ASAP7_75t_L g691 ( .A(n_133), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_133), .A2(n_150), .B1(n_634), .B2(n_714), .Y(n_719) );
INVx1_ASAP7_75t_L g1288 ( .A(n_134), .Y(n_1288) );
OAI22xp33_ASAP7_75t_L g1012 ( .A1(n_135), .A2(n_163), .B1(n_602), .B2(n_1013), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_136), .A2(n_228), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g790 ( .A(n_136), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g1274 ( .A1(n_137), .A2(n_185), .B1(n_1258), .B2(n_1262), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_138), .A2(n_261), .B1(n_841), .B2(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g860 ( .A(n_138), .Y(n_860) );
AOI22xp5_ASAP7_75t_L g1263 ( .A1(n_139), .A2(n_279), .B1(n_1264), .B2(n_1267), .Y(n_1263) );
INVx1_ASAP7_75t_L g1484 ( .A(n_140), .Y(n_1484) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_141), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g568 ( .A1(n_141), .A2(n_569), .B1(n_577), .B2(n_578), .C(n_581), .Y(n_568) );
XOR2xp5_ASAP7_75t_L g1081 ( .A(n_143), .B(n_1082), .Y(n_1081) );
CKINVDCx5p33_ASAP7_75t_R g964 ( .A(n_144), .Y(n_964) );
INVx1_ASAP7_75t_L g1106 ( .A(n_145), .Y(n_1106) );
INVxp67_ASAP7_75t_SL g625 ( .A(n_146), .Y(n_625) );
INVx1_ASAP7_75t_L g707 ( .A(n_147), .Y(n_707) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_147), .A2(n_153), .B1(n_549), .B2(n_731), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_148), .A2(n_221), .B1(n_761), .B2(n_765), .Y(n_760) );
INVx1_ASAP7_75t_L g795 ( .A(n_148), .Y(n_795) );
INVx1_ASAP7_75t_L g1327 ( .A(n_149), .Y(n_1327) );
INVx1_ASAP7_75t_L g683 ( .A(n_150), .Y(n_683) );
INVx1_ASAP7_75t_L g1090 ( .A(n_151), .Y(n_1090) );
INVx1_ASAP7_75t_L g1233 ( .A(n_152), .Y(n_1233) );
INVx1_ASAP7_75t_L g702 ( .A(n_153), .Y(n_702) );
INVx1_ASAP7_75t_L g979 ( .A(n_154), .Y(n_979) );
INVx1_ASAP7_75t_L g1089 ( .A(n_155), .Y(n_1089) );
INVx1_ASAP7_75t_L g799 ( .A(n_156), .Y(n_799) );
INVx1_ASAP7_75t_L g1087 ( .A(n_157), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_158), .A2(n_242), .B1(n_901), .B2(n_902), .Y(n_900) );
INVx1_ASAP7_75t_L g909 ( .A(n_158), .Y(n_909) );
INVx1_ASAP7_75t_L g933 ( .A(n_159), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_159), .A2(n_162), .B1(n_848), .B2(n_950), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_160), .A2(n_187), .B1(n_713), .B2(n_714), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_160), .A2(n_187), .B1(n_549), .B2(n_651), .Y(n_725) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_161), .Y(n_508) );
INVx1_ASAP7_75t_L g934 ( .A(n_162), .Y(n_934) );
INVx1_ASAP7_75t_L g1001 ( .A(n_163), .Y(n_1001) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_164), .Y(n_965) );
INVx1_ASAP7_75t_L g905 ( .A(n_166), .Y(n_905) );
INVx1_ASAP7_75t_L g1101 ( .A(n_167), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_167), .A2(n_191), .B1(n_839), .B2(n_1122), .Y(n_1121) );
INVxp33_ASAP7_75t_SL g1026 ( .A(n_168), .Y(n_1026) );
AOI22xp33_ASAP7_75t_SL g1048 ( .A1(n_168), .A2(n_204), .B1(n_1041), .B2(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g564 ( .A(n_169), .Y(n_564) );
AOI22x1_ASAP7_75t_SL g913 ( .A1(n_170), .A2(n_914), .B1(n_951), .B2(n_952), .Y(n_913) );
INVx1_ASAP7_75t_L g951 ( .A(n_170), .Y(n_951) );
INVxp67_ASAP7_75t_SL g1512 ( .A(n_172), .Y(n_1512) );
AOI221xp5_ASAP7_75t_L g1534 ( .A1(n_172), .A2(n_198), .B1(n_901), .B2(n_1535), .C(n_1536), .Y(n_1534) );
CKINVDCx5p33_ASAP7_75t_R g1577 ( .A(n_173), .Y(n_1577) );
INVx1_ASAP7_75t_L g918 ( .A(n_175), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_175), .A2(n_230), .B1(n_714), .B2(n_823), .Y(n_939) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_176), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_176), .B(n_288), .Y(n_1245) );
AND3x2_ASAP7_75t_L g1261 ( .A(n_176), .B(n_288), .C(n_1248), .Y(n_1261) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_178), .Y(n_352) );
INVx2_ASAP7_75t_L g301 ( .A(n_179), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_181), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g1578 ( .A(n_182), .Y(n_1578) );
INVx1_ASAP7_75t_L g967 ( .A(n_183), .Y(n_967) );
AOI21xp33_ASAP7_75t_L g994 ( .A1(n_183), .A2(n_451), .B(n_995), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_184), .A2(n_202), .B1(n_826), .B2(n_827), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_184), .A2(n_202), .B1(n_723), .B2(n_1173), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_186), .A2(n_209), .B1(n_1041), .B2(n_1043), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_186), .A2(n_209), .B1(n_1054), .B2(n_1056), .Y(n_1053) );
INVx1_ASAP7_75t_L g1606 ( .A(n_188), .Y(n_1606) );
CKINVDCx5p33_ASAP7_75t_R g922 ( .A(n_189), .Y(n_922) );
INVx1_ASAP7_75t_L g1248 ( .A(n_190), .Y(n_1248) );
INVx1_ASAP7_75t_L g1102 ( .A(n_191), .Y(n_1102) );
INVx1_ASAP7_75t_L g876 ( .A(n_192), .Y(n_876) );
CKINVDCx16_ASAP7_75t_R g605 ( .A(n_193), .Y(n_605) );
INVx1_ASAP7_75t_L g985 ( .A(n_194), .Y(n_985) );
INVx1_ASAP7_75t_L g879 ( .A(n_195), .Y(n_879) );
INVx1_ASAP7_75t_L g1583 ( .A(n_197), .Y(n_1583) );
OAI221xp5_ASAP7_75t_L g1593 ( .A1(n_197), .A2(n_540), .B1(n_775), .B2(n_1594), .C(n_1595), .Y(n_1593) );
INVxp67_ASAP7_75t_SL g1503 ( .A(n_198), .Y(n_1503) );
INVx1_ASAP7_75t_L g1584 ( .A(n_199), .Y(n_1584) );
OAI211xp5_ASAP7_75t_L g1598 ( .A1(n_199), .A2(n_542), .B(n_1599), .C(n_1604), .Y(n_1598) );
INVx1_ASAP7_75t_L g1209 ( .A(n_200), .Y(n_1209) );
AOI22xp33_ASAP7_75t_SL g936 ( .A1(n_201), .A2(n_253), .B1(n_517), .B2(n_714), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_201), .A2(n_253), .B1(n_846), .B2(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g1218 ( .A(n_203), .Y(n_1218) );
INVxp33_ASAP7_75t_L g1029 ( .A(n_204), .Y(n_1029) );
INVx1_ASAP7_75t_L g303 ( .A(n_205), .Y(n_303) );
INVx2_ASAP7_75t_L g323 ( .A(n_205), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_207), .A2(n_244), .B1(n_1130), .B2(n_1207), .Y(n_1206) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_207), .A2(n_244), .B1(n_1117), .B2(n_1118), .Y(n_1235) );
AOI22xp5_ASAP7_75t_L g1277 ( .A1(n_208), .A2(n_227), .B1(n_1264), .B2(n_1267), .Y(n_1277) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_210), .A2(n_542), .B1(n_1105), .B2(n_1108), .C(n_1114), .Y(n_1104) );
CKINVDCx5p33_ASAP7_75t_R g1196 ( .A(n_211), .Y(n_1196) );
INVx1_ASAP7_75t_L g1097 ( .A(n_212), .Y(n_1097) );
INVx1_ASAP7_75t_L g500 ( .A(n_213), .Y(n_500) );
AOI221xp5_ASAP7_75t_L g548 ( .A1(n_213), .A2(n_243), .B1(n_549), .B2(n_551), .C(n_554), .Y(n_548) );
INVx1_ASAP7_75t_L g1282 ( .A(n_214), .Y(n_1282) );
INVx1_ASAP7_75t_L g697 ( .A(n_215), .Y(n_697) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_216), .Y(n_317) );
INVx1_ASAP7_75t_L g1161 ( .A(n_217), .Y(n_1161) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_218), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g1551 ( .A(n_219), .Y(n_1551) );
CKINVDCx5p33_ASAP7_75t_R g1580 ( .A(n_220), .Y(n_1580) );
INVx1_ASAP7_75t_L g793 ( .A(n_221), .Y(n_793) );
INVx1_ASAP7_75t_L g816 ( .A(n_222), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_222), .A2(n_235), .B1(n_823), .B2(n_824), .Y(n_835) );
INVx1_ASAP7_75t_L g1205 ( .A(n_224), .Y(n_1205) );
OAI211xp5_ASAP7_75t_SL g1211 ( .A1(n_224), .A2(n_542), .B(n_1212), .C(n_1221), .Y(n_1211) );
INVx1_ASAP7_75t_L g786 ( .A(n_228), .Y(n_786) );
INVx1_ASAP7_75t_L g1509 ( .A(n_229), .Y(n_1509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_231), .Y(n_510) );
INVx1_ASAP7_75t_L g443 ( .A(n_233), .Y(n_443) );
INVx1_ASAP7_75t_L g809 ( .A(n_235), .Y(n_809) );
INVx1_ASAP7_75t_L g520 ( .A(n_236), .Y(n_520) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_236), .Y(n_577) );
OAI211xp5_ASAP7_75t_L g388 ( .A1(n_237), .A2(n_389), .B(n_394), .C(n_405), .Y(n_388) );
INVx1_ASAP7_75t_L g478 ( .A(n_237), .Y(n_478) );
INVx1_ASAP7_75t_L g617 ( .A(n_238), .Y(n_617) );
INVx1_ASAP7_75t_L g1158 ( .A(n_240), .Y(n_1158) );
INVx1_ASAP7_75t_L g701 ( .A(n_241), .Y(n_701) );
INVx1_ASAP7_75t_L g910 ( .A(n_242), .Y(n_910) );
AOI21xp33_ASAP7_75t_L g502 ( .A1(n_243), .A2(n_451), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g1249 ( .A(n_245), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_245), .B(n_1247), .Y(n_1269) );
INVx1_ASAP7_75t_L g1514 ( .A(n_246), .Y(n_1514) );
OAI211xp5_ASAP7_75t_L g1542 ( .A1(n_246), .A2(n_1543), .B(n_1545), .C(n_1552), .Y(n_1542) );
INVx1_ASAP7_75t_L g858 ( .A(n_247), .Y(n_858) );
INVx1_ASAP7_75t_L g1032 ( .A(n_248), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_248), .A2(n_269), .B1(n_627), .B2(n_855), .Y(n_1068) );
INVx1_ASAP7_75t_L g768 ( .A(n_249), .Y(n_768) );
INVx1_ASAP7_75t_L g1518 ( .A(n_250), .Y(n_1518) );
INVx1_ASAP7_75t_L g1028 ( .A(n_251), .Y(n_1028) );
INVx1_ASAP7_75t_L g1093 ( .A(n_252), .Y(n_1093) );
OAI211xp5_ASAP7_75t_L g333 ( .A1(n_254), .A2(n_334), .B(n_339), .C(n_346), .Y(n_333) );
INVx1_ASAP7_75t_L g439 ( .A(n_254), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g1569 ( .A1(n_256), .A2(n_1570), .B1(n_1571), .B2(n_1610), .Y(n_1569) );
CKINVDCx5p33_ASAP7_75t_R g1570 ( .A(n_256), .Y(n_1570) );
INVx1_ASAP7_75t_L g611 ( .A(n_257), .Y(n_611) );
INVx1_ASAP7_75t_L g807 ( .A(n_258), .Y(n_807) );
AO22x1_ASAP7_75t_L g1307 ( .A1(n_259), .A2(n_267), .B1(n_1262), .B2(n_1308), .Y(n_1307) );
CKINVDCx5p33_ASAP7_75t_R g1197 ( .A(n_260), .Y(n_1197) );
INVx1_ASAP7_75t_L g852 ( .A(n_261), .Y(n_852) );
INVx2_ASAP7_75t_L g300 ( .A(n_262), .Y(n_300) );
AO22x1_ASAP7_75t_L g1309 ( .A1(n_263), .A2(n_273), .B1(n_1264), .B2(n_1267), .Y(n_1309) );
NOR2xp33_ASAP7_75t_L g1162 ( .A(n_264), .B(n_1163), .Y(n_1162) );
CKINVDCx5p33_ASAP7_75t_R g970 ( .A(n_265), .Y(n_970) );
INVx1_ASAP7_75t_L g1152 ( .A(n_266), .Y(n_1152) );
CKINVDCx5p33_ASAP7_75t_R g1480 ( .A(n_268), .Y(n_1480) );
INVx1_ASAP7_75t_L g1033 ( .A(n_269), .Y(n_1033) );
INVx1_ASAP7_75t_L g687 ( .A(n_270), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_270), .A2(n_272), .B1(n_637), .B2(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g759 ( .A(n_271), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_271), .A2(n_278), .B1(n_582), .B2(n_587), .Y(n_783) );
INVx1_ASAP7_75t_L g684 ( .A(n_272), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_274), .Y(n_424) );
INVx1_ASAP7_75t_L g370 ( .A(n_276), .Y(n_370) );
BUFx3_ASAP7_75t_L g386 ( .A(n_276), .Y(n_386) );
BUFx3_ASAP7_75t_L g369 ( .A(n_277), .Y(n_369) );
INVx1_ASAP7_75t_L g379 ( .A(n_277), .Y(n_379) );
INVx1_ASAP7_75t_L g770 ( .A(n_278), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_280), .Y(n_398) );
XNOR2xp5_ASAP7_75t_L g1185 ( .A(n_281), .B(n_1186), .Y(n_1185) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_304), .B(n_1239), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_291), .Y(n_285) );
AND2x4_ASAP7_75t_L g1567 ( .A(n_286), .B(n_292), .Y(n_1567) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g1612 ( .A(n_287), .Y(n_1612) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_287), .B(n_289), .Y(n_1614) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_289), .B(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g313 ( .A(n_294), .B(n_314), .Y(n_313) );
OR2x6_ASAP7_75t_L g608 ( .A(n_294), .B(n_314), .Y(n_608) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g632 ( .A(n_295), .B(n_303), .Y(n_632) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g451 ( .A(n_296), .B(n_322), .Y(n_451) );
INVx8_ASAP7_75t_L g316 ( .A(n_297), .Y(n_316) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_298), .Y(n_453) );
OR2x6_ASAP7_75t_L g619 ( .A(n_298), .B(n_321), .Y(n_619) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_298), .B(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1597 ( .A(n_298), .Y(n_1597) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g326 ( .A(n_300), .Y(n_326) );
AND2x4_ASAP7_75t_L g331 ( .A(n_300), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g338 ( .A(n_300), .Y(n_338) );
INVx1_ASAP7_75t_L g345 ( .A(n_300), .Y(n_345) );
AND2x2_ASAP7_75t_L g350 ( .A(n_300), .B(n_301), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_301), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g332 ( .A(n_301), .Y(n_332) );
INVx1_ASAP7_75t_L g337 ( .A(n_301), .Y(n_337) );
INVx1_ASAP7_75t_L g354 ( .A(n_301), .Y(n_354) );
INVx1_ASAP7_75t_L g534 ( .A(n_301), .Y(n_534) );
AND2x4_ASAP7_75t_L g353 ( .A(n_302), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g855 ( .A(n_303), .B(n_357), .Y(n_855) );
OR2x2_ASAP7_75t_L g907 ( .A(n_303), .B(n_357), .Y(n_907) );
OAI22xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B1(n_954), .B2(n_955), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
XNOR2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_736), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
XNOR2x1_ASAP7_75t_L g309 ( .A(n_310), .B(n_603), .Y(n_309) );
XNOR2x1_ASAP7_75t_L g310 ( .A(n_311), .B(n_488), .Y(n_310) );
INVx1_ASAP7_75t_L g486 ( .A(n_312), .Y(n_486) );
OAI211xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_315), .B(n_360), .C(n_413), .Y(n_312) );
AOI31xp33_ASAP7_75t_L g850 ( .A1(n_313), .A2(n_851), .A3(n_856), .B(n_859), .Y(n_850) );
AOI31xp33_ASAP7_75t_L g1065 ( .A1(n_313), .A2(n_1066), .A3(n_1069), .B(n_1072), .Y(n_1065) );
AND2x4_ASAP7_75t_L g446 ( .A(n_314), .B(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g595 ( .A(n_314), .B(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g659 ( .A(n_314), .B(n_447), .Y(n_659) );
AOI211xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B(n_318), .C(n_333), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_316), .A2(n_616), .B1(n_617), .B2(n_618), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_316), .A2(n_618), .B1(n_686), .B2(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_316), .A2(n_806), .B1(n_860), .B2(n_861), .Y(n_859) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_316), .A2(n_861), .B1(n_877), .B2(n_912), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g1072 ( .A1(n_316), .A2(n_861), .B1(n_1028), .B2(n_1073), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g436 ( .A1(n_317), .A2(n_430), .B1(n_437), .B2(n_439), .Y(n_436) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .Y(n_319) );
AOI322xp5_ASAP7_75t_L g346 ( .A1(n_320), .A2(n_347), .A3(n_351), .B1(n_352), .B2(n_353), .C1(n_355), .C2(n_359), .Y(n_346) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g328 ( .A(n_321), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g612 ( .A(n_321), .B(n_532), .Y(n_612) );
AND2x4_ASAP7_75t_L g614 ( .A(n_321), .B(n_329), .Y(n_614) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g343 ( .A(n_323), .Y(n_343) );
INVx2_ASAP7_75t_L g459 ( .A(n_324), .Y(n_459) );
BUFx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g466 ( .A(n_325), .Y(n_466) );
INVx1_ASAP7_75t_L g494 ( .A(n_325), .Y(n_494) );
INVx1_ASAP7_75t_L g523 ( .A(n_326), .Y(n_523) );
AND2x4_ASAP7_75t_L g532 ( .A(n_326), .B(n_533), .Y(n_532) );
INVx5_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_328), .A2(n_612), .B1(n_857), .B2(n_858), .Y(n_856) );
AOI22xp33_ASAP7_75t_SL g908 ( .A1(n_328), .A2(n_612), .B1(n_909), .B2(n_910), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_328), .A2(n_612), .B1(n_933), .B2(n_934), .Y(n_932) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g462 ( .A(n_331), .Y(n_462) );
INVx3_ASAP7_75t_L g470 ( .A(n_331), .Y(n_470) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_331), .Y(n_829) );
AND2x4_ASAP7_75t_L g344 ( .A(n_332), .B(n_345), .Y(n_344) );
OAI221xp5_ASAP7_75t_L g1225 ( .A1(n_334), .A2(n_1103), .B1(n_1196), .B2(n_1197), .C(n_1226), .Y(n_1225) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g456 ( .A(n_336), .Y(n_456) );
INVx3_ASAP7_75t_L g501 ( .A(n_336), .Y(n_501) );
INVx2_ASAP7_75t_L g511 ( .A(n_336), .Y(n_511) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_337), .B(n_338), .Y(n_477) );
INVx1_ASAP7_75t_L g357 ( .A(n_338), .Y(n_357) );
NAND4xp25_ASAP7_75t_SL g609 ( .A(n_339), .B(n_610), .C(n_615), .D(n_620), .Y(n_609) );
NAND4xp25_ASAP7_75t_SL g695 ( .A(n_339), .B(n_696), .C(n_699), .D(n_706), .Y(n_695) );
CKINVDCx11_ASAP7_75t_R g339 ( .A(n_340), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g851 ( .A1(n_340), .A2(n_755), .B(n_852), .C(n_853), .Y(n_851) );
AOI211xp5_ASAP7_75t_L g904 ( .A1(n_340), .A2(n_824), .B(n_905), .C(n_906), .Y(n_904) );
NOR3xp33_ASAP7_75t_L g928 ( .A(n_340), .B(n_929), .C(n_931), .Y(n_928) );
AOI211xp5_ASAP7_75t_L g1066 ( .A1(n_340), .A2(n_755), .B(n_1067), .C(n_1068), .Y(n_1066) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVxp67_ASAP7_75t_L g358 ( .A(n_342), .Y(n_358) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g484 ( .A(n_343), .B(n_485), .Y(n_484) );
BUFx3_ASAP7_75t_L g544 ( .A(n_344), .Y(n_544) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_344), .Y(n_624) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_344), .Y(n_644) );
BUFx2_ASAP7_75t_L g705 ( .A(n_344), .Y(n_705) );
BUFx3_ASAP7_75t_L g1486 ( .A(n_344), .Y(n_1486) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g713 ( .A(n_348), .Y(n_713) );
INVx2_ASAP7_75t_SL g995 ( .A(n_348), .Y(n_995) );
INVx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_349), .Y(n_517) );
AND2x4_ASAP7_75t_L g541 ( .A(n_349), .B(n_531), .Y(n_541) );
BUFx2_ASAP7_75t_L g754 ( .A(n_349), .Y(n_754) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx3_ASAP7_75t_L g504 ( .A(n_350), .Y(n_504) );
AOI322xp5_ASAP7_75t_L g394 ( .A1(n_352), .A2(n_359), .A3(n_395), .B1(n_397), .B2(n_398), .C1(n_399), .C2(n_403), .Y(n_394) );
INVx2_ASAP7_75t_L g627 ( .A(n_353), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_353), .A2(n_355), .B1(n_700), .B2(n_701), .C1(n_702), .C2(n_703), .Y(n_699) );
INVx2_ASAP7_75t_L g854 ( .A(n_353), .Y(n_854) );
INVx2_ASAP7_75t_L g930 ( .A(n_353), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_354), .A2(n_520), .B1(n_521), .B2(n_522), .Y(n_519) );
INVx1_ASAP7_75t_L g763 ( .A(n_354), .Y(n_763) );
HB1xp67_ASAP7_75t_L g1006 ( .A(n_354), .Y(n_1006) );
AOI222xp33_ASAP7_75t_L g620 ( .A1(n_355), .A2(n_621), .B1(n_622), .B2(n_625), .C1(n_626), .C2(n_628), .Y(n_620) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI31xp33_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_371), .A3(n_388), .B(n_408), .Y(n_360) );
INVx4_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_363), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_363), .A2(n_682), .B1(n_683), .B2(n_684), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_363), .A2(n_381), .B1(n_806), .B2(n_807), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_363), .A2(n_673), .B1(n_879), .B2(n_880), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_363), .A2(n_381), .B1(n_1028), .B2(n_1029), .Y(n_1027) );
AND2x6_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
AND2x4_ASAP7_75t_L g670 ( .A(n_364), .B(n_671), .Y(n_670) );
AND2x4_ASAP7_75t_L g682 ( .A(n_364), .B(n_671), .Y(n_682) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g665 ( .A(n_365), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g375 ( .A(n_366), .Y(n_375) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_366), .Y(n_383) );
AND2x2_ASAP7_75t_L g417 ( .A(n_366), .B(n_410), .Y(n_417) );
INVx2_ASAP7_75t_L g448 ( .A(n_366), .Y(n_448) );
INVx1_ASAP7_75t_L g444 ( .A(n_367), .Y(n_444) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_367), .Y(n_649) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_367), .Y(n_658) );
INVx1_ASAP7_75t_L g1057 ( .A(n_367), .Y(n_1057) );
INVx2_ASAP7_75t_L g1131 ( .A(n_367), .Y(n_1131) );
BUFx6f_ASAP7_75t_L g1533 ( .A(n_367), .Y(n_1533) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g427 ( .A(n_368), .Y(n_427) );
INVx1_ASAP7_75t_L g557 ( .A(n_368), .Y(n_557) );
INVx1_ASAP7_75t_L g600 ( .A(n_368), .Y(n_600) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_368), .Y(n_724) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx2_ASAP7_75t_L g387 ( .A(n_369), .Y(n_387) );
AND2x2_ASAP7_75t_L g393 ( .A(n_369), .B(n_386), .Y(n_393) );
INVx1_ASAP7_75t_L g377 ( .A(n_370), .Y(n_377) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
INVx1_ASAP7_75t_L g397 ( .A(n_373), .Y(n_397) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g390 ( .A(n_374), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
AND2x6_ASAP7_75t_L g673 ( .A(n_374), .B(n_396), .Y(n_673) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x6_ASAP7_75t_L g403 ( .A(n_375), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g431 ( .A(n_376), .Y(n_431) );
INVx1_ASAP7_75t_L g1195 ( .A(n_376), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1561 ( .A(n_376), .B(n_591), .Y(n_1561) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x2_ASAP7_75t_L g435 ( .A(n_377), .B(n_378), .Y(n_435) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g396 ( .A(n_379), .B(n_386), .Y(n_396) );
INVx4_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_381), .A2(n_617), .B1(n_669), .B2(n_670), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_381), .A2(n_673), .B1(n_686), .B2(n_687), .C(n_688), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_381), .A2(n_682), .B1(n_876), .B2(n_877), .Y(n_875) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
AND2x2_ASAP7_75t_SL g399 ( .A(n_382), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g813 ( .A(n_382), .B(n_400), .Y(n_813) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx6_ASAP7_75t_L g553 ( .A(n_384), .Y(n_553) );
INVx2_ASAP7_75t_L g588 ( .A(n_384), .Y(n_588) );
AND2x2_ASAP7_75t_L g596 ( .A(n_384), .B(n_574), .Y(n_596) );
BUFx2_ASAP7_75t_L g654 ( .A(n_384), .Y(n_654) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g404 ( .A(n_385), .Y(n_404) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g402 ( .A(n_387), .Y(n_402) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI211xp5_ASAP7_75t_L g661 ( .A1(n_390), .A2(n_406), .B(n_662), .C(n_663), .Y(n_661) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_391), .Y(n_810) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_391), .Y(n_872) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_391), .Y(n_1060) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g406 ( .A(n_392), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g550 ( .A(n_392), .Y(n_550) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_392), .Y(n_692) );
INVx1_ASAP7_75t_L g798 ( .A(n_392), .Y(n_798) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_393), .Y(n_583) );
INVx2_ASAP7_75t_L g423 ( .A(n_395), .Y(n_423) );
INVx2_ASAP7_75t_SL g963 ( .A(n_395), .Y(n_963) );
INVx1_ASAP7_75t_L g978 ( .A(n_395), .Y(n_978) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_SL g442 ( .A(n_396), .Y(n_442) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_396), .Y(n_556) );
BUFx2_ASAP7_75t_L g648 ( .A(n_396), .Y(n_648) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_396), .Y(n_849) );
BUFx3_ASAP7_75t_L g1055 ( .A(n_396), .Y(n_1055) );
BUFx6f_ASAP7_75t_L g1174 ( .A(n_396), .Y(n_1174) );
HB1xp67_ASAP7_75t_L g1554 ( .A(n_396), .Y(n_1554) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_398), .A2(n_464), .B1(n_467), .B2(n_471), .Y(n_463) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g666 ( .A(n_401), .Y(n_666) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g571 ( .A(n_402), .Y(n_571) );
INVx3_ASAP7_75t_L g667 ( .A(n_403), .Y(n_667) );
AOI222xp33_ASAP7_75t_L g808 ( .A1(n_403), .A2(n_809), .B1(n_810), .B2(n_811), .C1(n_812), .C2(n_814), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_403), .A2(n_813), .B1(n_922), .B2(n_923), .Y(n_921) );
AOI222xp33_ASAP7_75t_L g1030 ( .A1(n_403), .A2(n_813), .B1(n_945), .B2(n_1031), .C1(n_1032), .C2(n_1033), .Y(n_1030) );
BUFx3_ASAP7_75t_L g580 ( .A(n_404), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_405), .B(n_917), .C(n_921), .Y(n_916) );
CKINVDCx8_ASAP7_75t_R g405 ( .A(n_406), .Y(n_405) );
INVx5_ASAP7_75t_L g804 ( .A(n_406), .Y(n_804) );
AOI211xp5_ASAP7_75t_L g870 ( .A1(n_406), .A2(n_871), .B(n_872), .C(n_873), .Y(n_870) );
OAI21xp33_ASAP7_75t_L g690 ( .A1(n_407), .A2(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_SL g676 ( .A(n_408), .Y(n_676) );
OAI31xp33_ASAP7_75t_L g915 ( .A1(n_408), .A2(n_916), .A3(n_924), .B(n_926), .Y(n_915) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
AND2x4_ASAP7_75t_L g694 ( .A(n_409), .B(n_411), .Y(n_694) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g447 ( .A(n_410), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g1010 ( .A(n_411), .Y(n_1010) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g418 ( .A(n_412), .Y(n_418) );
OR2x6_ASAP7_75t_L g450 ( .A(n_412), .B(n_451), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_449), .Y(n_413) );
OAI33xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_419), .A3(n_428), .B1(n_436), .B2(n_440), .B3(n_445), .Y(n_414) );
INVx1_ASAP7_75t_SL g646 ( .A(n_415), .Y(n_646) );
OAI33xp33_ASAP7_75t_L g961 ( .A1(n_415), .A2(n_962), .A3(n_966), .B1(n_971), .B2(n_977), .B3(n_982), .Y(n_961) );
OAI33xp33_ASAP7_75t_L g1574 ( .A1(n_415), .A2(n_982), .A3(n_1575), .B1(n_1579), .B2(n_1582), .B3(n_1585), .Y(n_1574) );
OR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
OR2x6_ASAP7_75t_L g559 ( .A(n_416), .B(n_418), .Y(n_559) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g728 ( .A(n_417), .Y(n_728) );
INVx2_ASAP7_75t_SL g1537 ( .A(n_417), .Y(n_1537) );
INVx2_ASAP7_75t_L g546 ( .A(n_418), .Y(n_546) );
AND2x4_ASAP7_75t_L g631 ( .A(n_418), .B(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g727 ( .A(n_418), .B(n_728), .Y(n_727) );
AND2x4_ASAP7_75t_L g821 ( .A(n_418), .B(n_632), .Y(n_821) );
BUFx2_ASAP7_75t_L g1154 ( .A(n_418), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_424), .B2(n_425), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_420), .A2(n_424), .B1(n_458), .B2(n_460), .Y(n_457) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_423), .A2(n_564), .B1(n_565), .B2(n_567), .Y(n_563) );
INVx2_ASAP7_75t_SL g1129 ( .A(n_423), .Y(n_1129) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g566 ( .A(n_427), .Y(n_566) );
OR2x2_ASAP7_75t_L g1562 ( .A(n_427), .B(n_591), .Y(n_1562) );
OAI22xp33_ASAP7_75t_SL g428 ( .A1(n_429), .A2(n_430), .B1(n_432), .B2(n_433), .Y(n_428) );
OAI22xp33_ASAP7_75t_L g452 ( .A1(n_429), .A2(n_432), .B1(n_453), .B2(n_454), .Y(n_452) );
OAI22xp33_ASAP7_75t_L g966 ( .A1(n_430), .A2(n_967), .B1(n_968), .B2(n_970), .Y(n_966) );
OAI22xp33_ASAP7_75t_L g1579 ( .A1(n_430), .A2(n_968), .B1(n_1580), .B2(n_1581), .Y(n_1579) );
OAI22xp33_ASAP7_75t_L g1582 ( .A1(n_430), .A2(n_1203), .B1(n_1583), .B2(n_1584), .Y(n_1582) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g972 ( .A(n_431), .Y(n_972) );
INVx1_ASAP7_75t_L g1016 ( .A(n_431), .Y(n_1016) );
HB1xp67_ASAP7_75t_L g1531 ( .A(n_431), .Y(n_1531) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g975 ( .A(n_434), .Y(n_975) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g438 ( .A(n_435), .Y(n_438) );
BUFx2_ASAP7_75t_L g969 ( .A(n_435), .Y(n_969) );
BUFx4f_ASAP7_75t_L g1204 ( .A(n_435), .Y(n_1204) );
BUFx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x6_ASAP7_75t_L g602 ( .A(n_438), .B(n_590), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g1192 ( .A1(n_438), .A2(n_1193), .B1(n_1196), .B2(n_1197), .C(n_1198), .Y(n_1192) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_440) );
INVx2_ASAP7_75t_L g594 ( .A(n_442), .Y(n_594) );
INVx1_ASAP7_75t_L g901 ( .A(n_442), .Y(n_901) );
INVx4_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g547 ( .A1(n_446), .A2(n_548), .B1(n_558), .B2(n_560), .C(n_568), .Y(n_547) );
AOI33xp33_ASAP7_75t_L g836 ( .A1(n_446), .A2(n_837), .A3(n_838), .B1(n_843), .B2(n_845), .B3(n_847), .Y(n_836) );
AOI33xp33_ASAP7_75t_L g940 ( .A1(n_446), .A2(n_837), .A3(n_941), .B1(n_944), .B2(n_946), .B3(n_949), .Y(n_940) );
AOI33xp33_ASAP7_75t_L g1052 ( .A1(n_446), .A2(n_837), .A3(n_1053), .B1(n_1058), .B2(n_1061), .B3(n_1064), .Y(n_1052) );
BUFx4f_ASAP7_75t_L g1132 ( .A(n_446), .Y(n_1132) );
BUFx4f_ASAP7_75t_L g1182 ( .A(n_446), .Y(n_1182) );
INVx2_ASAP7_75t_L g1559 ( .A(n_447), .Y(n_1559) );
AND2x4_ASAP7_75t_L g574 ( .A(n_448), .B(n_575), .Y(n_574) );
OAI33xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_452), .A3(n_457), .B1(n_463), .B2(n_472), .B3(n_479), .Y(n_449) );
OAI33xp33_ASAP7_75t_L g1501 ( .A1(n_450), .A2(n_1502), .A3(n_1508), .B1(n_1513), .B2(n_1517), .B3(n_1522), .Y(n_1501) );
OAI22xp33_ASAP7_75t_L g472 ( .A1(n_453), .A2(n_473), .B1(n_474), .B2(n_478), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g1100 ( .A1(n_453), .A2(n_476), .B1(n_1101), .B2(n_1102), .C(n_1103), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g1105 ( .A1(n_453), .A2(n_501), .B1(n_1090), .B2(n_1106), .C(n_1107), .Y(n_1105) );
BUFx2_ASAP7_75t_L g1226 ( .A(n_453), .Y(n_1226) );
OAI22xp33_ASAP7_75t_L g1508 ( .A1(n_453), .A2(n_1509), .B1(n_1510), .B2(n_1512), .Y(n_1508) );
OAI22xp33_ASAP7_75t_L g1517 ( .A1(n_453), .A2(n_1518), .B1(n_1519), .B2(n_1521), .Y(n_1517) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_456), .B(n_519), .Y(n_518) );
OR2x6_ASAP7_75t_L g775 ( .A(n_456), .B(n_525), .Y(n_775) );
OR2x2_ASAP7_75t_L g1234 ( .A(n_456), .B(n_525), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_458), .A2(n_964), .B1(n_965), .B2(n_990), .Y(n_989) );
OAI22xp5_ASAP7_75t_L g1502 ( .A1(n_458), .A2(n_1503), .B1(n_1504), .B2(n_1507), .Y(n_1502) );
OAI22xp5_ASAP7_75t_L g1513 ( .A1(n_458), .A2(n_1514), .B1(n_1515), .B2(n_1516), .Y(n_1513) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g894 ( .A(n_460), .Y(n_894) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g536 ( .A(n_461), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g773 ( .A(n_462), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_464), .A2(n_1097), .B1(n_1098), .B2(n_1099), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1594 ( .A1(n_464), .A2(n_828), .B1(n_1577), .B2(n_1578), .Y(n_1594) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g1215 ( .A(n_466), .Y(n_1215) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g718 ( .A(n_469), .Y(n_718) );
INVx2_ASAP7_75t_L g1044 ( .A(n_469), .Y(n_1044) );
INVx3_ASAP7_75t_L g1112 ( .A(n_469), .Y(n_1112) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g497 ( .A(n_470), .Y(n_497) );
INVx3_ASAP7_75t_L g991 ( .A(n_470), .Y(n_991) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g993 ( .A(n_476), .Y(n_993) );
BUFx3_ASAP7_75t_L g1511 ( .A(n_476), .Y(n_1511) );
OAI221xp5_ASAP7_75t_L g1595 ( .A1(n_476), .A2(n_1103), .B1(n_1580), .B2(n_1581), .C(n_1596), .Y(n_1595) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI33xp33_ASAP7_75t_L g630 ( .A1(n_480), .A2(n_631), .A3(n_633), .B1(n_636), .B2(n_640), .B3(n_642), .Y(n_630) );
AOI33xp33_ASAP7_75t_L g819 ( .A1(n_480), .A2(n_820), .A3(n_822), .B1(n_825), .B2(n_830), .B3(n_835), .Y(n_819) );
AOI33xp33_ASAP7_75t_L g935 ( .A1(n_480), .A2(n_631), .A3(n_936), .B1(n_937), .B2(n_938), .B3(n_939), .Y(n_935) );
INVx6_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx5_ASAP7_75t_L g720 ( .A(n_481), .Y(n_720) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g573 ( .A(n_482), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g590 ( .A(n_483), .B(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g1483 ( .A(n_483), .B(n_531), .Y(n_1483) );
BUFx2_ASAP7_75t_L g514 ( .A(n_484), .Y(n_514) );
INVx2_ASAP7_75t_L g758 ( .A(n_484), .Y(n_758) );
NAND4xp25_ASAP7_75t_L g489 ( .A(n_490), .B(n_547), .C(n_585), .D(n_597), .Y(n_489) );
OAI31xp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_528), .A3(n_539), .B(n_545), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_499), .B1(n_505), .B2(n_509), .C(n_515), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_495), .B1(n_496), .B2(n_498), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_493), .A2(n_506), .B1(n_507), .B2(n_508), .Y(n_505) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g998 ( .A(n_494), .Y(n_998) );
INVx1_ASAP7_75t_L g1110 ( .A(n_494), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_495), .A2(n_498), .B1(n_555), .B2(n_557), .Y(n_554) );
INVx2_ASAP7_75t_L g641 ( .A(n_496), .Y(n_641) );
INVx2_ASAP7_75t_SL g711 ( .A(n_496), .Y(n_711) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g507 ( .A(n_497), .Y(n_507) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_497), .Y(n_752) );
INVx1_ASAP7_75t_L g1506 ( .A(n_497), .Y(n_1506) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g1520 ( .A(n_501), .Y(n_1520) );
BUFx2_ASAP7_75t_L g634 ( .A(n_503), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_503), .B(n_747), .Y(n_746) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g513 ( .A(n_504), .Y(n_513) );
INVx2_ASAP7_75t_SL g1047 ( .A(n_504), .Y(n_1047) );
AOI222xp33_ASAP7_75t_L g585 ( .A1(n_506), .A2(n_516), .B1(n_586), .B2(n_592), .C1(n_593), .C2(n_595), .Y(n_585) );
INVx1_ASAP7_75t_L g639 ( .A(n_507), .Y(n_639) );
INVx2_ASAP7_75t_L g889 ( .A(n_507), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_508), .A2(n_510), .B1(n_598), .B2(n_601), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_512), .Y(n_509) );
BUFx3_ASAP7_75t_L g823 ( .A(n_513), .Y(n_823) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_518), .C(n_524), .Y(n_515) );
NAND2x1p5_ASAP7_75t_L g1498 ( .A(n_522), .B(n_1496), .Y(n_1498) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OR2x6_ASAP7_75t_L g765 ( .A(n_523), .B(n_525), .Y(n_765) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g747 ( .A(n_525), .Y(n_747) );
INVx1_ASAP7_75t_L g764 ( .A(n_525), .Y(n_764) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_530), .A2(n_536), .B1(n_767), .B2(n_768), .Y(n_766) );
INVx3_ASAP7_75t_L g1117 ( .A(n_530), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_530), .A2(n_536), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx2_ASAP7_75t_L g538 ( .A(n_531), .Y(n_538) );
INVx1_ASAP7_75t_L g638 ( .A(n_532), .Y(n_638) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_532), .Y(n_751) );
BUFx2_ASAP7_75t_L g826 ( .A(n_532), .Y(n_826) );
BUFx6f_ASAP7_75t_L g833 ( .A(n_532), .Y(n_833) );
BUFx2_ASAP7_75t_L g893 ( .A(n_532), .Y(n_893) );
BUFx6f_ASAP7_75t_L g1042 ( .A(n_532), .Y(n_1042) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx3_ASAP7_75t_L g1118 ( .A(n_536), .Y(n_1118) );
AND2x4_ASAP7_75t_L g543 ( .A(n_537), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
CKINVDCx6p67_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g769 ( .A1(n_541), .A2(n_770), .B1(n_771), .B2(n_772), .C(n_774), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g1148 ( .A1(n_541), .A2(n_774), .B1(n_1149), .B2(n_1151), .C(n_1152), .Y(n_1148) );
INVx8_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI221xp5_ASAP7_75t_SL g749 ( .A1(n_543), .A2(n_750), .B1(n_753), .B2(n_759), .C(n_760), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g1138 ( .A1(n_543), .A2(n_1139), .B1(n_1140), .B2(n_1143), .C(n_1144), .Y(n_1138) );
INVx1_ASAP7_75t_L g756 ( .A(n_544), .Y(n_756) );
INVx1_ASAP7_75t_L g776 ( .A(n_545), .Y(n_776) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp67_ASAP7_75t_L g745 ( .A(n_546), .B(n_746), .Y(n_745) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g782 ( .A(n_550), .Y(n_782) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_553), .Y(n_562) );
INVx2_ASAP7_75t_L g652 ( .A(n_553), .Y(n_652) );
INVx2_ASAP7_75t_L g671 ( .A(n_553), .Y(n_671) );
INVx1_ASAP7_75t_L g731 ( .A(n_553), .Y(n_731) );
INVx2_ASAP7_75t_L g840 ( .A(n_553), .Y(n_840) );
INVx1_ASAP7_75t_L g1178 ( .A(n_553), .Y(n_1178) );
INVx1_ASAP7_75t_L g942 ( .A(n_555), .Y(n_942) );
INVx1_ASAP7_75t_L g1124 ( .A(n_555), .Y(n_1124) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
BUFx3_ASAP7_75t_L g844 ( .A(n_556), .Y(n_844) );
AND2x4_ASAP7_75t_L g1544 ( .A(n_556), .B(n_1528), .Y(n_1544) );
INVx1_ASAP7_75t_L g943 ( .A(n_557), .Y(n_943) );
INVx1_ASAP7_75t_L g950 ( .A(n_557), .Y(n_950) );
OAI22xp33_ASAP7_75t_L g962 ( .A1(n_557), .A2(n_963), .B1(n_964), .B2(n_965), .Y(n_962) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_559), .Y(n_837) );
CKINVDCx5p33_ASAP7_75t_R g1120 ( .A(n_559), .Y(n_1120) );
OAI22xp5_ASAP7_75t_SL g1191 ( .A1(n_559), .A2(n_1192), .B1(n_1199), .B2(n_1200), .Y(n_1191) );
INVx4_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g899 ( .A(n_562), .Y(n_899) );
INVx1_ASAP7_75t_L g886 ( .A(n_565), .Y(n_886) );
INVx1_ASAP7_75t_L g902 ( .A(n_565), .Y(n_902) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g794 ( .A(n_569), .Y(n_794) );
INVx1_ASAP7_75t_L g1085 ( .A(n_569), .Y(n_1085) );
INVx2_ASAP7_75t_L g1168 ( .A(n_569), .Y(n_1168) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g1547 ( .A(n_571), .Y(n_1547) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
OR2x6_ASAP7_75t_L g578 ( .A(n_573), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g584 ( .A(n_573), .Y(n_584) );
INVx1_ASAP7_75t_L g1541 ( .A(n_574), .Y(n_1541) );
AND2x4_ASAP7_75t_L g1546 ( .A(n_574), .B(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g792 ( .A(n_578), .Y(n_792) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_579), .B(n_1541), .Y(n_1550) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g1166 ( .A(n_581), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
INVx1_ASAP7_75t_L g1063 ( .A(n_582), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g1180 ( .A(n_582), .Y(n_1180) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g656 ( .A(n_583), .Y(n_656) );
INVx2_ASAP7_75t_SL g920 ( .A(n_583), .Y(n_920) );
BUFx3_ASAP7_75t_L g945 ( .A(n_583), .Y(n_945) );
BUFx4f_ASAP7_75t_L g1122 ( .A(n_583), .Y(n_1122) );
AND2x4_ASAP7_75t_L g1527 ( .A(n_583), .B(n_1528), .Y(n_1527) );
AND2x2_ASAP7_75t_L g796 ( .A(n_584), .B(n_797), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_586), .A2(n_593), .B1(n_789), .B2(n_790), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g1088 ( .A1(n_586), .A2(n_593), .B1(n_1089), .B2(n_1090), .C(n_1091), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_586), .A2(n_593), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_587), .Y(n_1059) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g846 ( .A(n_588), .Y(n_846) );
AND2x2_ASAP7_75t_L g593 ( .A(n_589), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x6_ASAP7_75t_L g599 ( .A(n_590), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_590), .B(n_600), .Y(n_1013) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_590), .B(n_1016), .Y(n_1015) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_590), .B(n_1018), .Y(n_1017) );
INVx2_ASAP7_75t_L g1528 ( .A(n_591), .Y(n_1528) );
OR2x6_ASAP7_75t_L g744 ( .A(n_595), .B(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g1476 ( .A(n_595), .Y(n_1476) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_598), .A2(n_601), .B1(n_786), .B2(n_787), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_598), .A2(n_601), .B1(n_1160), .B2(n_1161), .Y(n_1159) );
CKINVDCx6p67_ASAP7_75t_R g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g780 ( .A(n_600), .Y(n_780) );
CKINVDCx6p67_ASAP7_75t_R g601 ( .A(n_602), .Y(n_601) );
OA22x2_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_677), .B1(n_678), .B2(n_735), .Y(n_603) );
INVx1_ASAP7_75t_L g735 ( .A(n_604), .Y(n_735) );
XNOR2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
AOI211xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_609), .B(n_629), .C(n_660), .Y(n_606) );
AOI221x1_ASAP7_75t_L g679 ( .A1(n_607), .A2(n_680), .B1(n_693), .B2(n_695), .C(n_708), .Y(n_679) );
CKINVDCx16_ASAP7_75t_R g607 ( .A(n_608), .Y(n_607) );
AOI31xp33_ASAP7_75t_L g903 ( .A1(n_608), .A2(n_904), .A3(n_908), .B(n_911), .Y(n_903) );
AO21x1_ASAP7_75t_SL g927 ( .A1(n_608), .A2(n_928), .B(n_932), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_612), .A2(n_614), .B1(n_697), .B2(n_698), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g1069 ( .A1(n_612), .A2(n_614), .B1(n_1070), .B2(n_1071), .Y(n_1069) );
INVx4_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx5_ASAP7_75t_L g861 ( .A(n_619), .Y(n_861) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g824 ( .A(n_623), .Y(n_824) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_624), .Y(n_635) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_630), .B(n_645), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_631), .B(n_710), .C(n_712), .Y(n_709) );
BUFx2_ASAP7_75t_SL g1103 ( .A(n_632), .Y(n_1103) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_SL g715 ( .A(n_644), .Y(n_715) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_644), .Y(n_896) );
AOI33xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .A3(n_650), .B1(n_653), .B2(n_657), .B3(n_659), .Y(n_645) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g1557 ( .A(n_652), .Y(n_1557) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g1535 ( .A(n_656), .Y(n_1535) );
NAND3xp33_ASAP7_75t_L g729 ( .A(n_659), .B(n_730), .C(n_732), .Y(n_729) );
AOI33xp33_ASAP7_75t_L g778 ( .A1(n_659), .A2(n_726), .A3(n_779), .B1(n_781), .B2(n_783), .B3(n_784), .Y(n_778) );
NAND3xp33_ASAP7_75t_L g897 ( .A(n_659), .B(n_898), .C(n_900), .Y(n_897) );
INVx1_ASAP7_75t_L g982 ( .A(n_659), .Y(n_982) );
AOI31xp33_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_668), .A3(n_672), .B(n_676), .Y(n_660) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g689 ( .A(n_665), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_670), .A2(n_673), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_673), .A2(n_682), .B1(n_816), .B2(n_817), .Y(n_815) );
CKINVDCx6p67_ASAP7_75t_R g925 ( .A(n_673), .Y(n_925) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g734 ( .A(n_679), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_685), .Y(n_680) );
INVx1_ASAP7_75t_L g842 ( .A(n_692), .Y(n_842) );
BUFx6f_ASAP7_75t_L g948 ( .A(n_692), .Y(n_948) );
AND2x4_ASAP7_75t_L g1539 ( .A(n_692), .B(n_1540), .Y(n_1539) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI211x1_ASAP7_75t_SL g802 ( .A1(n_694), .A2(n_803), .B(n_818), .C(n_850), .Y(n_802) );
AO211x2_ASAP7_75t_L g868 ( .A1(n_694), .A2(n_869), .B(n_881), .C(n_903), .Y(n_868) );
INVx1_ASAP7_75t_L g1035 ( .A(n_694), .Y(n_1035) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND4xp25_ASAP7_75t_L g708 ( .A(n_709), .B(n_716), .C(n_721), .D(n_729), .Y(n_708) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .C(n_720), .Y(n_716) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_720), .B(n_888), .C(n_890), .Y(n_887) );
AOI33xp33_ASAP7_75t_L g1037 ( .A1(n_720), .A2(n_1038), .A3(n_1040), .B1(n_1045), .B2(n_1048), .B3(n_1051), .Y(n_1037) );
CKINVDCx8_ASAP7_75t_R g1522 ( .A(n_720), .Y(n_1522) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .C(n_726), .Y(n_721) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g980 ( .A(n_724), .Y(n_980) );
INVx1_ASAP7_75t_L g1126 ( .A(n_724), .Y(n_1126) );
NAND3xp33_ASAP7_75t_L g882 ( .A(n_726), .B(n_883), .C(n_884), .Y(n_882) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B1(n_865), .B2(n_953), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AOI21x1_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_800), .B(n_864), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g864 ( .A(n_740), .B(n_801), .Y(n_864) );
XOR2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_799), .Y(n_740) );
NOR3xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_748), .C(n_777), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_744), .B(n_985), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_744), .B(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1163 ( .A(n_744), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_744), .B(n_1209), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1589 ( .A(n_744), .B(n_1590), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_747), .B(n_1006), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_747), .B(n_1006), .Y(n_1115) );
AOI31xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_766), .A3(n_769), .B(n_776), .Y(n_748) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g1107 ( .A(n_757), .Y(n_1107) );
INVx2_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g1220 ( .A(n_758), .Y(n_1220) );
NAND2x1p5_ASAP7_75t_L g761 ( .A(n_762), .B(n_764), .Y(n_761) );
NAND2x1_ASAP7_75t_SL g1495 ( .A(n_762), .B(n_1496), .Y(n_1495) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
CKINVDCx11_ASAP7_75t_R g1008 ( .A(n_765), .Y(n_1008) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
OAI31xp33_ASAP7_75t_L g1523 ( .A1(n_776), .A2(n_1524), .A3(n_1542), .B(n_1560), .Y(n_1523) );
NAND4xp25_ASAP7_75t_L g777 ( .A(n_778), .B(n_785), .C(n_788), .D(n_791), .Y(n_777) );
AOI221xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_794), .B2(n_795), .C(n_796), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g1084 ( .A1(n_792), .A2(n_796), .B1(n_1085), .B2(n_1086), .C(n_1087), .Y(n_1084) );
AOI22xp5_ASAP7_75t_L g1167 ( .A1(n_792), .A2(n_1168), .B1(n_1169), .B2(n_1170), .Y(n_1167) );
NOR3xp33_ASAP7_75t_L g960 ( .A(n_796), .B(n_961), .C(n_983), .Y(n_960) );
BUFx2_ASAP7_75t_L g1188 ( .A(n_796), .Y(n_1188) );
NOR3xp33_ASAP7_75t_L g1573 ( .A(n_796), .B(n_1574), .C(n_1588), .Y(n_1573) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g863 ( .A(n_802), .Y(n_863) );
NAND4xp25_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .C(n_808), .D(n_815), .Y(n_803) );
NAND4xp25_ASAP7_75t_L g1023 ( .A(n_804), .B(n_1024), .C(n_1027), .D(n_1030), .Y(n_1023) );
BUFx4f_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g874 ( .A(n_813), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_836), .Y(n_818) );
BUFx3_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NAND3xp33_ASAP7_75t_L g891 ( .A(n_821), .B(n_892), .C(n_895), .Y(n_891) );
INVx2_ASAP7_75t_L g1039 ( .A(n_821), .Y(n_1039) );
INVx2_ASAP7_75t_SL g827 ( .A(n_828), .Y(n_827) );
INVx4_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
BUFx3_ASAP7_75t_L g834 ( .A(n_829), .Y(n_834) );
INVx2_ASAP7_75t_SL g1000 ( .A(n_829), .Y(n_1000) );
INVx2_ASAP7_75t_SL g1050 ( .A(n_829), .Y(n_1050) );
INVx2_ASAP7_75t_SL g1098 ( .A(n_829), .Y(n_1098) );
INVx2_ASAP7_75t_SL g1601 ( .A(n_829), .Y(n_1601) );
INVx3_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_SL g832 ( .A(n_833), .Y(n_832) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_833), .B(n_1483), .Y(n_1491) );
AOI33xp33_ASAP7_75t_L g1171 ( .A1(n_837), .A2(n_1172), .A3(n_1175), .B1(n_1179), .B2(n_1181), .B3(n_1182), .Y(n_1171) );
BUFx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_840), .Y(n_947) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
BUFx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
BUFx4f_ASAP7_75t_L g885 ( .A(n_849), .Y(n_885) );
INVx1_ASAP7_75t_L g1018 ( .A(n_849), .Y(n_1018) );
INVx1_ASAP7_75t_L g953 ( .A(n_865), .Y(n_953) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
XNOR2x1_ASAP7_75t_L g866 ( .A(n_867), .B(n_913), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g869 ( .A(n_870), .B(n_875), .C(n_878), .Y(n_869) );
NAND4xp25_ASAP7_75t_L g881 ( .A(n_882), .B(n_887), .C(n_891), .D(n_897), .Y(n_881) );
INVx1_ASAP7_75t_L g1217 ( .A(n_894), .Y(n_1217) );
AND4x1_ASAP7_75t_L g914 ( .A(n_915), .B(n_927), .C(n_935), .D(n_940), .Y(n_914) );
NAND4xp25_ASAP7_75t_L g952 ( .A(n_915), .B(n_927), .C(n_935), .D(n_940), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
XNOR2xp5_ASAP7_75t_L g955 ( .A(n_956), .B(n_1076), .Y(n_955) );
AOI22xp33_ASAP7_75t_SL g956 ( .A1(n_957), .A2(n_1019), .B1(n_1020), .B2(n_1075), .Y(n_956) );
INVx1_ASAP7_75t_L g1075 ( .A(n_957), .Y(n_1075) );
HB1xp67_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
AND4x1_ASAP7_75t_L g959 ( .A(n_960), .B(n_984), .C(n_986), .D(n_1011), .Y(n_959) );
INVx2_ASAP7_75t_SL g968 ( .A(n_969), .Y(n_968) );
OAI21xp33_ASAP7_75t_SL g992 ( .A1(n_970), .A2(n_993), .B(n_994), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_973), .B1(n_974), .B2(n_976), .Y(n_971) );
OAI221xp5_ASAP7_75t_L g1200 ( .A1(n_972), .A2(n_1201), .B1(n_1202), .B2(n_1205), .C(n_1206), .Y(n_1200) );
INVx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_978), .A2(n_979), .B1(n_980), .B2(n_981), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g1585 ( .A1(n_978), .A2(n_1532), .B1(n_1586), .B2(n_1587), .Y(n_1585) );
OAI22xp33_ASAP7_75t_L g1575 ( .A1(n_980), .A2(n_1576), .B1(n_1577), .B2(n_1578), .Y(n_1575) );
OAI31xp33_ASAP7_75t_L g986 ( .A1(n_987), .A2(n_988), .A3(n_996), .B(n_1009), .Y(n_986) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
BUFx3_ASAP7_75t_L g1232 ( .A(n_991), .Y(n_1232) );
AND2x4_ASAP7_75t_L g1482 ( .A(n_991), .B(n_1483), .Y(n_1482) );
OAI221xp5_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_999), .B1(n_1000), .B2(n_1001), .C(n_1002), .Y(n_997) );
INVx1_ASAP7_75t_L g1229 ( .A(n_998), .Y(n_1229) );
OAI221xp5_ASAP7_75t_L g1599 ( .A1(n_998), .A2(n_1600), .B1(n_1601), .B2(n_1602), .C(n_1603), .Y(n_1599) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1005), .B1(n_1007), .B2(n_1008), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_1005), .A2(n_1008), .B1(n_1222), .B2(n_1223), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1604 ( .A1(n_1005), .A2(n_1008), .B1(n_1605), .B2(n_1606), .Y(n_1604) );
AOI22xp5_ASAP7_75t_L g1114 ( .A1(n_1008), .A2(n_1086), .B1(n_1087), .B2(n_1115), .Y(n_1114) );
OAI31xp33_ASAP7_75t_L g1094 ( .A1(n_1009), .A2(n_1095), .A3(n_1104), .B(n_1116), .Y(n_1094) );
OAI31xp33_ASAP7_75t_L g1591 ( .A1(n_1009), .A2(n_1592), .A3(n_1593), .B(n_1598), .Y(n_1591) );
BUFx8_ASAP7_75t_SL g1009 ( .A(n_1010), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1014), .Y(n_1011) );
INVx2_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1022), .Y(n_1074) );
AOI211x1_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1034), .B(n_1036), .C(n_1065), .Y(n_1022) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1052), .Y(n_1036) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
BUFx3_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
BUFx3_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1047), .Y(n_1142) );
BUFx2_ASAP7_75t_L g1150 ( .A(n_1047), .Y(n_1150) );
AND2x4_ASAP7_75t_L g1489 ( .A(n_1047), .B(n_1483), .Y(n_1489) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx2_ASAP7_75t_SL g1576 ( .A(n_1055), .Y(n_1576) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
AOI22xp5_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1078), .B1(n_1183), .B2(n_1184), .Y(n_1076) );
INVxp67_ASAP7_75t_SL g1077 ( .A(n_1078), .Y(n_1077) );
INVxp67_ASAP7_75t_SL g1078 ( .A(n_1079), .Y(n_1078) );
AOI22xp5_ASAP7_75t_L g1079 ( .A1(n_1080), .A2(n_1081), .B1(n_1133), .B2(n_1134), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
NAND4xp75_ASAP7_75t_SL g1082 ( .A(n_1083), .B(n_1092), .C(n_1094), .D(n_1119), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1088), .Y(n_1083) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1085), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_1089), .A2(n_1109), .B1(n_1111), .B2(n_1113), .Y(n_1108) );
BUFx2_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1112), .Y(n_1515) );
AOI33xp33_ASAP7_75t_L g1119 ( .A1(n_1120), .A2(n_1121), .A3(n_1123), .B1(n_1127), .B2(n_1128), .B3(n_1132), .Y(n_1119) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
CKINVDCx5p33_ASAP7_75t_R g1199 ( .A(n_1132), .Y(n_1199) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
XNOR2xp5_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
NOR4xp75_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1155), .C(n_1162), .D(n_1164), .Y(n_1136) );
AOI31xp33_ASAP7_75t_SL g1137 ( .A1(n_1138), .A2(n_1145), .A3(n_1148), .B(n_1153), .Y(n_1137) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
CKINVDCx8_ASAP7_75t_R g1153 ( .A(n_1154), .Y(n_1153) );
OAI31xp33_ASAP7_75t_L g1210 ( .A1(n_1154), .A2(n_1211), .A3(n_1224), .B(n_1235), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1159), .Y(n_1155) );
NAND3xp33_ASAP7_75t_SL g1164 ( .A(n_1165), .B(n_1167), .C(n_1171), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
BUFx2_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
BUFx3_ASAP7_75t_L g1207 ( .A(n_1174), .Y(n_1207) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
HB1xp67_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
AND4x1_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1208), .C(n_1210), .D(n_1236), .Y(n_1186) );
NOR3xp33_ASAP7_75t_SL g1187 ( .A(n_1188), .B(n_1189), .C(n_1191), .Y(n_1187) );
BUFx2_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
BUFx2_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
OAI221xp5_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1216), .B1(n_1217), .B2(n_1218), .C(n_1219), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_1228), .A2(n_1230), .B1(n_1231), .B2(n_1233), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
CKINVDCx5p33_ASAP7_75t_R g1231 ( .A(n_1232), .Y(n_1231) );
NOR2xp33_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1238), .Y(n_1236) );
OAI21xp5_ASAP7_75t_SL g1239 ( .A1(n_1240), .A2(n_1250), .B(n_1465), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
OAI22xp33_ASAP7_75t_L g1326 ( .A1(n_1242), .A2(n_1327), .B1(n_1328), .B2(n_1329), .Y(n_1326) );
BUFx3_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
OAI22xp33_ASAP7_75t_L g1281 ( .A1(n_1243), .A2(n_1282), .B1(n_1283), .B2(n_1284), .Y(n_1281) );
OAI22xp5_ASAP7_75t_L g1287 ( .A1(n_1243), .A2(n_1284), .B1(n_1288), .B2(n_1289), .Y(n_1287) );
OAI22xp33_ASAP7_75t_L g1334 ( .A1(n_1243), .A2(n_1335), .B1(n_1336), .B2(n_1337), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1246), .Y(n_1244) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1245), .Y(n_1266) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1245), .B(n_1269), .Y(n_1284) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1246), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1249), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1249), .Y(n_1260) );
NOR4xp25_ASAP7_75t_L g1250 ( .A(n_1251), .B(n_1392), .C(n_1427), .D(n_1456), .Y(n_1250) );
NAND3xp33_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1338), .C(n_1364), .Y(n_1251) );
OAI21xp5_ASAP7_75t_L g1252 ( .A1(n_1253), .A2(n_1299), .B(n_1320), .Y(n_1252) );
AOI22xp5_ASAP7_75t_L g1253 ( .A1(n_1254), .A2(n_1290), .B1(n_1294), .B2(n_1298), .Y(n_1253) );
NOR2xp33_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1270), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1255), .B(n_1312), .Y(n_1319) );
NOR2xp33_ASAP7_75t_L g1360 ( .A(n_1255), .B(n_1361), .Y(n_1360) );
INVx3_ASAP7_75t_L g1375 ( .A(n_1255), .Y(n_1375) );
NOR2xp33_ASAP7_75t_L g1394 ( .A(n_1255), .B(n_1300), .Y(n_1394) );
AOI21xp5_ASAP7_75t_L g1411 ( .A1(n_1255), .A2(n_1412), .B(n_1413), .Y(n_1411) );
AOI211xp5_ASAP7_75t_L g1428 ( .A1(n_1255), .A2(n_1404), .B(n_1429), .C(n_1434), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1255), .B(n_1356), .Y(n_1460) );
CKINVDCx5p33_ASAP7_75t_R g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1256), .Y(n_1298) );
INVx1_ASAP7_75t_SL g1305 ( .A(n_1256), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1256), .B(n_1312), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1256), .B(n_1306), .Y(n_1342) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1256), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1358 ( .A(n_1256), .B(n_1272), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1366 ( .A(n_1256), .B(n_1367), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1256), .B(n_1343), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1256), .B(n_1272), .Y(n_1418) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1256), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1263), .Y(n_1256) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1258), .Y(n_1323) );
AND2x4_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1261), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1259), .B(n_1261), .Y(n_1308) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
AND2x4_ASAP7_75t_L g1262 ( .A(n_1260), .B(n_1261), .Y(n_1262) );
INVx2_ASAP7_75t_L g1325 ( .A(n_1262), .Y(n_1325) );
AND2x4_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1266), .Y(n_1264) );
OAI21xp33_ASAP7_75t_SL g1613 ( .A1(n_1265), .A2(n_1612), .B(n_1614), .Y(n_1613) );
AND2x4_ASAP7_75t_L g1267 ( .A(n_1266), .B(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1279), .Y(n_1270) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1271), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1271), .B(n_1292), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1271), .B(n_1302), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1275), .Y(n_1271) );
INVx3_ASAP7_75t_L g1297 ( .A(n_1272), .Y(n_1297) );
INVx4_ASAP7_75t_L g1343 ( .A(n_1272), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1272), .B(n_1292), .Y(n_1401) );
AND2x4_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1274), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1275), .B(n_1354), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_1275), .B(n_1285), .Y(n_1384) );
OR2x2_ASAP7_75t_L g1405 ( .A(n_1275), .B(n_1406), .Y(n_1405) );
NOR2xp33_ASAP7_75t_L g1414 ( .A(n_1275), .B(n_1285), .Y(n_1414) );
OR2x2_ASAP7_75t_L g1463 ( .A(n_1275), .B(n_1374), .Y(n_1463) );
BUFx3_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1276), .B(n_1292), .Y(n_1291) );
INVx2_ASAP7_75t_L g1295 ( .A(n_1276), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1276), .B(n_1302), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1276), .B(n_1346), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1276), .B(n_1374), .Y(n_1412) );
OR2x2_ASAP7_75t_L g1421 ( .A(n_1276), .B(n_1410), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1278), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1279), .B(n_1297), .Y(n_1296) );
AOI21xp5_ASAP7_75t_L g1380 ( .A1(n_1279), .A2(n_1342), .B(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1279), .Y(n_1406) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1279), .B(n_1368), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1285), .Y(n_1279) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1280), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1280), .B(n_1286), .Y(n_1302) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1280), .Y(n_1374) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1284), .Y(n_1330) );
HB1xp67_ASAP7_75t_L g1337 ( .A(n_1284), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1285), .B(n_1295), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1285), .B(n_1293), .Y(n_1346) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1285), .Y(n_1354) );
INVx2_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1286), .B(n_1293), .Y(n_1292) );
AOI21xp33_ASAP7_75t_SL g1423 ( .A1(n_1290), .A2(n_1424), .B(n_1425), .Y(n_1423) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1292), .B(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1292), .Y(n_1410) );
OR2x2_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1296), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1295), .B(n_1346), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1295), .B(n_1343), .Y(n_1368) );
NOR2x1_ASAP7_75t_L g1388 ( .A(n_1295), .B(n_1374), .Y(n_1388) );
NAND4xp25_ASAP7_75t_L g1389 ( .A(n_1295), .B(n_1318), .C(n_1348), .D(n_1390), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1295), .B(n_1400), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1295), .B(n_1302), .Y(n_1455) );
INVx2_ASAP7_75t_L g1318 ( .A(n_1297), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1297), .B(n_1345), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1297), .B(n_1301), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1297), .B(n_1414), .Y(n_1440) );
OR2x2_ASAP7_75t_L g1457 ( .A(n_1297), .B(n_1363), .Y(n_1457) );
OAI221xp5_ASAP7_75t_L g1299 ( .A1(n_1300), .A2(n_1303), .B1(n_1310), .B2(n_1313), .C(n_1314), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1302), .B(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1302), .Y(n_1391) );
OAI321xp33_ASAP7_75t_L g1383 ( .A1(n_1303), .A2(n_1371), .A3(n_1384), .B1(n_1385), .B2(n_1386), .C(n_1389), .Y(n_1383) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1304), .B(n_1378), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1306), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1305), .B(n_1369), .Y(n_1385) );
CKINVDCx6p67_ASAP7_75t_R g1312 ( .A(n_1306), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1306), .B(n_1349), .Y(n_1348) );
OAI221xp5_ASAP7_75t_L g1442 ( .A1(n_1306), .A2(n_1373), .B1(n_1439), .B2(n_1443), .C(n_1444), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1458 ( .A(n_1306), .B(n_1459), .Y(n_1458) );
OR2x6_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1309), .Y(n_1306) );
NOR2xp33_ASAP7_75t_L g1362 ( .A(n_1310), .B(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1311), .B(n_1343), .Y(n_1443) );
NAND2xp5_ASAP7_75t_L g1444 ( .A(n_1311), .B(n_1445), .Y(n_1444) );
AND2x4_ASAP7_75t_SL g1356 ( .A(n_1312), .B(n_1349), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1312), .B(n_1333), .Y(n_1369) );
OR2x2_ASAP7_75t_L g1396 ( .A(n_1312), .B(n_1349), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1312), .B(n_1417), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_1312), .B(n_1353), .Y(n_1422) );
NOR2xp33_ASAP7_75t_L g1436 ( .A(n_1312), .B(n_1437), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1312), .B(n_1426), .Y(n_1453) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1316), .Y(n_1314) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1319), .Y(n_1317) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1319), .Y(n_1425) );
NOR2xp33_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1331), .Y(n_1320) );
OAI31xp33_ASAP7_75t_L g1338 ( .A1(n_1321), .A2(n_1339), .A3(n_1360), .B(n_1362), .Y(n_1338) );
AOI221xp5_ASAP7_75t_L g1364 ( .A1(n_1321), .A2(n_1365), .B1(n_1369), .B2(n_1370), .C(n_1383), .Y(n_1364) );
BUFx3_ASAP7_75t_L g1426 ( .A(n_1321), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1447 ( .A(n_1321), .B(n_1331), .Y(n_1447) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1321), .Y(n_1459) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
NOR3xp33_ASAP7_75t_L g1357 ( .A(n_1331), .B(n_1358), .C(n_1359), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1408 ( .A(n_1331), .B(n_1375), .Y(n_1408) );
INVx2_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1332), .B(n_1342), .Y(n_1341) );
OAI322xp33_ASAP7_75t_L g1370 ( .A1(n_1332), .A2(n_1371), .A3(n_1373), .B1(n_1375), .B2(n_1376), .C1(n_1379), .C2(n_1380), .Y(n_1370) );
INVx2_ASAP7_75t_L g1378 ( .A(n_1332), .Y(n_1378) );
NAND3xp33_ASAP7_75t_L g1454 ( .A(n_1332), .B(n_1382), .C(n_1455), .Y(n_1454) );
INVx2_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
INVx2_ASAP7_75t_SL g1349 ( .A(n_1333), .Y(n_1349) );
OAI221xp5_ASAP7_75t_L g1339 ( .A1(n_1340), .A2(n_1343), .B1(n_1344), .B2(n_1347), .C(n_1350), .Y(n_1339) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1341), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1342), .B(n_1343), .Y(n_1464) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1343), .Y(n_1353) );
NOR2xp33_ASAP7_75t_L g1372 ( .A(n_1343), .B(n_1349), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1343), .B(n_1388), .Y(n_1387) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1344), .B(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
OAI21xp5_ASAP7_75t_L g1461 ( .A1(n_1345), .A2(n_1462), .B(n_1464), .Y(n_1461) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1346), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1346), .B(n_1382), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1424 ( .A(n_1346), .B(n_1368), .Y(n_1424) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1451 ( .A(n_1349), .B(n_1375), .Y(n_1451) );
AOI21xp5_ASAP7_75t_L g1350 ( .A1(n_1351), .A2(n_1356), .B(n_1357), .Y(n_1350) );
INVxp67_ASAP7_75t_SL g1351 ( .A(n_1352), .Y(n_1351) );
NAND3xp33_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1354), .C(n_1355), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1353), .B(n_1414), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1359), .B(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1361), .Y(n_1434) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1367), .Y(n_1452) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1369), .Y(n_1415) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
NOR2xp33_ASAP7_75t_L g1397 ( .A(n_1375), .B(n_1398), .Y(n_1397) );
O2A1O1Ixp33_ASAP7_75t_L g1450 ( .A1(n_1375), .A2(n_1395), .B(n_1426), .C(n_1451), .Y(n_1450) );
OAI221xp5_ASAP7_75t_L g1409 ( .A1(n_1376), .A2(n_1410), .B1(n_1411), .B2(n_1415), .C(n_1416), .Y(n_1409) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
NOR2xp33_ASAP7_75t_L g1417 ( .A(n_1384), .B(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
AOI31xp33_ASAP7_75t_L g1392 ( .A1(n_1393), .A2(n_1402), .A3(n_1419), .B(n_1426), .Y(n_1392) );
AOI21xp5_ASAP7_75t_L g1393 ( .A1(n_1394), .A2(n_1395), .B(n_1397), .Y(n_1393) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
O2A1O1Ixp33_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1404), .B(n_1407), .C(n_1409), .Y(n_1402) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
AOI21xp33_ASAP7_75t_L g1419 ( .A1(n_1420), .A2(n_1422), .B(n_1423), .Y(n_1419) );
OAI221xp5_ASAP7_75t_L g1456 ( .A1(n_1421), .A2(n_1457), .B1(n_1458), .B2(n_1460), .C(n_1461), .Y(n_1456) );
INVx2_ASAP7_75t_L g1437 ( .A(n_1426), .Y(n_1437) );
OAI221xp5_ASAP7_75t_SL g1427 ( .A1(n_1428), .A2(n_1435), .B1(n_1438), .B2(n_1439), .C(n_1441), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1430), .B(n_1432), .Y(n_1429) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
INVxp67_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
AOI21xp5_ASAP7_75t_SL g1441 ( .A1(n_1442), .A2(n_1446), .B(n_1448), .Y(n_1441) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
OAI221xp5_ASAP7_75t_L g1448 ( .A1(n_1449), .A2(n_1450), .B1(n_1452), .B2(n_1453), .C(n_1454), .Y(n_1448) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
HB1xp67_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1470), .Y(n_1563) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
INVx5_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
AND2x4_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1476), .Y(n_1473) );
INVx3_ASAP7_75t_L g1496 ( .A(n_1475), .Y(n_1496) );
NOR3xp33_ASAP7_75t_L g1477 ( .A(n_1478), .B(n_1492), .C(n_1501), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1487), .Y(n_1478) );
AOI22xp33_ASAP7_75t_L g1479 ( .A1(n_1480), .A2(n_1481), .B1(n_1484), .B2(n_1485), .Y(n_1479) );
OAI221xp5_ASAP7_75t_L g1552 ( .A1(n_1480), .A2(n_1490), .B1(n_1532), .B2(n_1553), .C(n_1555), .Y(n_1552) );
BUFx2_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
AND2x6_ASAP7_75t_L g1485 ( .A(n_1483), .B(n_1486), .Y(n_1485) );
NAND2x1p5_ASAP7_75t_L g1500 ( .A(n_1486), .B(n_1496), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g1487 ( .A1(n_1488), .A2(n_1489), .B1(n_1490), .B2(n_1491), .Y(n_1487) );
INVx2_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
INVx2_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
BUFx4f_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
BUFx2_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx2_ASAP7_75t_SL g1504 ( .A(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
OAI221xp5_ASAP7_75t_L g1529 ( .A1(n_1507), .A2(n_1509), .B1(n_1530), .B2(n_1532), .C(n_1534), .Y(n_1529) );
BUFx3_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
BUFx6f_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
INVx2_ASAP7_75t_SL g1532 ( .A(n_1533), .Y(n_1532) );
BUFx2_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_SL g1540 ( .A(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
AOI22xp33_ASAP7_75t_L g1545 ( .A1(n_1546), .A2(n_1548), .B1(n_1549), .B2(n_1551), .Y(n_1545) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
BUFx2_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
BUFx2_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVxp67_ASAP7_75t_SL g1568 ( .A(n_1569), .Y(n_1568) );
INVxp67_ASAP7_75t_L g1610 ( .A(n_1571), .Y(n_1610) );
HB1xp67_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
AND4x1_ASAP7_75t_L g1572 ( .A(n_1573), .B(n_1589), .C(n_1591), .D(n_1607), .Y(n_1572) );
INVx2_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
NOR2xp33_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1609), .Y(n_1607) );
endmodule