module fake_aes_452_n_1012 (n_117, n_44, n_133, n_149, n_81, n_69, n_214, n_204, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_96, n_39, n_1012);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_96;
input n_39;
output n_1012;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_230;
wire n_274;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_666;
wire n_621;
wire n_880;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_1006;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_859;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_991;
wire n_843;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g216 ( .A(n_84), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_209), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_52), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_158), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_109), .Y(n_220) );
BUFx5_ASAP7_75t_L g221 ( .A(n_142), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_92), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_98), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_20), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_200), .Y(n_225) );
BUFx3_ASAP7_75t_L g226 ( .A(n_28), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_201), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_137), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_165), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_189), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_35), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_12), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_49), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_85), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_102), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_103), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_205), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_134), .Y(n_238) );
BUFx10_ASAP7_75t_L g239 ( .A(n_204), .Y(n_239) );
INVxp33_ASAP7_75t_SL g240 ( .A(n_68), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_170), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_101), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_36), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_157), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_160), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_44), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_71), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_106), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_86), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_207), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_67), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_198), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_69), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_178), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_171), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_57), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_130), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_11), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_72), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_21), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_194), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_155), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_24), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_122), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_81), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_182), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_13), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_188), .Y(n_268) );
INVxp67_ASAP7_75t_SL g269 ( .A(n_192), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_166), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_186), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_27), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_73), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_58), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_196), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_120), .B(n_11), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_126), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_148), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_108), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_173), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_149), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_121), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_60), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_175), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_131), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_115), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_195), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_4), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_193), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_163), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_41), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_138), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_174), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_51), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_23), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_113), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_214), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_50), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_4), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_199), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_0), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_79), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_29), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_215), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_119), .B(n_104), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_168), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_10), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_78), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_20), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_51), .Y(n_310) );
CKINVDCx16_ASAP7_75t_R g311 ( .A(n_127), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_76), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_107), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_187), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_128), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_151), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_95), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_206), .Y(n_318) );
BUFx5_ASAP7_75t_L g319 ( .A(n_191), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_24), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_45), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_129), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_203), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_15), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_6), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_2), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_172), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_87), .Y(n_328) );
CKINVDCx14_ASAP7_75t_R g329 ( .A(n_66), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_31), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_52), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_70), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_88), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_59), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_190), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_222), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_218), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_230), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_217), .Y(n_339) );
CKINVDCx8_ASAP7_75t_R g340 ( .A(n_311), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_233), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_230), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_221), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_218), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_274), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_233), .B(n_1), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_246), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_246), .B(n_1), .Y(n_348) );
OA21x2_ASAP7_75t_L g349 ( .A1(n_223), .A2(n_65), .B(n_64), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_226), .B(n_2), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_226), .B(n_3), .Y(n_351) );
INVx4_ASAP7_75t_L g352 ( .A(n_227), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_241), .Y(n_353) );
OAI22x1_ASAP7_75t_R g354 ( .A1(n_224), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_354) );
INVx5_ASAP7_75t_L g355 ( .A(n_222), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_288), .A2(n_9), .B1(n_5), .B2(n_8), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_245), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_301), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_221), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_301), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_252), .Y(n_361) );
INVx6_ASAP7_75t_L g362 ( .A(n_239), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_291), .B(n_8), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_291), .A2(n_10), .B1(n_12), .B2(n_13), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_222), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_221), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_288), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_266), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_320), .B(n_14), .Y(n_369) );
AND2x6_ASAP7_75t_L g370 ( .A(n_249), .B(n_285), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_267), .B(n_14), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_341), .B(n_294), .Y(n_372) );
NAND2xp33_ASAP7_75t_L g373 ( .A(n_370), .B(n_221), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_343), .Y(n_374) );
NAND2xp33_ASAP7_75t_L g375 ( .A(n_370), .B(n_221), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_341), .A2(n_229), .B1(n_328), .B2(n_234), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_343), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_359), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
OR2x6_ASAP7_75t_L g380 ( .A(n_346), .B(n_232), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_350), .Y(n_381) );
AND2x6_ASAP7_75t_L g382 ( .A(n_350), .B(n_249), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_359), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_359), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g385 ( .A1(n_364), .A2(n_263), .B1(n_224), .B2(n_309), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_346), .A2(n_234), .B1(n_328), .B2(n_229), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_352), .B(n_318), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_350), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_366), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_351), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_352), .B(n_329), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_338), .B(n_260), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_366), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_352), .B(n_329), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_362), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_366), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_337), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
NAND2xp33_ASAP7_75t_SL g399 ( .A(n_347), .B(n_306), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_336), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_337), .Y(n_401) );
INVx4_ASAP7_75t_SL g402 ( .A(n_370), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_337), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_355), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_348), .A2(n_272), .B1(n_295), .B2(n_283), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_337), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_362), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_355), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_355), .Y(n_409) );
AND3x1_ASAP7_75t_L g410 ( .A(n_364), .B(n_303), .C(n_299), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_370), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_338), .B(n_239), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_342), .B(n_231), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_340), .B(n_219), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_344), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_362), .B(n_240), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_362), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_397), .Y(n_418) );
NAND2xp33_ASAP7_75t_L g419 ( .A(n_382), .B(n_370), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_391), .B(n_363), .Y(n_420) );
INVx4_ASAP7_75t_L g421 ( .A(n_382), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_397), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_382), .A2(n_351), .B1(n_363), .B2(n_367), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_380), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_394), .B(n_369), .Y(n_425) );
AO221x1_ASAP7_75t_L g426 ( .A1(n_376), .A2(n_354), .B1(n_353), .B2(n_357), .C(n_339), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_401), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_401), .Y(n_428) );
NOR2x1p5_ASAP7_75t_L g429 ( .A(n_372), .B(n_361), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_372), .B(n_368), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_382), .A2(n_367), .B1(n_344), .B2(n_370), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_380), .B(n_371), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_380), .A2(n_356), .B1(n_256), .B2(n_258), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_387), .B(n_345), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_392), .B(n_344), .Y(n_435) );
AND2x6_ASAP7_75t_SL g436 ( .A(n_380), .B(n_354), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_417), .B(n_235), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_413), .B(n_344), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_412), .B(n_345), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_403), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_416), .B(n_370), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_382), .B(n_370), .Y(n_442) );
NOR2x2_ASAP7_75t_L g443 ( .A(n_386), .B(n_263), .Y(n_443) );
NAND2x1_ASAP7_75t_L g444 ( .A(n_379), .B(n_349), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_379), .B(n_358), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_381), .B(n_360), .Y(n_446) );
NAND2x1_ASAP7_75t_L g447 ( .A(n_381), .B(n_349), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_415), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g450 ( .A(n_411), .B(n_298), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_381), .A2(n_388), .B(n_390), .Y(n_451) );
AOI22x1_ASAP7_75t_R g452 ( .A1(n_410), .A2(n_324), .B1(n_326), .B2(n_310), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_395), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_386), .B(n_321), .Y(n_455) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_411), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_381), .B(n_360), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_407), .Y(n_458) );
INVx2_ASAP7_75t_SL g459 ( .A(n_407), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_406), .Y(n_460) );
O2A1O1Ixp5_ASAP7_75t_L g461 ( .A1(n_388), .A2(n_269), .B(n_220), .C(n_225), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_390), .B(n_216), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_415), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_390), .A2(n_331), .B(n_330), .C(n_228), .Y(n_464) );
NOR2xp33_ASAP7_75t_SL g465 ( .A(n_411), .B(n_325), .Y(n_465) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_414), .B(n_349), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_377), .Y(n_467) );
OAI22xp33_ASAP7_75t_L g468 ( .A1(n_385), .A2(n_334), .B1(n_307), .B2(n_243), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_378), .Y(n_469) );
BUFx4_ASAP7_75t_L g470 ( .A(n_399), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_405), .B(n_236), .Y(n_471) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_374), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_389), .B(n_378), .Y(n_473) );
NAND2xp33_ASAP7_75t_L g474 ( .A(n_383), .B(n_319), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_402), .B(n_251), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_383), .B(n_237), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_384), .Y(n_477) );
OAI22xp33_ASAP7_75t_L g478 ( .A1(n_393), .A2(n_243), .B1(n_244), .B2(n_242), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_396), .Y(n_479) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_398), .B(n_247), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_398), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_404), .Y(n_482) );
NOR2xp67_ASAP7_75t_SL g483 ( .A(n_402), .B(n_255), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_404), .B(n_285), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_373), .A2(n_250), .B1(n_253), .B2(n_248), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_408), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_375), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_409), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_SL g489 ( .A1(n_409), .A2(n_276), .B(n_223), .C(n_238), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_400), .A2(n_257), .B1(n_259), .B2(n_254), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_400), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_444), .A2(n_262), .B(n_261), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_468), .A2(n_265), .B(n_268), .C(n_264), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_432), .B(n_271), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_424), .B(n_270), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_450), .B(n_273), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_430), .Y(n_497) );
NOR2x1_ASAP7_75t_L g498 ( .A(n_421), .B(n_275), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_424), .A2(n_277), .B1(n_279), .B2(n_278), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_472), .Y(n_500) );
CKINVDCx8_ASAP7_75t_R g501 ( .A(n_436), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_461), .A2(n_282), .B(n_284), .C(n_280), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_472), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_471), .A2(n_290), .B1(n_292), .B2(n_286), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_445), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_461), .A2(n_297), .B(n_304), .C(n_296), .Y(n_506) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_421), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_427), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_420), .B(n_287), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_441), .A2(n_312), .B(n_308), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_446), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_471), .A2(n_313), .B1(n_317), .B2(n_316), .Y(n_512) );
INVx5_ASAP7_75t_L g513 ( .A(n_456), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_425), .B(n_289), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_433), .A2(n_327), .B1(n_322), .B2(n_300), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_456), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_448), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_457), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g519 ( .A1(n_489), .A2(n_293), .B(n_335), .C(n_305), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_423), .A2(n_315), .B1(n_323), .B2(n_314), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_465), .B(n_332), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_454), .Y(n_522) );
AO32x2_ASAP7_75t_L g523 ( .A1(n_489), .A2(n_319), .A3(n_365), .B1(n_336), .B2(n_222), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_455), .B(n_16), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_460), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_429), .B(n_16), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_456), .Y(n_527) );
OR2x6_ASAP7_75t_SL g528 ( .A(n_443), .B(n_281), .Y(n_528) );
INVx4_ASAP7_75t_L g529 ( .A(n_456), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_434), .B(n_333), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_464), .A2(n_17), .B(n_18), .C(n_19), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_439), .B(n_319), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_462), .A2(n_355), .B(n_302), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_435), .Y(n_534) );
BUFx3_ASAP7_75t_L g535 ( .A(n_484), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_426), .B(n_18), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_439), .B(n_319), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_473), .B(n_438), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_477), .B(n_19), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_462), .A2(n_355), .B(n_302), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_476), .A2(n_418), .B(n_428), .C(n_422), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_431), .B(n_302), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_440), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_449), .Y(n_544) );
AO32x2_ASAP7_75t_L g545 ( .A1(n_453), .A2(n_458), .A3(n_459), .B1(n_488), .B2(n_482), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_437), .B(n_22), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_487), .A2(n_463), .B(n_419), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_476), .A2(n_365), .B1(n_336), .B2(n_27), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_467), .B(n_25), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_466), .A2(n_365), .B(n_336), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_442), .A2(n_479), .B(n_469), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_470), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_485), .B(n_25), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_478), .B(n_26), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_490), .A2(n_26), .B1(n_29), .B2(n_30), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_478), .B(n_32), .Y(n_556) );
OA22x2_ASAP7_75t_L g557 ( .A1(n_452), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_557) );
INVx3_ASAP7_75t_L g558 ( .A(n_481), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_486), .B(n_33), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_480), .B(n_34), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_475), .Y(n_561) );
OR2x6_ASAP7_75t_SL g562 ( .A(n_483), .B(n_37), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_474), .B(n_38), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_491), .B(n_39), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_423), .A2(n_40), .B1(n_41), .B2(n_42), .Y(n_565) );
INVx2_ASAP7_75t_SL g566 ( .A(n_430), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_423), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_432), .A2(n_45), .B1(n_46), .B2(n_47), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_472), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_455), .B(n_46), .Y(n_570) );
NOR2xp33_ASAP7_75t_R g571 ( .A(n_436), .B(n_47), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_468), .A2(n_48), .B1(n_49), .B2(n_53), .C(n_54), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_472), .Y(n_573) );
CKINVDCx14_ASAP7_75t_R g574 ( .A(n_430), .Y(n_574) );
OR2x6_ASAP7_75t_L g575 ( .A(n_424), .B(n_48), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_432), .B(n_53), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_430), .B(n_54), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_432), .B(n_55), .Y(n_578) );
AND2x4_ASAP7_75t_SL g579 ( .A(n_424), .B(n_55), .Y(n_579) );
OA22x2_ASAP7_75t_L g580 ( .A1(n_426), .A2(n_56), .B1(n_57), .B2(n_58), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_444), .A2(n_75), .B(n_74), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_423), .A2(n_56), .B1(n_59), .B2(n_60), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_444), .A2(n_146), .B(n_213), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_472), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_455), .B(n_61), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_432), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_432), .B(n_63), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_444), .A2(n_77), .B(n_80), .Y(n_588) );
OAI21xp33_ASAP7_75t_SL g589 ( .A1(n_472), .A2(n_82), .B(n_83), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_472), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_472), .Y(n_591) );
CKINVDCx8_ASAP7_75t_R g592 ( .A(n_436), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_421), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_423), .A2(n_89), .B1(n_90), .B2(n_91), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_500), .B(n_93), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_544), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g597 ( .A1(n_589), .A2(n_94), .B(n_96), .C(n_97), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_543), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_589), .B(n_99), .C(n_100), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_573), .B(n_105), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_550), .A2(n_110), .B(n_111), .Y(n_601) );
BUFx12f_ASAP7_75t_L g602 ( .A(n_575), .Y(n_602) );
AO31x2_ASAP7_75t_L g603 ( .A1(n_541), .A2(n_112), .A3(n_114), .B(n_116), .Y(n_603) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_575), .A2(n_117), .B1(n_118), .B2(n_123), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_547), .A2(n_124), .B(n_125), .Y(n_605) );
AOI221xp5_ASAP7_75t_SL g606 ( .A1(n_493), .A2(n_132), .B1(n_133), .B2(n_135), .C(n_136), .Y(n_606) );
BUFx8_ASAP7_75t_L g607 ( .A(n_536), .Y(n_607) );
NAND3x1_ASAP7_75t_L g608 ( .A(n_528), .B(n_139), .C(n_140), .Y(n_608) );
AOI211x1_ASAP7_75t_L g609 ( .A1(n_565), .A2(n_141), .B(n_143), .C(n_144), .Y(n_609) );
NAND2x1p5_ASAP7_75t_L g610 ( .A(n_552), .B(n_145), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_551), .A2(n_147), .B(n_150), .Y(n_611) );
AO31x2_ASAP7_75t_L g612 ( .A1(n_502), .A2(n_152), .A3(n_153), .B(n_154), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_567), .Y(n_613) );
AO31x2_ASAP7_75t_L g614 ( .A1(n_506), .A2(n_156), .A3(n_159), .B(n_161), .Y(n_614) );
AOI221xp5_ASAP7_75t_SL g615 ( .A1(n_577), .A2(n_162), .B1(n_164), .B2(n_167), .C(n_169), .Y(n_615) );
BUFx10_ASAP7_75t_L g616 ( .A(n_579), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_592), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_524), .B(n_176), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_510), .A2(n_177), .B(n_179), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_570), .B(n_180), .Y(n_620) );
AO22x2_ASAP7_75t_L g621 ( .A1(n_526), .A2(n_181), .B1(n_183), .B2(n_184), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_584), .B(n_185), .Y(n_622) );
INVx5_ASAP7_75t_L g623 ( .A(n_507), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_590), .A2(n_591), .B1(n_511), .B2(n_505), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_568), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_586), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_508), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_585), .B(n_197), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_517), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_522), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_525), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_539), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_574), .B(n_202), .Y(n_633) );
OAI22x1_ASAP7_75t_L g634 ( .A1(n_515), .A2(n_208), .B1(n_210), .B2(n_211), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_531), .A2(n_212), .B(n_587), .C(n_578), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_518), .B(n_495), .Y(n_636) );
AOI31xp67_ASAP7_75t_L g637 ( .A1(n_542), .A2(n_548), .A3(n_532), .B(n_537), .Y(n_637) );
AOI222xp33_ASAP7_75t_L g638 ( .A1(n_572), .A2(n_534), .B1(n_555), .B2(n_512), .C1(n_504), .C2(n_576), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_553), .A2(n_556), .B(n_554), .C(n_519), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_593), .B(n_535), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_499), .B(n_494), .Y(n_641) );
BUFx3_ASAP7_75t_L g642 ( .A(n_562), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_530), .A2(n_514), .B(n_509), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_557), .Y(n_644) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_581), .A2(n_588), .B(n_583), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_546), .B(n_559), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_549), .Y(n_647) );
NOR2xp67_ASAP7_75t_SL g648 ( .A(n_513), .B(n_507), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_558), .Y(n_649) );
OA21x2_ASAP7_75t_L g650 ( .A1(n_563), .A2(n_540), .B(n_533), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_520), .A2(n_580), .B1(n_560), .B2(n_498), .Y(n_651) );
INVx4_ASAP7_75t_SL g652 ( .A(n_571), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_561), .A2(n_496), .B(n_521), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_545), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_545), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_545), .Y(n_656) );
INVx3_ASAP7_75t_L g657 ( .A(n_529), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_564), .A2(n_593), .B(n_529), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_516), .A2(n_527), .B(n_523), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_516), .A2(n_527), .B(n_523), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_516), .A2(n_527), .B(n_523), .Y(n_661) );
AO32x2_ASAP7_75t_L g662 ( .A1(n_565), .A2(n_582), .A3(n_567), .B1(n_555), .B2(n_594), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_541), .A2(n_461), .B(n_451), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_544), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_500), .Y(n_665) );
NOR2xp67_ASAP7_75t_L g666 ( .A(n_566), .B(n_376), .Y(n_666) );
AO31x2_ASAP7_75t_L g667 ( .A1(n_541), .A2(n_506), .A3(n_502), .B(n_550), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_501), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_500), .Y(n_669) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_513), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_492), .A2(n_447), .B(n_444), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_500), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_492), .A2(n_447), .B(n_444), .Y(n_673) );
NOR2xp67_ASAP7_75t_L g674 ( .A(n_566), .B(n_376), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_500), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_500), .Y(n_676) );
AO31x2_ASAP7_75t_L g677 ( .A1(n_541), .A2(n_506), .A3(n_502), .B(n_550), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_500), .B(n_432), .Y(n_678) );
AOI21xp5_ASAP7_75t_SL g679 ( .A1(n_575), .A2(n_421), .B(n_472), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_500), .B(n_432), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_497), .Y(n_681) );
AO31x2_ASAP7_75t_L g682 ( .A1(n_541), .A2(n_506), .A3(n_502), .B(n_550), .Y(n_682) );
NAND3x1_ASAP7_75t_L g683 ( .A(n_536), .B(n_386), .C(n_364), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_497), .B(n_566), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_541), .A2(n_461), .B(n_451), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_497), .B(n_430), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_500), .A2(n_423), .B1(n_538), .B2(n_503), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_501), .Y(n_688) );
AO31x2_ASAP7_75t_L g689 ( .A1(n_541), .A2(n_506), .A3(n_502), .B(n_550), .Y(n_689) );
AND2x6_ASAP7_75t_L g690 ( .A(n_503), .B(n_569), .Y(n_690) );
NAND2x1p5_ASAP7_75t_L g691 ( .A(n_497), .B(n_552), .Y(n_691) );
AO31x2_ASAP7_75t_L g692 ( .A1(n_541), .A2(n_506), .A3(n_502), .B(n_550), .Y(n_692) );
AO31x2_ASAP7_75t_L g693 ( .A1(n_541), .A2(n_506), .A3(n_502), .B(n_550), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_686), .B(n_681), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_625), .B(n_626), .Y(n_695) );
AOI21x1_ASAP7_75t_L g696 ( .A1(n_659), .A2(n_661), .B(n_660), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_596), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_664), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_613), .B(n_598), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_627), .Y(n_700) );
BUFx2_ASAP7_75t_L g701 ( .A(n_691), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_636), .B(n_665), .Y(n_702) );
CKINVDCx11_ASAP7_75t_R g703 ( .A(n_652), .Y(n_703) );
OR2x6_ASAP7_75t_L g704 ( .A(n_679), .B(n_602), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_687), .B(n_641), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_669), .B(n_672), .Y(n_706) );
NAND2x1p5_ASAP7_75t_L g707 ( .A(n_648), .B(n_623), .Y(n_707) );
AOI21x1_ASAP7_75t_L g708 ( .A1(n_654), .A2(n_655), .B(n_656), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_624), .B(n_638), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_644), .A2(n_674), .B1(n_666), .B2(n_642), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_643), .A2(n_673), .B(n_671), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_675), .B(n_676), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_678), .B(n_680), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_623), .B(n_670), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_632), .B(n_647), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_629), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_621), .A2(n_620), .B1(n_628), .B2(n_618), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_630), .Y(n_718) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_631), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_690), .Y(n_720) );
NOR2x1_ASAP7_75t_R g721 ( .A(n_617), .B(n_668), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_649), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_690), .A2(n_607), .B1(n_646), .B2(n_621), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_651), .B(n_663), .Y(n_724) );
OA21x2_ASAP7_75t_L g725 ( .A1(n_615), .A2(n_606), .B(n_645), .Y(n_725) );
AND2x4_ASAP7_75t_L g726 ( .A(n_640), .B(n_657), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_688), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_599), .A2(n_683), .B1(n_604), .B2(n_597), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_640), .Y(n_729) );
CKINVDCx11_ASAP7_75t_R g730 ( .A(n_652), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_610), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_616), .B(n_633), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_608), .Y(n_733) );
OAI21x1_ASAP7_75t_SL g734 ( .A1(n_619), .A2(n_658), .B(n_595), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_600), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_667), .B(n_692), .Y(n_736) );
INVx4_ASAP7_75t_L g737 ( .A(n_650), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_667), .B(n_693), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_653), .B(n_622), .Y(n_739) );
OAI21x1_ASAP7_75t_L g740 ( .A1(n_611), .A2(n_601), .B(n_605), .Y(n_740) );
BUFx2_ASAP7_75t_L g741 ( .A(n_634), .Y(n_741) );
AO31x2_ASAP7_75t_L g742 ( .A1(n_637), .A2(n_603), .A3(n_609), .B(n_692), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_677), .B(n_692), .Y(n_743) );
O2A1O1Ixp33_ASAP7_75t_L g744 ( .A1(n_662), .A2(n_677), .B(n_682), .C(n_689), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_662), .A2(n_682), .B1(n_689), .B2(n_614), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_689), .B(n_612), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_662), .A2(n_612), .B1(n_614), .B2(n_603), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_614), .B(n_603), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_598), .Y(n_749) );
AOI21xp33_ASAP7_75t_SL g750 ( .A1(n_617), .A2(n_376), .B(n_580), .Y(n_750) );
BUFx2_ASAP7_75t_L g751 ( .A(n_681), .Y(n_751) );
AOI21x1_ASAP7_75t_L g752 ( .A1(n_659), .A2(n_661), .B(n_660), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_636), .B(n_644), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_598), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_598), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_598), .Y(n_756) );
BUFx6f_ASAP7_75t_L g757 ( .A(n_670), .Y(n_757) );
INVx3_ASAP7_75t_L g758 ( .A(n_623), .Y(n_758) );
AO21x2_ASAP7_75t_L g759 ( .A1(n_659), .A2(n_661), .B(n_660), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_598), .Y(n_760) );
OR2x2_ASAP7_75t_L g761 ( .A(n_686), .B(n_497), .Y(n_761) );
OAI21xp5_ASAP7_75t_L g762 ( .A1(n_663), .A2(n_685), .B(n_639), .Y(n_762) );
INVxp67_ASAP7_75t_SL g763 ( .A(n_636), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_625), .B(n_626), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_598), .Y(n_765) );
BUFx3_ASAP7_75t_L g766 ( .A(n_684), .Y(n_766) );
OA21x2_ASAP7_75t_L g767 ( .A1(n_659), .A2(n_661), .B(n_660), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_596), .Y(n_768) );
NAND2x1_ASAP7_75t_L g769 ( .A(n_648), .B(n_679), .Y(n_769) );
INVx2_ASAP7_75t_SL g770 ( .A(n_616), .Y(n_770) );
CKINVDCx6p67_ASAP7_75t_R g771 ( .A(n_602), .Y(n_771) );
INVx3_ASAP7_75t_L g772 ( .A(n_623), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_598), .Y(n_773) );
BUFx4f_ASAP7_75t_SL g774 ( .A(n_602), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_598), .Y(n_775) );
NOR2x1_ASAP7_75t_SL g776 ( .A(n_602), .B(n_575), .Y(n_776) );
AND2x4_ASAP7_75t_L g777 ( .A(n_636), .B(n_644), .Y(n_777) );
CKINVDCx6p67_ASAP7_75t_R g778 ( .A(n_602), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_596), .Y(n_779) );
INVx3_ASAP7_75t_L g780 ( .A(n_623), .Y(n_780) );
A2O1A1Ixp33_ASAP7_75t_L g781 ( .A1(n_643), .A2(n_639), .B(n_589), .C(n_635), .Y(n_781) );
NOR2x1_ASAP7_75t_SL g782 ( .A(n_602), .B(n_575), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_598), .Y(n_783) );
INVx4_ASAP7_75t_L g784 ( .A(n_602), .Y(n_784) );
INVx2_ASAP7_75t_SL g785 ( .A(n_616), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_596), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_684), .B(n_686), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_598), .Y(n_788) );
OA21x2_ASAP7_75t_L g789 ( .A1(n_762), .A2(n_748), .B(n_746), .Y(n_789) );
INVxp67_ASAP7_75t_L g790 ( .A(n_761), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_763), .B(n_697), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_737), .Y(n_792) );
INVx1_ASAP7_75t_SL g793 ( .A(n_751), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_709), .B(n_695), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_698), .B(n_768), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_709), .B(n_695), .Y(n_796) );
BUFx3_ASAP7_75t_L g797 ( .A(n_707), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_699), .Y(n_798) );
BUFx12f_ASAP7_75t_L g799 ( .A(n_703), .Y(n_799) );
INVx3_ASAP7_75t_L g800 ( .A(n_769), .Y(n_800) );
OR2x2_ASAP7_75t_L g801 ( .A(n_764), .B(n_713), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_733), .B(n_720), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_779), .B(n_786), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_708), .Y(n_804) );
AOI21x1_ASAP7_75t_L g805 ( .A1(n_696), .A2(n_752), .B(n_711), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_764), .B(n_787), .Y(n_806) );
OA21x2_ASAP7_75t_L g807 ( .A1(n_762), .A2(n_746), .B(n_747), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_713), .B(n_724), .Y(n_808) );
NOR2xp33_ASAP7_75t_SL g809 ( .A(n_774), .B(n_771), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_724), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_700), .B(n_716), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_718), .B(n_719), .Y(n_812) );
BUFx2_ASAP7_75t_L g813 ( .A(n_737), .Y(n_813) );
INVx3_ASAP7_75t_L g814 ( .A(n_757), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_749), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_715), .B(n_754), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_715), .B(n_755), .Y(n_817) );
OAI22xp33_ASAP7_75t_L g818 ( .A1(n_717), .A2(n_694), .B1(n_704), .B2(n_766), .Y(n_818) );
BUFx2_ASAP7_75t_L g819 ( .A(n_741), .Y(n_819) );
AOI21xp5_ASAP7_75t_SL g820 ( .A1(n_717), .A2(n_781), .B(n_705), .Y(n_820) );
OR2x2_ASAP7_75t_L g821 ( .A(n_705), .B(n_702), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_756), .B(n_760), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_765), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_773), .B(n_775), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_783), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_706), .B(n_712), .Y(n_826) );
BUFx3_ASAP7_75t_L g827 ( .A(n_707), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_788), .B(n_753), .Y(n_828) );
BUFx4f_ASAP7_75t_SL g829 ( .A(n_778), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_736), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_767), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_736), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_738), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_777), .B(n_723), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_722), .B(n_745), .Y(n_835) );
OR2x2_ASAP7_75t_L g836 ( .A(n_743), .B(n_780), .Y(n_836) );
OR2x6_ASAP7_75t_L g837 ( .A(n_704), .B(n_734), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_759), .Y(n_838) );
BUFx2_ASAP7_75t_L g839 ( .A(n_758), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_742), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_742), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_744), .Y(n_842) );
AND2x4_ASAP7_75t_L g843 ( .A(n_772), .B(n_780), .Y(n_843) );
BUFx2_ASAP7_75t_L g844 ( .A(n_701), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_725), .Y(n_845) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_729), .Y(n_846) );
OAI21xp5_ASAP7_75t_L g847 ( .A1(n_750), .A2(n_728), .B(n_739), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_735), .Y(n_848) );
INVx2_ASAP7_75t_SL g849 ( .A(n_714), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_740), .Y(n_850) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_726), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_804), .Y(n_852) );
OR2x2_ASAP7_75t_L g853 ( .A(n_836), .B(n_704), .Y(n_853) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_791), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_831), .Y(n_855) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_791), .Y(n_856) );
OR2x2_ASAP7_75t_L g857 ( .A(n_836), .B(n_710), .Y(n_857) );
BUFx3_ASAP7_75t_L g858 ( .A(n_813), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_835), .B(n_731), .Y(n_859) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_812), .Y(n_860) );
AO21x2_ASAP7_75t_L g861 ( .A1(n_805), .A2(n_732), .B(n_782), .Y(n_861) );
AND2x4_ASAP7_75t_L g862 ( .A(n_792), .B(n_776), .Y(n_862) );
OR2x2_ASAP7_75t_L g863 ( .A(n_821), .B(n_770), .Y(n_863) );
INVxp67_ASAP7_75t_L g864 ( .A(n_813), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_816), .B(n_785), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_830), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_832), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_812), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_816), .B(n_784), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_817), .B(n_784), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_817), .B(n_730), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_798), .B(n_721), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_810), .B(n_727), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_810), .B(n_833), .Y(n_874) );
AO21x2_ASAP7_75t_L g875 ( .A1(n_847), .A2(n_845), .B(n_850), .Y(n_875) );
BUFx2_ASAP7_75t_L g876 ( .A(n_792), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_822), .B(n_824), .Y(n_877) );
OR2x2_ASAP7_75t_L g878 ( .A(n_801), .B(n_808), .Y(n_878) );
NOR2x1_ASAP7_75t_L g879 ( .A(n_837), .B(n_797), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_822), .B(n_824), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_842), .B(n_798), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_808), .B(n_794), .Y(n_882) );
INVx2_ASAP7_75t_SL g883 ( .A(n_792), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_842), .B(n_815), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_815), .B(n_823), .Y(n_885) );
AND2x4_ASAP7_75t_L g886 ( .A(n_837), .B(n_800), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_823), .B(n_825), .Y(n_887) );
AND2x4_ASAP7_75t_L g888 ( .A(n_837), .B(n_800), .Y(n_888) );
INVx2_ASAP7_75t_SL g889 ( .A(n_797), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_811), .B(n_795), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_795), .B(n_803), .Y(n_891) );
OR2x2_ASAP7_75t_L g892 ( .A(n_801), .B(n_794), .Y(n_892) );
BUFx2_ASAP7_75t_L g893 ( .A(n_837), .Y(n_893) );
INVx3_ASAP7_75t_L g894 ( .A(n_886), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_855), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_877), .B(n_807), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_854), .A2(n_818), .B1(n_796), .B2(n_837), .Y(n_897) );
INVx5_ASAP7_75t_L g898 ( .A(n_862), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g899 ( .A(n_871), .B(n_809), .Y(n_899) );
INVxp67_ASAP7_75t_SL g900 ( .A(n_864), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_877), .B(n_807), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_852), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_881), .B(n_819), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_880), .B(n_807), .Y(n_904) );
AND2x4_ASAP7_75t_SL g905 ( .A(n_856), .B(n_800), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_884), .B(n_807), .Y(n_906) );
AND2x2_ASAP7_75t_SL g907 ( .A(n_893), .B(n_819), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_884), .B(n_820), .Y(n_908) );
OR2x2_ASAP7_75t_L g909 ( .A(n_860), .B(n_806), .Y(n_909) );
OR2x2_ASAP7_75t_L g910 ( .A(n_868), .B(n_826), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_891), .B(n_789), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_874), .B(n_820), .Y(n_912) );
BUFx2_ASAP7_75t_L g913 ( .A(n_858), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_891), .B(n_789), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_890), .B(n_789), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_874), .B(n_789), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_885), .B(n_840), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_885), .B(n_887), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_887), .B(n_841), .Y(n_919) );
INVxp67_ASAP7_75t_L g920 ( .A(n_869), .Y(n_920) );
NAND2xp33_ASAP7_75t_L g921 ( .A(n_879), .B(n_793), .Y(n_921) );
AND2x4_ASAP7_75t_L g922 ( .A(n_886), .B(n_838), .Y(n_922) );
NAND2xp5_ASAP7_75t_SL g923 ( .A(n_862), .B(n_839), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_866), .B(n_867), .Y(n_924) );
BUFx2_ASAP7_75t_L g925 ( .A(n_876), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_882), .A2(n_790), .B1(n_848), .B2(n_828), .C(n_846), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_895), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_896), .B(n_901), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_896), .B(n_883), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_918), .B(n_882), .Y(n_930) );
AND2x4_ASAP7_75t_L g931 ( .A(n_894), .B(n_888), .Y(n_931) );
INVx4_ASAP7_75t_L g932 ( .A(n_898), .Y(n_932) );
OR2x2_ASAP7_75t_L g933 ( .A(n_901), .B(n_878), .Y(n_933) );
NAND2x1_ASAP7_75t_L g934 ( .A(n_913), .B(n_879), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_902), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_904), .B(n_892), .Y(n_936) );
NAND2xp5_ASAP7_75t_SL g937 ( .A(n_898), .B(n_862), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_902), .Y(n_938) );
AND2x2_ASAP7_75t_SL g939 ( .A(n_905), .B(n_893), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_915), .B(n_911), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_918), .B(n_892), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_914), .B(n_875), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_914), .B(n_875), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_916), .B(n_875), .Y(n_944) );
OR2x6_ASAP7_75t_L g945 ( .A(n_913), .B(n_888), .Y(n_945) );
AND2x4_ASAP7_75t_L g946 ( .A(n_894), .B(n_888), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_903), .B(n_864), .Y(n_947) );
INVx1_ASAP7_75t_SL g948 ( .A(n_910), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_916), .B(n_875), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_906), .B(n_859), .Y(n_950) );
AND2x2_ASAP7_75t_SL g951 ( .A(n_905), .B(n_853), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_933), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_927), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_927), .Y(n_954) );
NAND2x1_ASAP7_75t_L g955 ( .A(n_932), .B(n_925), .Y(n_955) );
OR2x2_ASAP7_75t_L g956 ( .A(n_936), .B(n_903), .Y(n_956) );
AND2x2_ASAP7_75t_SL g957 ( .A(n_939), .B(n_905), .Y(n_957) );
OAI32xp33_ASAP7_75t_L g958 ( .A1(n_948), .A2(n_920), .A3(n_899), .B1(n_909), .B2(n_897), .Y(n_958) );
OR2x2_ASAP7_75t_L g959 ( .A(n_928), .B(n_908), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_928), .B(n_906), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_935), .Y(n_961) );
AOI21xp5_ASAP7_75t_L g962 ( .A1(n_937), .A2(n_921), .B(n_923), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_940), .B(n_917), .Y(n_963) );
OR2x2_ASAP7_75t_L g964 ( .A(n_941), .B(n_908), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_950), .B(n_912), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_940), .B(n_917), .Y(n_966) );
OR2x2_ASAP7_75t_L g967 ( .A(n_930), .B(n_919), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_942), .B(n_924), .Y(n_968) );
OAI21xp5_ASAP7_75t_L g969 ( .A1(n_939), .A2(n_870), .B(n_869), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_938), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_943), .B(n_922), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_970), .Y(n_972) );
OAI21xp5_ASAP7_75t_L g973 ( .A1(n_962), .A2(n_870), .B(n_939), .Y(n_973) );
AOI22xp5_ASAP7_75t_L g974 ( .A1(n_957), .A2(n_897), .B1(n_944), .B2(n_949), .Y(n_974) );
INVx2_ASAP7_75t_L g975 ( .A(n_953), .Y(n_975) );
OAI321xp33_ASAP7_75t_L g976 ( .A1(n_969), .A2(n_945), .A3(n_947), .B1(n_949), .B2(n_926), .C(n_872), .Y(n_976) );
INVx2_ASAP7_75t_L g977 ( .A(n_953), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_952), .B(n_929), .Y(n_978) );
AOI221x1_ASAP7_75t_L g979 ( .A1(n_961), .A2(n_932), .B1(n_873), .B2(n_848), .C(n_865), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_954), .Y(n_980) );
AOI21xp33_ASAP7_75t_L g981 ( .A1(n_958), .A2(n_861), .B(n_863), .Y(n_981) );
AOI21xp5_ASAP7_75t_L g982 ( .A1(n_955), .A2(n_951), .B(n_934), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_954), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_964), .A2(n_907), .B1(n_834), .B2(n_946), .Y(n_984) );
OAI21xp33_ASAP7_75t_L g985 ( .A1(n_974), .A2(n_958), .B(n_959), .Y(n_985) );
AOI32xp33_ASAP7_75t_L g986 ( .A1(n_976), .A2(n_960), .A3(n_963), .B1(n_966), .B2(n_932), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_973), .A2(n_955), .B1(n_951), .B2(n_956), .Y(n_987) );
OAI21xp5_ASAP7_75t_L g988 ( .A1(n_979), .A2(n_907), .B(n_951), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_981), .A2(n_965), .B1(n_971), .B2(n_968), .C(n_960), .Y(n_989) );
O2A1O1Ixp33_ASAP7_75t_SL g990 ( .A1(n_982), .A2(n_934), .B(n_967), .C(n_889), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_984), .A2(n_945), .B1(n_898), .B2(n_966), .Y(n_991) );
OAI21xp33_ASAP7_75t_SL g992 ( .A1(n_978), .A2(n_963), .B(n_945), .Y(n_992) );
NAND2xp5_ASAP7_75t_SL g993 ( .A(n_975), .B(n_898), .Y(n_993) );
AOI21xp33_ASAP7_75t_L g994 ( .A1(n_972), .A2(n_861), .B(n_865), .Y(n_994) );
OAI211xp5_ASAP7_75t_L g995 ( .A1(n_980), .A2(n_898), .B(n_900), .C(n_857), .Y(n_995) );
NAND3xp33_ASAP7_75t_L g996 ( .A(n_986), .B(n_989), .C(n_985), .Y(n_996) );
NOR3xp33_ASAP7_75t_L g997 ( .A(n_987), .B(n_992), .C(n_990), .Y(n_997) );
NOR3xp33_ASAP7_75t_L g998 ( .A(n_995), .B(n_991), .C(n_988), .Y(n_998) );
NAND3xp33_ASAP7_75t_SL g999 ( .A(n_997), .B(n_829), .C(n_799), .Y(n_999) );
AOI31xp33_ASAP7_75t_L g1000 ( .A1(n_996), .A2(n_799), .A3(n_994), .B(n_993), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_999), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g1002 ( .A(n_1001), .B(n_1000), .Y(n_1002) );
XNOR2xp5_ASAP7_75t_L g1003 ( .A(n_1001), .B(n_998), .Y(n_1003) );
XNOR2xp5_ASAP7_75t_L g1004 ( .A(n_1003), .B(n_851), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_1002), .B(n_977), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g1006 ( .A1(n_1005), .A2(n_861), .B1(n_802), .B2(n_844), .Y(n_1006) );
AOI21xp5_ASAP7_75t_L g1007 ( .A1(n_1004), .A2(n_843), .B(n_849), .Y(n_1007) );
AOI21xp5_ASAP7_75t_L g1008 ( .A1(n_1007), .A2(n_843), .B(n_849), .Y(n_1008) );
AOI22xp5_ASAP7_75t_L g1009 ( .A1(n_1006), .A2(n_802), .B1(n_843), .B2(n_827), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_1008), .B(n_931), .Y(n_1010) );
AO21x2_ASAP7_75t_L g1011 ( .A1(n_1010), .A2(n_1009), .B(n_983), .Y(n_1011) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_1011), .A2(n_983), .B(n_814), .Y(n_1012) );
endmodule