module fake_jpeg_8429_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_34),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_48),
.B1(n_18),
.B2(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_54),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_18),
.B1(n_33),
.B2(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_60),
.B1(n_47),
.B2(n_48),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_35),
.C(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx2_ASAP7_75t_SL g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_18),
.B1(n_33),
.B2(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g77 ( 
.A(n_61),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_64),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_21),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_35),
.B1(n_23),
.B2(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_75),
.Y(n_102)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_79),
.Y(n_120)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_85),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_94),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_46),
.Y(n_111)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_72),
.A2(n_80),
.B1(n_94),
.B2(n_48),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_123),
.B1(n_98),
.B2(n_84),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_31),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_112),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_67),
.B(n_38),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_43),
.C(n_45),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_22),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_22),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_89),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_39),
.B1(n_67),
.B2(n_46),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_89),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_137),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_39),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_154),
.C(n_114),
.Y(n_156)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_131),
.B(n_132),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_102),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_134),
.A2(n_143),
.B(n_146),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_136),
.A2(n_128),
.B1(n_141),
.B2(n_155),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_148),
.Y(n_158)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_68),
.B1(n_76),
.B2(n_87),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_141),
.A2(n_155),
.B1(n_105),
.B2(n_109),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_118),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_103),
.B(n_43),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_68),
.B1(n_76),
.B2(n_41),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_147),
.B1(n_115),
.B2(n_124),
.Y(n_165)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_41),
.B1(n_74),
.B2(n_25),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_22),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_107),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_151),
.B(n_152),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_103),
.A2(n_20),
.B(n_25),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_32),
.B(n_38),
.Y(n_153)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_99),
.B(n_45),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_41),
.C(n_52),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_36),
.B1(n_38),
.B2(n_19),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_156),
.B(n_186),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_170),
.Y(n_195)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_166),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_105),
.B1(n_99),
.B2(n_108),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_162),
.A2(n_167),
.B(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_178),
.B1(n_138),
.B2(n_152),
.Y(n_187)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_151),
.A2(n_126),
.B(n_125),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_179),
.B1(n_183),
.B2(n_147),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_177),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_118),
.C(n_121),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_185),
.C(n_56),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_136),
.B1(n_153),
.B2(n_144),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_143),
.B1(n_100),
.B2(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_0),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_105),
.B1(n_104),
.B2(n_74),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_113),
.Y(n_182)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_127),
.B1(n_122),
.B2(n_113),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_28),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_28),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_59),
.C(n_52),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_187),
.B(n_190),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_188),
.A2(n_189),
.B1(n_208),
.B2(n_165),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_143),
.B1(n_145),
.B2(n_100),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_184),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_202),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_205),
.B1(n_160),
.B2(n_169),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_199),
.C(n_201),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_100),
.B1(n_81),
.B2(n_61),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_198),
.A2(n_200),
.B1(n_207),
.B2(n_169),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_70),
.C(n_45),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_70),
.B1(n_17),
.B2(n_26),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_45),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_158),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_174),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_171),
.B1(n_183),
.B2(n_164),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_29),
.B1(n_30),
.B2(n_17),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_45),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_214),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_215),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_158),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_215),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_182),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_209),
.A2(n_171),
.B(n_164),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_221),
.B(n_237),
.Y(n_247)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_167),
.B(n_168),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_225),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_204),
.Y(n_223)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_235),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_234),
.B1(n_239),
.B2(n_201),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_193),
.A2(n_168),
.B1(n_163),
.B2(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_188),
.A2(n_176),
.B1(n_181),
.B2(n_29),
.Y(n_236)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_176),
.B(n_13),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_242),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_205),
.A2(n_192),
.B1(n_213),
.B2(n_207),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_196),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_194),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_216),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_255),
.Y(n_270)
);

XOR2x1_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_210),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_249),
.A2(n_259),
.B1(n_264),
.B2(n_32),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_220),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_252),
.A2(n_241),
.B1(n_233),
.B2(n_229),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_216),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_28),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_251),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_234),
.C(n_239),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_221),
.C(n_232),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_227),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_265),
.A2(n_231),
.B(n_240),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_276),
.C(n_281),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_255),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_274),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_218),
.B1(n_219),
.B2(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_223),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_219),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_275),
.B(n_247),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_32),
.C(n_28),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_252),
.A2(n_24),
.B1(n_30),
.B2(n_19),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_258),
.A2(n_26),
.B1(n_24),
.B2(n_19),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_26),
.B1(n_24),
.B2(n_28),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_0),
.C(n_1),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_0),
.C(n_1),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_265),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_3),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_247),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_270),
.C(n_10),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_283),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_256),
.Y(n_287)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_251),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_291),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_270),
.B(n_8),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_246),
.B1(n_253),
.B2(n_4),
.Y(n_295)
);

OAI321xp33_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_296),
.A3(n_3),
.B1(n_6),
.B2(n_8),
.C(n_9),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_289),
.Y(n_306)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_276),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_14),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_298),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_16),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_310),
.B(n_285),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_308),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_284),
.C(n_297),
.Y(n_310)
);

OAI21x1_ASAP7_75t_SL g311 ( 
.A1(n_285),
.A2(n_11),
.B(n_12),
.Y(n_311)
);

OR2x6_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_11),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_292),
.Y(n_313)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_319),
.B(n_303),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_320),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_12),
.B(n_14),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_307),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_312),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_310),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_327),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_313),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_314),
.B(n_321),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_331),
.A2(n_332),
.B(n_323),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_330),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_316),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_326),
.B(n_306),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_15),
.B(n_330),
.Y(n_340)
);


endmodule