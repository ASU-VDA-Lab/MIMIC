module fake_netlist_5_1020_n_7696 (n_137, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_649, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_631, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_637, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_645, n_539, n_175, n_538, n_262, n_238, n_639, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_7696);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_639;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_7696;

wire n_924;
wire n_6643;
wire n_6122;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_977;
wire n_4706;
wire n_5567;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_6579;
wire n_7164;
wire n_5287;
wire n_6546;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_790;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_5978;
wire n_2395;
wire n_5161;
wire n_5776;
wire n_6551;
wire n_5512;
wire n_5207;
wire n_2347;
wire n_6786;
wire n_7206;
wire n_7303;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_7461;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_6649;
wire n_7154;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_6810;
wire n_7660;
wire n_671;
wire n_6276;
wire n_6072;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_7686;
wire n_4211;
wire n_7024;
wire n_3448;
wire n_7205;
wire n_6742;
wire n_3019;
wire n_2096;
wire n_6694;
wire n_877;
wire n_3776;
wire n_7616;
wire n_2530;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_7486;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_6090;
wire n_6580;
wire n_7010;
wire n_5480;
wire n_6549;
wire n_668;
wire n_6913;
wire n_2147;
wire n_3010;
wire n_7315;
wire n_7004;
wire n_2770;
wire n_4131;
wire n_5402;
wire n_2584;
wire n_5851;
wire n_3188;
wire n_5509;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_7641;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_1242;
wire n_3283;
wire n_7468;
wire n_5469;
wire n_2323;
wire n_6431;
wire n_5744;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_731;
wire n_5202;
wire n_5648;
wire n_7667;
wire n_1314;
wire n_1512;
wire n_6931;
wire n_1490;
wire n_6618;
wire n_6408;
wire n_3214;
wire n_7523;
wire n_1517;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_5922;
wire n_1449;
wire n_6698;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_5848;
wire n_5406;
wire n_6085;
wire n_3947;
wire n_3490;
wire n_7421;
wire n_7306;
wire n_6214;
wire n_7493;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_6939;
wire n_882;
wire n_2384;
wire n_7528;
wire n_3156;
wire n_696;
wire n_3376;
wire n_7562;
wire n_5037;
wire n_4468;
wire n_5661;
wire n_6991;
wire n_3653;
wire n_5562;
wire n_3702;
wire n_1040;
wire n_4976;
wire n_6586;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_6096;
wire n_2276;
wire n_6707;
wire n_5852;
wire n_2089;
wire n_3420;
wire n_6920;
wire n_6868;
wire n_1561;
wire n_1165;
wire n_5144;
wire n_1034;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_845;
wire n_7402;
wire n_4255;
wire n_1796;
wire n_5577;
wire n_901;
wire n_4484;
wire n_7592;
wire n_3668;
wire n_7152;
wire n_6512;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_5689;
wire n_5894;
wire n_2079;
wire n_2238;
wire n_1151;
wire n_1405;
wire n_7463;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_6725;
wire n_7613;
wire n_2859;
wire n_1075;
wire n_3395;
wire n_7083;
wire n_4917;
wire n_7086;
wire n_7349;
wire n_6464;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_7647;
wire n_5825;
wire n_2968;
wire n_7316;
wire n_1585;
wire n_6820;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_4421;
wire n_6098;
wire n_7019;
wire n_6686;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_6561;
wire n_6584;
wire n_7452;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3735;
wire n_3349;
wire n_7323;
wire n_2248;
wire n_7195;
wire n_6701;
wire n_7478;
wire n_3007;
wire n_1000;
wire n_6769;
wire n_7683;
wire n_6592;
wire n_5686;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_6191;
wire n_6062;
wire n_2258;
wire n_748;
wire n_1667;
wire n_1058;
wire n_838;
wire n_3983;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_5909;
wire n_1385;
wire n_7575;
wire n_793;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_6043;
wire n_2987;
wire n_1527;
wire n_6271;
wire n_7171;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_6793;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_7127;
wire n_5397;
wire n_4471;
wire n_6550;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_5709;
wire n_7568;
wire n_3208;
wire n_6021;
wire n_3331;
wire n_4983;
wire n_2379;
wire n_5695;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_5860;
wire n_6926;
wire n_3649;
wire n_4302;
wire n_7589;
wire n_6928;
wire n_2514;
wire n_5862;
wire n_6304;
wire n_5189;
wire n_6956;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_7026;
wire n_1027;
wire n_4160;
wire n_6782;
wire n_2293;
wire n_5854;
wire n_5516;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_7002;
wire n_1412;
wire n_3981;
wire n_7141;
wire n_5936;
wire n_6126;
wire n_1199;
wire n_1038;
wire n_1841;
wire n_6027;
wire n_6598;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_6342;
wire n_1711;
wire n_870;
wire n_6638;
wire n_1891;
wire n_7308;
wire n_5254;
wire n_3526;
wire n_6900;
wire n_2546;
wire n_965;
wire n_3790;
wire n_7264;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_7457;
wire n_4613;
wire n_4649;
wire n_7617;
wire n_1888;
wire n_6269;
wire n_5615;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_5902;
wire n_4028;
wire n_5479;
wire n_1690;
wire n_3819;
wire n_6013;
wire n_7357;
wire n_2449;
wire n_5083;
wire n_6927;
wire n_1194;
wire n_6503;
wire n_5888;
wire n_2297;
wire n_4186;
wire n_7310;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_5698;
wire n_5592;
wire n_7521;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_7593;
wire n_6256;
wire n_2876;
wire n_4099;
wire n_7406;
wire n_7600;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_5870;
wire n_1464;
wire n_4295;
wire n_5303;
wire n_1444;
wire n_7076;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_6982;
wire n_1680;
wire n_4697;
wire n_7286;
wire n_7137;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_6727;
wire n_3317;
wire n_7539;
wire n_1121;
wire n_7229;
wire n_4391;
wire n_949;
wire n_5954;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1001;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_6097;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_7125;
wire n_6677;
wire n_1195;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_6624;
wire n_7121;
wire n_2796;
wire n_757;
wire n_6466;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_6008;
wire n_3095;
wire n_2805;
wire n_1145;
wire n_5624;
wire n_4918;
wire n_5714;
wire n_5806;
wire n_3856;
wire n_1153;
wire n_741;
wire n_7624;
wire n_4898;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_6221;
wire n_7160;
wire n_4002;
wire n_1163;
wire n_6805;
wire n_6185;
wire n_1207;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_6568;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_6004;
wire n_940;
wire n_6351;
wire n_7552;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_6901;
wire n_2947;
wire n_978;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_4801;
wire n_7183;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_6411;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_3378;
wire n_5435;
wire n_1431;
wire n_6873;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_5745;
wire n_7139;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_6594;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_962;
wire n_723;
wire n_2536;
wire n_6387;
wire n_1336;
wire n_7223;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_6179;
wire n_7338;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_6019;
wire n_6222;
wire n_7165;
wire n_3505;
wire n_6223;
wire n_4610;
wire n_6435;
wire n_3730;
wire n_4489;
wire n_7235;
wire n_974;
wire n_727;
wire n_5210;
wire n_6976;
wire n_4967;
wire n_6486;
wire n_5657;
wire n_957;
wire n_6889;
wire n_6083;
wire n_4992;
wire n_6844;
wire n_3001;
wire n_7404;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_6295;
wire n_3597;
wire n_1612;
wire n_4198;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_5857;
wire n_4534;
wire n_4500;
wire n_7437;
wire n_5014;
wire n_6241;
wire n_3185;
wire n_1300;
wire n_6087;
wire n_1127;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_6846;
wire n_4329;
wire n_1006;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_5756;
wire n_2231;
wire n_6041;
wire n_2017;
wire n_2604;
wire n_6994;
wire n_4257;
wire n_3453;
wire n_7449;
wire n_7329;
wire n_2390;
wire n_5708;
wire n_3213;
wire n_6790;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_7194;
wire n_6273;
wire n_3474;
wire n_3984;
wire n_6807;
wire n_5927;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3888;
wire n_3422;
wire n_5638;
wire n_7115;
wire n_4189;
wire n_5670;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_5584;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_5965;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_948;
wire n_5751;
wire n_5664;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_5641;
wire n_4037;
wire n_6218;
wire n_7281;
wire n_2922;
wire n_3499;
wire n_3275;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_6824;
wire n_1552;
wire n_6189;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_6993;
wire n_3683;
wire n_6037;
wire n_7245;
wire n_3642;
wire n_3808;
wire n_3286;
wire n_5963;
wire n_5980;
wire n_824;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_815;
wire n_4594;
wire n_6153;
wire n_3424;
wire n_5970;
wire n_1381;
wire n_6418;
wire n_1037;
wire n_6564;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_7192;
wire n_3171;
wire n_6671;
wire n_1437;
wire n_6591;
wire n_6266;
wire n_7161;
wire n_7580;
wire n_7153;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_6517;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_7350;
wire n_5690;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_6967;
wire n_5885;
wire n_2254;
wire n_6433;
wire n_1382;
wire n_925;
wire n_3546;
wire n_7535;
wire n_6893;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_950;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_7178;
wire n_7480;
wire n_2443;
wire n_1811;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_7632;
wire n_3244;
wire n_6501;
wire n_6028;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_968;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_5362;
wire n_6709;
wire n_4355;
wire n_3494;
wire n_6798;
wire n_5702;
wire n_5050;
wire n_885;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_683;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_721;
wire n_4572;
wire n_3073;
wire n_1157;
wire n_5527;
wire n_6986;
wire n_802;
wire n_5609;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_5266;
wire n_7471;
wire n_3178;
wire n_873;
wire n_5355;
wire n_2334;
wire n_6745;
wire n_690;
wire n_4521;
wire n_4488;
wire n_5977;
wire n_6811;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_6209;
wire n_2263;
wire n_6875;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_6853;
wire n_4519;
wire n_5551;
wire n_7594;
wire n_3715;
wire n_7340;
wire n_6699;
wire n_6073;
wire n_972;
wire n_5767;
wire n_6324;
wire n_3040;
wire n_1938;
wire n_5640;
wire n_2499;
wire n_1200;
wire n_3568;
wire n_5655;
wire n_5475;
wire n_3737;
wire n_1185;
wire n_991;
wire n_6138;
wire n_7603;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_5692;
wire n_4856;
wire n_7494;
wire n_2997;
wire n_5921;
wire n_4400;
wire n_5168;
wire n_943;
wire n_3326;
wire n_6477;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_883;
wire n_6159;
wire n_6283;
wire n_7396;
wire n_5322;
wire n_856;
wire n_7116;
wire n_1793;
wire n_4352;
wire n_7519;
wire n_4441;
wire n_6943;
wire n_918;
wire n_4761;
wire n_6827;
wire n_6173;
wire n_942;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_6312;
wire n_2533;
wire n_2364;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_6997;
wire n_5418;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_1096;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_7664;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_6300;
wire n_2043;
wire n_2751;
wire n_6131;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_6537;
wire n_5933;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_7023;
wire n_1807;
wire n_2618;
wire n_7428;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_763;
wire n_6783;
wire n_4748;
wire n_7465;
wire n_2295;
wire n_3931;
wire n_1219;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_7149;
wire n_2795;
wire n_6459;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_5644;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_6869;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_7117;
wire n_789;
wire n_4247;
wire n_4933;
wire n_6977;
wire n_4018;
wire n_3900;
wire n_1105;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_6313;
wire n_3872;
wire n_4336;
wire n_6569;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_6555;
wire n_3877;
wire n_6639;
wire n_7516;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_1102;
wire n_7596;
wire n_4052;
wire n_5864;
wire n_6536;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_6490;
wire n_2633;
wire n_6961;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_1164;
wire n_2097;
wire n_5460;
wire n_7628;
wire n_4304;
wire n_6761;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_6294;
wire n_6767;
wire n_4431;
wire n_7427;
wire n_4192;
wire n_6802;
wire n_7527;
wire n_5570;
wire n_3736;
wire n_6326;
wire n_4805;
wire n_4885;
wire n_5983;
wire n_1661;
wire n_5804;
wire n_6376;
wire n_3565;
wire n_6167;
wire n_4701;
wire n_2575;
wire n_5910;
wire n_7411;
wire n_7101;
wire n_5040;
wire n_6730;
wire n_6948;
wire n_861;
wire n_6582;
wire n_1658;
wire n_1904;
wire n_6996;
wire n_1345;
wire n_1899;
wire n_6974;
wire n_6765;
wire n_7577;
wire n_1003;
wire n_6921;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_1726;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_6898;
wire n_6710;
wire n_5717;
wire n_7162;
wire n_5464;
wire n_6565;
wire n_1657;
wire n_5886;
wire n_768;
wire n_7080;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3639;
wire n_7302;
wire n_6533;
wire n_708;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_6960;
wire n_6426;
wire n_6634;
wire n_7180;
wire n_1915;
wire n_5610;
wire n_1109;
wire n_5239;
wire n_6836;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_6972;
wire n_2924;
wire n_7111;
wire n_7549;
wire n_4111;
wire n_808;
wire n_2484;
wire n_797;
wire n_5785;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_6344;
wire n_5305;
wire n_5994;
wire n_4538;
wire n_6093;
wire n_766;
wire n_6010;
wire n_7247;
wire n_1117;
wire n_6833;
wire n_2754;
wire n_687;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_7481;
wire n_5204;
wire n_7292;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_7150;
wire n_2866;
wire n_3561;
wire n_7687;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_6265;
wire n_1650;
wire n_1137;
wire n_6821;
wire n_3934;
wire n_4985;
wire n_6373;
wire n_6988;
wire n_5788;
wire n_3922;
wire n_3846;
wire n_7692;
wire n_5897;
wire n_6887;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_1999;
wire n_6676;
wire n_2372;
wire n_3673;
wire n_6347;
wire n_6492;
wire n_7016;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_5795;
wire n_7072;
wire n_5508;
wire n_5582;
wire n_4022;
wire n_7374;
wire n_7440;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_7547;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_7201;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_5746;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_6648;
wire n_4601;
wire n_2687;
wire n_1120;
wire n_1890;
wire n_714;
wire n_4220;
wire n_1944;
wire n_909;
wire n_5630;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_7513;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_7413;
wire n_4403;
wire n_1981;
wire n_7540;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_5504;
wire n_7622;
wire n_7005;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_7353;
wire n_6219;
wire n_1889;
wire n_6965;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_6720;
wire n_1569;
wire n_2188;
wire n_6032;
wire n_7174;
wire n_6205;
wire n_6362;
wire n_6402;
wire n_756;
wire n_1429;
wire n_4644;
wire n_7166;
wire n_4456;
wire n_5060;
wire n_7607;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_7591;
wire n_5775;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_7282;
wire n_6491;
wire n_2898;
wire n_2717;
wire n_7151;
wire n_6229;
wire n_1861;
wire n_760;
wire n_5731;
wire n_5581;
wire n_3628;
wire n_3691;
wire n_6668;
wire n_7446;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_7053;
wire n_5831;
wire n_2573;
wire n_7473;
wire n_4435;
wire n_2939;
wire n_6835;
wire n_6419;
wire n_6039;
wire n_3807;
wire n_5884;
wire n_2447;
wire n_4764;
wire n_886;
wire n_5653;
wire n_6258;
wire n_7070;
wire n_1221;
wire n_5394;
wire n_6755;
wire n_2774;
wire n_7276;
wire n_7351;
wire n_1707;
wire n_853;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_751;
wire n_6084;
wire n_4827;
wire n_7412;
wire n_7157;
wire n_6436;
wire n_2488;
wire n_7666;
wire n_6472;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_704;
wire n_7211;
wire n_4399;
wire n_6531;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_771;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_7368;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_6567;
wire n_5889;
wire n_6771;
wire n_2526;
wire n_6389;
wire n_2703;
wire n_2167;
wire n_5764;
wire n_5428;
wire n_6910;
wire n_6442;
wire n_3391;
wire n_6102;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_6441;
wire n_5543;
wire n_816;
wire n_5678;
wire n_5935;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_7677;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_5950;
wire n_2173;
wire n_1842;
wire n_871;
wire n_3738;
wire n_685;
wire n_5995;
wire n_6162;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_6331;
wire n_1555;
wire n_6006;
wire n_3245;
wire n_4417;
wire n_6109;
wire n_6278;
wire n_6787;
wire n_6872;
wire n_4899;
wire n_796;
wire n_6208;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_6632;
wire n_1012;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_7027;
wire n_3509;
wire n_3352;
wire n_5671;
wire n_3076;
wire n_6990;
wire n_3535;
wire n_2182;
wire n_6349;
wire n_3251;
wire n_1061;
wire n_2931;
wire n_7631;
wire n_6830;
wire n_5185;
wire n_1193;
wire n_6359;
wire n_3118;
wire n_3511;
wire n_1226;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_7498;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_7377;
wire n_781;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_6301;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_5945;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_6744;
wire n_4981;
wire n_3125;
wire n_3114;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_6439;
wire n_7381;
wire n_5565;
wire n_4081;
wire n_1103;
wire n_3132;
wire n_4407;
wire n_7291;
wire n_3951;
wire n_4894;
wire n_5780;
wire n_5643;
wire n_3238;
wire n_3210;
wire n_5846;
wire n_2036;
wire n_7430;
wire n_3267;
wire n_4995;
wire n_695;
wire n_5524;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_6104;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_6475;
wire n_3884;
wire n_6465;
wire n_3726;
wire n_6496;
wire n_805;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_6998;
wire n_6145;
wire n_3577;
wire n_2820;
wire n_7305;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_3347;
wire n_1074;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_7075;
wire n_7545;
wire n_1448;
wire n_4288;
wire n_6076;
wire n_3567;
wire n_6194;
wire n_7695;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_6092;
wire n_7275;
wire n_5401;
wire n_6357;
wire n_5843;
wire n_4241;
wire n_3321;
wire n_7537;
wire n_3212;
wire n_666;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_7489;
wire n_5106;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_6335;
wire n_1186;
wire n_5883;
wire n_6985;
wire n_5319;
wire n_1018;
wire n_2247;
wire n_7451;
wire n_6238;
wire n_713;
wire n_1622;
wire n_1180;
wire n_3705;
wire n_6548;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_2268;
wire n_3778;
wire n_5706;
wire n_5337;
wire n_6366;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_7236;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_7269;
wire n_5223;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_6602;
wire n_4419;
wire n_4477;
wire n_6620;
wire n_3179;
wire n_6502;
wire n_3256;
wire n_7560;
wire n_667;
wire n_7326;
wire n_7060;
wire n_2386;
wire n_1501;
wire n_7572;
wire n_3086;
wire n_1007;
wire n_6885;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_1099;
wire n_2568;
wire n_5364;
wire n_6529;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_1021;
wire n_5895;
wire n_4639;
wire n_6951;
wire n_3713;
wire n_3663;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_7169;
wire n_6423;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_7140;
wire n_7233;
wire n_819;
wire n_5088;
wire n_2302;
wire n_6558;
wire n_5457;
wire n_7352;
wire n_951;
wire n_7134;
wire n_5532;
wire n_1494;
wire n_2069;
wire n_6950;
wire n_7246;
wire n_6525;
wire n_7650;
wire n_3434;
wire n_1806;
wire n_933;
wire n_6631;
wire n_6892;
wire n_1563;
wire n_7663;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_755;
wire n_7056;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_6683;
wire n_2482;
wire n_2677;
wire n_6292;
wire n_5544;
wire n_3832;
wire n_3987;
wire n_7339;
wire n_902;
wire n_5987;
wire n_6180;
wire n_5352;
wire n_5824;
wire n_4991;
wire n_5538;
wire n_6658;
wire n_6264;
wire n_6925;
wire n_5919;
wire n_1698;
wire n_2329;
wire n_1098;
wire n_2142;
wire n_6176;
wire n_5410;
wire n_3332;
wire n_7146;
wire n_1135;
wire n_3048;
wire n_3937;
wire n_6124;
wire n_7672;
wire n_2203;
wire n_4525;
wire n_1243;
wire n_3782;
wire n_7482;
wire n_6864;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_7090;
wire n_3786;
wire n_7158;
wire n_2888;
wire n_7156;
wire n_5742;
wire n_3638;
wire n_5992;
wire n_6494;
wire n_5503;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_6199;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_5958;
wire n_6614;
wire n_3022;
wire n_4264;
wire n_7504;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_7360;
wire n_7681;
wire n_7301;
wire n_5129;
wire n_2149;
wire n_1078;
wire n_7375;
wire n_7102;
wire n_5500;
wire n_3060;
wire n_4276;
wire n_7366;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_5654;
wire n_2408;
wire n_7025;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_6947;
wire n_1723;
wire n_5107;
wire n_5999;
wire n_4485;
wire n_7309;
wire n_4626;
wire n_1036;
wire n_1097;
wire n_6863;
wire n_6637;
wire n_798;
wire n_6100;
wire n_6735;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_6358;
wire n_1852;
wire n_5602;
wire n_3089;
wire n_6050;
wire n_2470;
wire n_7244;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_1391;
wire n_670;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_7610;
wire n_663;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_5903;
wire n_6371;
wire n_813;
wire n_1284;
wire n_7043;
wire n_3440;
wire n_6171;
wire n_6510;
wire n_1748;
wire n_4569;
wire n_6468;
wire n_2699;
wire n_4897;
wire n_888;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_2615;
wire n_3940;
wire n_1064;
wire n_5842;
wire n_858;
wire n_6352;
wire n_2985;
wire n_691;
wire n_5722;
wire n_7534;
wire n_5636;
wire n_5065;
wire n_2753;
wire n_7287;
wire n_1582;
wire n_7032;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_5492;
wire n_3141;
wire n_5084;
wire n_6850;
wire n_5667;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_7119;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_6354;
wire n_5918;
wire n_7634;
wire n_4503;
wire n_3507;
wire n_6959;
wire n_3821;
wire n_6909;
wire n_2700;
wire n_1211;
wire n_6332;
wire n_3367;
wire n_4464;
wire n_7006;
wire n_5877;
wire n_907;
wire n_3096;
wire n_6306;
wire n_7682;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_6434;
wire n_2356;
wire n_6751;
wire n_7068;
wire n_892;
wire n_4556;
wire n_6322;
wire n_5454;
wire n_2620;
wire n_6667;
wire n_7526;
wire n_1581;
wire n_6530;
wire n_4089;
wire n_7376;
wire n_6156;
wire n_5913;
wire n_7268;
wire n_7044;
wire n_5621;
wire n_2919;
wire n_4327;
wire n_953;
wire n_4218;
wire n_6429;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_7239;
wire n_2757;
wire n_963;
wire n_1052;
wire n_954;
wire n_5573;
wire n_6405;
wire n_6613;
wire n_4353;
wire n_2042;
wire n_6248;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_6088;
wire n_5529;
wire n_6894;
wire n_1856;
wire n_7267;
wire n_4959;
wire n_4161;
wire n_5800;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_6204;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_1156;
wire n_794;
wire n_7387;
wire n_7431;
wire n_7654;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_686;
wire n_2837;
wire n_847;
wire n_4844;
wire n_6296;
wire n_2979;
wire n_5257;
wire n_6290;
wire n_6288;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_702;
wire n_2548;
wire n_822;
wire n_5645;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_5779;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_6140;
wire n_1779;
wire n_7441;
wire n_4738;
wire n_6211;
wire n_1369;
wire n_3909;
wire n_6307;
wire n_6164;
wire n_3207;
wire n_3944;
wire n_7394;
wire n_809;
wire n_4434;
wire n_4837;
wire n_7022;
wire n_3042;
wire n_1942;
wire n_6860;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_5697;
wire n_7188;
wire n_1810;
wire n_7573;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_7087;
wire n_2222;
wire n_3510;
wire n_6147;
wire n_3218;
wire n_2667;
wire n_6515;
wire n_6011;
wire n_6645;
wire n_3150;
wire n_747;
wire n_6984;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_851;
wire n_843;
wire n_7193;
wire n_705;
wire n_3775;
wire n_4133;
wire n_6897;
wire n_7256;
wire n_678;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_6460;
wire n_4379;
wire n_7128;
wire n_7595;
wire n_2181;
wire n_1829;
wire n_6183;
wire n_7522;
wire n_5882;
wire n_4030;
wire n_7436;
wire n_4490;
wire n_3138;
wire n_7380;
wire n_7012;
wire n_4397;
wire n_1710;
wire n_7502;
wire n_1128;
wire n_2928;
wire n_7335;
wire n_7103;
wire n_1734;
wire n_4820;
wire n_6246;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_6383;
wire n_4938;
wire n_7020;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_677;
wire n_2723;
wire n_5672;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_5548;
wire n_5601;
wire n_7248;
wire n_7662;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_6099;
wire n_3158;
wire n_5693;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_6904;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_7533;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_878;
wire n_6626;
wire n_6563;
wire n_5486;
wire n_6611;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_5599;
wire n_906;
wire n_6116;
wire n_919;
wire n_7186;
wire n_4356;
wire n_6819;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_6473;
wire n_1586;
wire n_4291;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_6310;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_7429;
wire n_3545;
wire n_6688;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_1614;
wire n_2339;
wire n_7148;
wire n_5782;
wire n_6714;
wire n_4637;
wire n_7017;
wire n_7250;
wire n_7462;
wire n_7658;
wire n_4935;
wire n_6365;
wire n_4785;
wire n_3820;
wire n_3454;
wire n_3426;
wire n_5608;
wire n_3741;
wire n_3410;
wire n_7401;
wire n_6828;
wire n_2029;
wire n_995;
wire n_1609;
wire n_5298;
wire n_6355;
wire n_5596;
wire n_1887;
wire n_4413;
wire n_1073;
wire n_6777;
wire n_5728;
wire n_2346;
wire n_662;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_1215;
wire n_1592;
wire n_6420;
wire n_6945;
wire n_2882;
wire n_1721;
wire n_7356;
wire n_2338;
wire n_5726;
wire n_7288;
wire n_7637;
wire n_7124;
wire n_3672;
wire n_7294;
wire n_5290;
wire n_3197;
wire n_7018;
wire n_3109;
wire n_2721;
wire n_7321;
wire n_1043;
wire n_5095;
wire n_3002;
wire n_6754;
wire n_6583;
wire n_6622;
wire n_6936;
wire n_5324;
wire n_3897;
wire n_1159;
wire n_7691;
wire n_5928;
wire n_3845;
wire n_7108;
wire n_6882;
wire n_2081;
wire n_7585;
wire n_4570;
wire n_7386;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_5911;
wire n_7362;
wire n_7417;
wire n_2418;
wire n_7187;
wire n_5589;
wire n_5841;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_7544;
wire n_3458;
wire n_5712;
wire n_1420;
wire n_3330;
wire n_1132;
wire n_4606;
wire n_6166;
wire n_4774;
wire n_2477;
wire n_6966;
wire n_3887;
wire n_7542;
wire n_6781;
wire n_7255;
wire n_4093;
wire n_1486;
wire n_7120;
wire n_7218;
wire n_4672;
wire n_7147;
wire n_3519;
wire n_7221;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_4766;
wire n_5633;
wire n_2896;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_6980;
wire n_1927;
wire n_5583;
wire n_1349;
wire n_4460;
wire n_3645;
wire n_1031;
wire n_3223;
wire n_3929;
wire n_6064;
wire n_6110;
wire n_6237;
wire n_834;
wire n_7196;
wire n_2255;
wire n_2272;
wire n_893;
wire n_6341;
wire n_1965;
wire n_1902;
wire n_6590;
wire n_1941;
wire n_5501;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_6697;
wire n_874;
wire n_5652;
wire n_6453;
wire n_6135;
wire n_7559;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_7081;
wire n_3189;
wire n_2066;
wire n_6449;
wire n_993;
wire n_3154;
wire n_1551;
wire n_6141;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_7584;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_6983;
wire n_970;
wire n_1935;
wire n_6036;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_7222;
wire n_3242;
wire n_6071;
wire n_3525;
wire n_3486;
wire n_6808;
wire n_2405;
wire n_6724;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_4036;
wire n_6571;
wire n_921;
wire n_5100;
wire n_7470;
wire n_1795;
wire n_5849;
wire n_6251;
wire n_7400;
wire n_2578;
wire n_3483;
wire n_6635;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_1080;
wire n_1274;
wire n_7623;
wire n_3524;
wire n_5616;
wire n_7597;
wire n_5034;
wire n_6733;
wire n_1708;
wire n_7071;
wire n_5988;
wire n_6467;
wire n_6035;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_6522;
wire n_7109;
wire n_2092;
wire n_5959;
wire n_2075;
wire n_7645;
wire n_3658;
wire n_6732;
wire n_1776;
wire n_4807;
wire n_6562;
wire n_6150;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_890;
wire n_1919;
wire n_960;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_5917;
wire n_1252;
wire n_5754;
wire n_6016;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_7212;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_5628;
wire n_1808;
wire n_6726;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_7009;
wire n_6554;
wire n_967;
wire n_6689;
wire n_2731;
wire n_6143;
wire n_5614;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_7355;
wire n_3979;
wire n_7365;
wire n_4582;
wire n_2998;
wire n_6277;
wire n_4684;
wire n_7395;
wire n_5981;
wire n_6095;
wire n_7671;
wire n_6247;
wire n_4840;
wire n_3162;
wire n_983;
wire n_2760;
wire n_6880;
wire n_3377;
wire n_3749;
wire n_5720;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_762;
wire n_1283;
wire n_5325;
wire n_5696;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_6499;
wire n_6837;
wire n_4423;
wire n_4096;
wire n_7393;
wire n_2881;
wire n_6616;
wire n_1203;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_6946;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_5759;
wire n_4478;
wire n_5753;
wire n_2646;
wire n_5536;
wire n_1605;
wire n_7484;
wire n_5173;
wire n_6305;
wire n_1228;
wire n_6317;
wire n_3920;
wire n_4890;
wire n_5691;
wire n_5794;
wire n_5027;
wire n_5647;
wire n_7231;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_7272;
wire n_828;
wire n_779;
wire n_4106;
wire n_3717;
wire n_5738;
wire n_2743;
wire n_2675;
wire n_7649;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_7324;
wire n_945;
wire n_6693;
wire n_3743;
wire n_6734;
wire n_7135;
wire n_7014;
wire n_1932;
wire n_4721;
wire n_5597;
wire n_5635;
wire n_984;
wire n_694;
wire n_6382;
wire n_7328;
wire n_1983;
wire n_7635;
wire n_6404;
wire n_5975;
wire n_4029;
wire n_1594;
wire n_900;
wire n_3870;
wire n_6379;
wire n_7066;
wire n_4496;
wire n_3529;
wire n_7358;
wire n_1977;
wire n_1147;
wire n_2153;
wire n_6235;
wire n_4338;
wire n_7277;
wire n_6504;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_7265;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_6789;
wire n_7184;
wire n_6440;
wire n_6417;
wire n_1470;
wire n_2318;
wire n_1735;
wire n_833;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_7491;
wire n_5942;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_1201;
wire n_7690;
wire n_1114;
wire n_7219;
wire n_7479;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_669;
wire n_7270;
wire n_1176;
wire n_5940;
wire n_1149;
wire n_7390;
wire n_1020;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_5555;
wire n_6914;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_7182;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_5784;
wire n_6272;
wire n_6484;
wire n_661;
wire n_7674;
wire n_6236;
wire n_5576;
wire n_4668;
wire n_4953;
wire n_5466;
wire n_6958;
wire n_6840;
wire n_3898;
wire n_849;
wire n_6871;
wire n_1786;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_6768;
wire n_4759;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_7506;
wire n_2340;
wire n_3552;
wire n_875;
wire n_6717;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_7048;
wire n_5578;
wire n_2361;
wire n_1173;
wire n_1603;
wire n_1401;
wire n_969;
wire n_4113;
wire n_1998;
wire n_1019;
wire n_4686;
wire n_5530;
wire n_3759;
wire n_6196;
wire n_7416;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_5741;
wire n_5991;
wire n_3933;
wire n_7330;
wire n_3206;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_1702;
wire n_5221;
wire n_6992;
wire n_4183;
wire n_778;
wire n_4068;
wire n_1122;
wire n_4872;
wire n_6000;
wire n_4233;
wire n_7283;
wire n_3192;
wire n_7099;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_6448;
wire n_2649;
wire n_6655;
wire n_7304;
wire n_5792;
wire n_1187;
wire n_6657;
wire n_1929;
wire n_5575;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_1174;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_7626;
wire n_3742;
wire n_7474;
wire n_2252;
wire n_7612;
wire n_6113;
wire n_4819;
wire n_1685;
wire n_917;
wire n_1714;
wire n_6242;
wire n_7088;
wire n_6519;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_6842;
wire n_7588;
wire n_3390;
wire n_1573;
wire n_6206;
wire n_6414;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_6801;
wire n_774;
wire n_2493;
wire n_4930;
wire n_7680;
wire n_5276;
wire n_6308;
wire n_1059;
wire n_7398;
wire n_1133;
wire n_6906;
wire n_5078;
wire n_4537;
wire n_7230;
wire n_2885;
wire n_6629;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_6968;
wire n_4282;
wire n_6615;
wire n_3485;
wire n_4180;
wire n_7378;
wire n_665;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_5651;
wire n_2845;
wire n_6144;
wire n_4143;
wire n_4659;
wire n_6188;
wire n_2602;
wire n_5819;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_5998;
wire n_6398;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_5721;
wire n_5673;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_6415;
wire n_2994;
wire n_6857;
wire n_2401;
wire n_3135;
wire n_5476;
wire n_2003;
wire n_5856;
wire n_1457;
wire n_5446;
wire n_4895;
wire n_6722;
wire n_3573;
wire n_3148;
wire n_6428;
wire n_5944;
wire n_7618;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_6413;
wire n_7679;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_6361;
wire n_3438;
wire n_6231;
wire n_4098;
wire n_872;
wire n_5684;
wire n_5861;
wire n_1297;
wire n_5976;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_2184;
wire n_1184;
wire n_5312;
wire n_985;
wire n_5850;
wire n_3404;
wire n_3425;
wire n_3217;
wire n_5111;
wire n_5890;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_7167;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_7643;
wire n_676;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_6712;
wire n_1602;
wire n_1178;
wire n_5687;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_5839;
wire n_3397;
wire n_3740;
wire n_6953;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_703;
wire n_1318;
wire n_780;
wire n_2977;
wire n_6303;
wire n_6474;
wire n_6182;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_5674;
wire n_3600;
wire n_6573;
wire n_4134;
wire n_6053;
wire n_7234;
wire n_1388;
wire n_2836;
wire n_5682;
wire n_672;
wire n_6392;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_3239;
wire n_898;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_5612;
wire n_6125;
wire n_6599;
wire n_6685;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_6560;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_6253;
wire n_4740;
wire n_7382;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_7615;
wire n_5898;
wire n_1192;
wire n_2221;
wire n_3576;
wire n_1024;
wire n_7298;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_7581;
wire n_4049;
wire n_6641;
wire n_941;
wire n_3862;
wire n_5214;
wire n_5563;
wire n_5487;
wire n_6593;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_6673;
wire n_7172;
wire n_7074;
wire n_5497;
wire n_4724;
wire n_5832;
wire n_1238;
wire n_7190;
wire n_7112;
wire n_7678;
wire n_1772;
wire n_752;
wire n_1476;
wire n_1108;
wire n_5526;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_6367;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_6195;
wire n_862;
wire n_3584;
wire n_6356;
wire n_3756;
wire n_2889;
wire n_7001;
wire n_5593;
wire n_5021;
wire n_6514;
wire n_2772;
wire n_7369;
wire n_5444;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_6559;
wire n_7359;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_7144;
wire n_4833;
wire n_6841;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_5110;
wire n_6653;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_7450;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_5737;
wire n_786;
wire n_1142;
wire n_2579;
wire n_6923;
wire n_6825;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_6112;
wire n_2788;
wire n_6547;
wire n_2984;
wire n_6198;
wire n_7439;
wire n_3364;
wire n_5560;
wire n_6399;
wire n_1873;
wire n_3201;
wire n_6275;
wire n_1087;
wire n_5666;
wire n_6575;
wire n_3472;
wire n_6151;
wire n_2874;
wire n_5179;
wire n_7227;
wire n_7040;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_7325;
wire n_4968;
wire n_6469;
wire n_6756;
wire n_1272;
wire n_5030;
wire n_3949;
wire n_5961;
wire n_3543;
wire n_7191;
wire n_1247;
wire n_7459;
wire n_7096;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_5272;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_6826;
wire n_2360;
wire n_6015;
wire n_3254;
wire n_5361;
wire n_5683;
wire n_4171;
wire n_5847;
wire n_7551;
wire n_4045;
wire n_6678;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_5740;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_5729;
wire n_7485;
wire n_6748;
wire n_2030;
wire n_903;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_6752;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_6553;
wire n_2209;
wire n_7652;
wire n_6500;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_7051;
wire n_5152;
wire n_2321;
wire n_722;
wire n_3680;
wire n_6628;
wire n_844;
wire n_6297;
wire n_5905;
wire n_3497;
wire n_6975;
wire n_1601;
wire n_5409;
wire n_6329;
wire n_2940;
wire n_7536;
wire n_5688;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_979;
wire n_2841;
wire n_6293;
wire n_3322;
wire n_4576;
wire n_846;
wire n_2505;
wire n_2427;
wire n_7676;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_7553;
wire n_6905;
wire n_7425;
wire n_2594;
wire n_5798;
wire n_6381;
wire n_6521;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_5986;
wire n_3112;
wire n_2349;
wire n_6581;
wire n_1379;
wire n_3874;
wire n_6215;
wire n_7095;
wire n_5415;
wire n_4676;
wire n_5770;
wire n_7064;
wire n_5892;
wire n_4544;
wire n_2170;
wire n_1091;
wire n_6577;
wire n_6899;
wire n_5676;
wire n_7307;
wire n_6545;
wire n_5802;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_6370;
wire n_3266;
wire n_7210;
wire n_4646;
wire n_5769;
wire n_6065;
wire n_1130;
wire n_7039;
wire n_6987;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_6190;
wire n_6859;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_6309;
wire n_6623;
wire n_2426;
wire n_6527;
wire n_7443;
wire n_5341;
wire n_4320;
wire n_5930;
wire n_5814;
wire n_4881;
wire n_5979;
wire n_5271;
wire n_5089;
wire n_7015;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1505;
wire n_1181;
wire n_6929;
wire n_4012;
wire n_5518;
wire n_4636;
wire n_5637;
wire n_4584;
wire n_5622;
wire n_807;
wire n_3910;
wire n_4711;
wire n_835;
wire n_3319;
wire n_7348;
wire n_5240;
wire n_3335;
wire n_5813;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_5546;
wire n_927;
wire n_2689;
wire n_3259;
wire n_7143;
wire n_5482;
wire n_7312;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_7155;
wire n_3688;
wire n_6865;
wire n_3016;
wire n_1693;
wire n_5393;
wire n_2599;
wire n_6535;
wire n_904;
wire n_3338;
wire n_7213;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_5966;
wire n_1542;
wire n_7456;
wire n_5041;
wire n_7420;
wire n_1423;
wire n_1166;
wire n_1751;
wire n_5431;
wire n_1508;
wire n_785;
wire n_2200;
wire n_3261;
wire n_6482;
wire n_5026;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_5059;
wire n_5505;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_6605;
wire n_4250;
wire n_5329;
wire n_1055;
wire n_3596;
wire n_4699;
wire n_7007;
wire n_3906;
wire n_4127;
wire n_880;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_6018;
wire n_5908;
wire n_4202;
wire n_7168;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_688;
wire n_5939;
wire n_7177;
wire n_3766;
wire n_1353;
wire n_800;
wire n_2880;
wire n_7379;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_7444;
wire n_5931;
wire n_7435;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_915;
wire n_864;
wire n_7030;
wire n_5420;
wire n_1264;
wire n_6311;
wire n_4412;
wire n_3599;
wire n_3407;
wire n_6424;
wire n_6654;
wire n_6816;
wire n_6220;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_6740;
wire n_7122;
wire n_5835;
wire n_7049;
wire n_7567;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_6029;
wire n_1607;
wire n_6879;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_1118;
wire n_1686;
wire n_5679;
wire n_947;
wire n_3710;
wire n_5938;
wire n_6702;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_5891;
wire n_1230;
wire n_4144;
wire n_5724;
wire n_5774;
wire n_2165;
wire n_6452;
wire n_929;
wire n_3379;
wire n_4374;
wire n_6791;
wire n_3532;
wire n_1124;
wire n_5131;
wire n_7280;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_6915;
wire n_7110;
wire n_1104;
wire n_1294;
wire n_7511;
wire n_1257;
wire n_6856;
wire n_1182;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_7232;
wire n_4548;
wire n_7345;
wire n_5923;
wire n_5790;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_6451;
wire n_6364;
wire n_6552;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_6328;
wire n_4816;
wire n_1483;
wire n_6363;
wire n_2983;
wire n_7159;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_6132;
wire n_6578;
wire n_6406;
wire n_5598;
wire n_2085;
wire n_1669;
wire n_5306;
wire n_6978;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_2651;
wire n_4358;
wire n_7477;
wire n_5147;
wire n_3656;
wire n_6918;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_7363;
wire n_6612;
wire n_5677;
wire n_4168;
wire n_3446;
wire n_5997;
wire n_955;
wire n_5511;
wire n_5680;
wire n_3028;
wire n_4806;
wire n_4350;
wire n_1146;
wire n_7295;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_897;
wire n_5280;
wire n_6375;
wire n_6479;
wire n_1428;
wire n_6866;
wire n_1216;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_6170;
wire n_1931;
wire n_4187;
wire n_1070;
wire n_4166;
wire n_6447;
wire n_6263;
wire n_7093;
wire n_5206;
wire n_1030;
wire n_3222;
wire n_1071;
wire n_7466;
wire n_1267;
wire n_1801;
wire n_5419;
wire n_6130;
wire n_1513;
wire n_2970;
wire n_7651;
wire n_2235;
wire n_673;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_680;
wire n_1473;
wire n_3755;
wire n_5803;
wire n_4258;
wire n_6014;
wire n_4498;
wire n_6935;
wire n_1590;
wire n_7530;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_675;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_5985;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_6907;
wire n_6158;
wire n_7661;
wire n_6541;
wire n_3262;
wire n_6119;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_5896;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_889;
wire n_2358;
wire n_973;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_6226;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_7145;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_6338;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_7467;
wire n_736;
wire n_5097;
wire n_2750;
wire n_5730;
wire n_3899;
wire n_7550;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_5816;
wire n_4069;
wire n_2784;
wire n_7541;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_7241;
wire n_2557;
wire n_5300;
wire n_1248;
wire n_4850;
wire n_6625;
wire n_3781;
wire n_4912;
wire n_4813;
wire n_7464;
wire n_2590;
wire n_6302;
wire n_2330;
wire n_5748;
wire n_2942;
wire n_6759;
wire n_5525;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_6706;
wire n_944;
wire n_3889;
wire n_6139;
wire n_4256;
wire n_7434;
wire n_7636;
wire n_7054;
wire n_6999;
wire n_4224;
wire n_6403;
wire n_3508;
wire n_6483;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_6228;
wire n_857;
wire n_5650;
wire n_2636;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_7299;
wire n_4702;
wire n_6888;
wire n_4252;
wire n_4457;
wire n_6063;
wire n_971;
wire n_6800;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_6922;
wire n_3481;
wire n_5481;
wire n_6890;
wire n_7503;
wire n_2808;
wire n_6070;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_6651;
wire n_5821;
wire n_7091;
wire n_4491;
wire n_7273;
wire n_6647;
wire n_7296;
wire n_2930;
wire n_5733;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_5871;
wire n_7543;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_6184;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_7507;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_7555;
wire n_5707;
wire n_4001;
wire n_3047;
wire n_868;
wire n_2454;
wire n_4371;
wire n_5836;
wire n_914;
wire n_5281;
wire n_6716;
wire n_6422;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5521;
wire n_7578;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_7475;
wire n_4194;
wire n_759;
wire n_5585;
wire n_6397;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_7033;
wire n_6121;
wire n_1571;
wire n_3119;
wire n_7531;
wire n_4142;
wire n_4082;
wire n_1189;
wire n_5561;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_6981;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_6954;
wire n_3279;
wire n_2621;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_5875;
wire n_4262;
wire n_2671;
wire n_6646;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_7131;
wire n_6903;
wire n_1647;
wire n_4685;
wire n_6101;
wire n_5968;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_6941;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_5812;
wire n_6148;
wire n_5515;
wire n_6106;
wire n_6604;
wire n_4014;
wire n_7418;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_7688;
wire n_2913;
wire n_2336;
wire n_1233;
wire n_5607;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_6566;
wire n_1443;
wire n_946;
wire n_1539;
wire n_5734;
wire n_6081;
wire n_4892;
wire n_7204;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_689;
wire n_738;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_1279;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_6047;
wire n_2960;
wire n_1090;
wire n_5438;
wire n_4627;
wire n_758;
wire n_7354;
wire n_7448;
wire n_6244;
wire n_2290;
wire n_6861;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_1049;
wire n_2145;
wire n_5725;
wire n_1639;
wire n_3030;
wire n_1068;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_7571;
wire n_5163;
wire n_2039;
wire n_5768;
wire n_4961;
wire n_7556;
wire n_3753;
wire n_7640;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_7422;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_6588;
wire n_3396;
wire n_1445;
wire n_7050;
wire n_4023;
wire n_4420;
wire n_5685;
wire n_1923;
wire n_5773;
wire n_7136;
wire n_7318;
wire n_6055;
wire n_5138;
wire n_1017;
wire n_5374;
wire n_6108;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_6165;
wire n_1828;
wire n_6621;
wire n_2320;
wire n_1045;
wire n_7175;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_6323;
wire n_1033;
wire n_4396;
wire n_5127;
wire n_6587;
wire n_4367;
wire n_6480;
wire n_2087;
wire n_6731;
wire n_5485;
wire n_5766;
wire n_5216;
wire n_6597;
wire n_1009;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_6933;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_6881;
wire n_1578;
wire n_7289;
wire n_5805;
wire n_7665;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_6216;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_6817;
wire n_7170;
wire n_7314;
wire n_2725;
wire n_6949;
wire n_6509;
wire n_5175;
wire n_3883;
wire n_7260;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_773;
wire n_7263;
wire n_743;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_6911;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_5900;
wire n_3466;
wire n_4962;
wire n_1237;
wire n_6327;
wire n_2595;
wire n_761;
wire n_6607;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_7509;
wire n_7209;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_6401;
wire n_5554;
wire n_6227;
wire n_7240;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_5427;
wire n_5639;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_5417;
wire n_4614;
wire n_1265;
wire n_2681;
wire n_3103;
wire n_765;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_7609;
wire n_1015;
wire n_7278;
wire n_1651;
wire n_7630;
wire n_2775;
wire n_6416;
wire n_4693;
wire n_5488;
wire n_1101;
wire n_4326;
wire n_1106;
wire n_6695;
wire n_3557;
wire n_2230;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_6127;
wire n_7565;
wire n_2851;
wire n_4305;
wire n_5781;
wire n_1455;
wire n_6600;
wire n_767;
wire n_2490;
wire n_1407;
wire n_7410;
wire n_4213;
wire n_2849;
wire n_7097;
wire n_3692;
wire n_2204;
wire n_6421;
wire n_5747;
wire n_7414;
wire n_7495;
wire n_5969;
wire n_4929;
wire n_729;
wire n_1961;
wire n_4964;
wire n_911;
wire n_1430;
wire n_6079;
wire n_4802;
wire n_6192;
wire n_6458;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_6746;
wire n_2508;
wire n_4031;
wire n_7586;
wire n_6719;
wire n_2416;
wire n_5437;
wire n_5826;
wire n_7659;
wire n_3881;
wire n_2461;
wire n_6506;
wire n_2243;
wire n_4583;
wire n_6287;
wire n_6662;
wire n_4210;
wire n_5245;
wire n_7189;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_6851;
wire n_6687;
wire n_2890;
wire n_6884;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_716;
wire n_1630;
wire n_6780;
wire n_6513;
wire n_4891;
wire n_6619;
wire n_701;
wire n_1023;
wire n_5603;
wire n_6804;
wire n_803;
wire n_1092;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_5716;
wire n_3993;
wire n_4940;
wire n_6516;
wire n_5208;
wire n_7490;
wire n_1056;
wire n_3588;
wire n_6924;
wire n_2308;
wire n_4590;
wire n_7492;
wire n_5606;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_1029;
wire n_1206;
wire n_5456;
wire n_3160;
wire n_7073;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_6040;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_5727;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_7114;
wire n_1060;
wire n_5347;
wire n_2824;
wire n_3298;
wire n_3033;
wire n_6788;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_6393;
wire n_2333;
wire n_2916;
wire n_6249;
wire n_4297;
wire n_5833;
wire n_6849;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_7271;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_6572;
wire n_4172;
wire n_4791;
wire n_6739;
wire n_4536;
wire n_5149;
wire n_5967;
wire n_2463;
wire n_5151;
wire n_7569;
wire n_7003;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_6666;
wire n_2472;
wire n_4611;
wire n_6812;
wire n_4755;
wire n_5982;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_7419;
wire n_5827;
wire n_1560;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_6200;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_6123;
wire n_6934;
wire n_2589;
wire n_7094;
wire n_7500;
wire n_1301;
wire n_1363;
wire n_3482;
wire n_6082;
wire n_2233;
wire n_1312;
wire n_804;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_1504;
wire n_7129;
wire n_3956;
wire n_5758;
wire n_5323;
wire n_3572;
wire n_992;
wire n_4215;
wire n_6952;
wire n_4280;
wire n_7062;
wire n_3375;
wire n_4047;
wire n_5471;
wire n_842;
wire n_7642;
wire n_5434;
wire n_2082;
wire n_5941;
wire n_7045;
wire n_1643;
wire n_5879;
wire n_3167;
wire n_5558;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_7238;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_7126;
wire n_5669;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3078;
wire n_6979;
wire n_6203;
wire n_7405;
wire n_894;
wire n_3253;
wire n_7207;
wire n_4027;
wire n_831;
wire n_2280;
wire n_7454;
wire n_4599;
wire n_5830;
wire n_6796;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_5760;
wire n_6368;
wire n_3689;
wire n_6556;
wire n_2020;
wire n_4628;
wire n_5668;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_5878;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_5765;
wire n_3950;
wire n_4458;
wire n_6596;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_6870;
wire n_7639;
wire n_4476;
wire n_5613;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_7251;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_6080;
wire n_7059;
wire n_7035;
wire n_1848;
wire n_5571;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_6713;
wire n_5513;
wire n_6747;
wire n_6281;
wire n_4803;
wire n_5972;
wire n_4079;
wire n_4091;
wire n_681;
wire n_1638;
wire n_5916;
wire n_5984;
wire n_7029;
wire n_7317;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_6094;
wire n_2935;
wire n_6444;
wire n_5132;
wire n_830;
wire n_5191;
wire n_6333;
wire n_6262;
wire n_3085;
wire n_5869;
wire n_5925;
wire n_1655;
wire n_749;
wire n_6240;
wire n_5359;
wire n_6412;
wire n_2574;
wire n_1134;
wire n_5293;
wire n_1358;
wire n_7220;
wire n_717;
wire n_4316;
wire n_3697;
wire n_939;
wire n_7438;
wire n_1232;
wire n_734;
wire n_2638;
wire n_7515;
wire n_7574;
wire n_4044;
wire n_4062;
wire n_6684;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_7065;
wire n_1338;
wire n_5510;
wire n_6046;
wire n_2016;
wire n_1522;
wire n_6973;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_7285;
wire n_5200;
wire n_1653;
wire n_5659;
wire n_1506;
wire n_5618;
wire n_6325;
wire n_990;
wire n_2867;
wire n_1894;
wire n_975;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_6737;
wire n_6454;
wire n_4253;
wire n_5356;
wire n_6721;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_770;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_7008;
wire n_711;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_6111;
wire n_1834;
wire n_7505;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_6260;
wire n_7501;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_6665;
wire n_7566;
wire n_7055;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_5858;
wire n_5817;
wire n_6690;
wire n_3402;
wire n_5723;
wire n_5295;
wire n_6137;
wire n_4679;
wire n_4115;
wire n_6201;
wire n_726;
wire n_7113;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_818;
wire n_1970;
wire n_2766;
wire n_5627;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_7242;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_6461;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_6212;
wire n_3401;
wire n_6908;
wire n_3226;
wire n_6570;
wire n_1410;
wire n_707;
wire n_6498;
wire n_3902;
wire n_4730;
wire n_7228;
wire n_6692;
wire n_937;
wire n_6074;
wire n_2779;
wire n_7561;
wire n_1584;
wire n_6380;
wire n_3654;
wire n_2164;
wire n_5996;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_6045;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_6505;
wire n_2811;
wire n_3348;
wire n_7415;
wire n_5796;
wire n_7598;
wire n_6320;
wire n_6489;
wire n_6068;
wire n_895;
wire n_3358;
wire n_5791;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_6772;
wire n_1543;
wire n_1991;
wire n_2224;
wire n_6823;
wire n_6877;
wire n_732;
wire n_6806;
wire n_7426;
wire n_5906;
wire n_4743;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_6831;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_7217;
wire n_2692;
wire n_2008;
wire n_6284;
wire n_7058;
wire n_4654;
wire n_6157;
wire n_5423;
wire n_7497;
wire n_799;
wire n_6785;
wire n_1213;
wire n_6374;
wire n_6930;
wire n_4733;
wire n_3792;
wire n_6017;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_6838;
wire n_869;
wire n_5736;
wire n_6937;
wire n_6443;
wire n_3312;
wire n_6105;
wire n_1352;
wire n_2197;
wire n_7558;
wire n_2199;
wire n_5069;
wire n_7442;
wire n_5700;
wire n_6543;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_6091;
wire n_684;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_6674;
wire n_664;
wire n_2480;
wire n_6034;
wire n_7499;
wire n_2363;
wire n_4072;
wire n_916;
wire n_5579;
wire n_1115;
wire n_7085;
wire n_4781;
wire n_3606;
wire n_6652;
wire n_7098;
wire n_5004;
wire n_2550;
wire n_6762;
wire n_7341;
wire n_4424;
wire n_823;
wire n_725;
wire n_7611;
wire n_7391;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_5837;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_6895;
wire n_3878;
wire n_7646;
wire n_4450;
wire n_5642;
wire n_3553;
wire n_7224;
wire n_719;
wire n_5880;
wire n_6169;
wire n_4746;
wire n_7524;
wire n_5713;
wire n_6005;
wire n_1683;
wire n_1530;
wire n_997;
wire n_7627;
wire n_932;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_2996;
wire n_1268;
wire n_5793;
wire n_5591;
wire n_1320;
wire n_4050;
wire n_7496;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_5623;
wire n_1063;
wire n_5681;
wire n_4853;
wire n_981;
wire n_7399;
wire n_867;
wire n_2422;
wire n_6213;
wire n_2239;
wire n_6118;
wire n_5256;
wire n_2950;
wire n_7605;
wire n_5220;
wire n_5732;
wire n_3852;
wire n_5178;
wire n_812;
wire n_4520;
wire n_6814;
wire n_7342;
wire n_2057;
wire n_4008;
wire n_5507;
wire n_905;
wire n_7214;
wire n_7472;
wire n_5077;
wire n_782;
wire n_5872;
wire n_3858;
wire n_7408;
wire n_1901;
wire n_6115;
wire n_4502;
wire n_6858;
wire n_3032;
wire n_4851;
wire n_5735;
wire n_1330;
wire n_7254;
wire n_6944;
wire n_7384;
wire n_3072;
wire n_3313;
wire n_3081;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_769;
wire n_4571;
wire n_2006;
wire n_6430;
wire n_6193;
wire n_934;
wire n_5314;
wire n_6462;
wire n_1618;
wire n_826;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_6757;
wire n_6822;
wire n_2535;
wire n_4205;
wire n_5953;
wire n_2726;
wire n_7599;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_6779;
wire n_6518;
wire n_6797;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_1083;
wire n_5952;
wire n_4739;
wire n_5820;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_5718;
wire n_787;
wire n_6916;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_930;
wire n_3926;
wire n_6152;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_5777;
wire n_2764;
wire n_1498;
wire n_7046;
wire n_4225;
wire n_682;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_5926;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_6589;
wire n_7579;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_7173;
wire n_5951;
wire n_7092;
wire n_2442;
wire n_6197;
wire n_6971;
wire n_928;
wire n_1943;
wire n_7460;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_6154;
wire n_7344;
wire n_1396;
wire n_1348;
wire n_6020;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_5701;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_7079;
wire n_5120;
wire n_5470;
wire n_4565;
wire n_7675;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_5797;
wire n_6696;
wire n_4839;
wire n_5222;
wire n_5743;
wire n_1028;
wire n_4016;
wire n_6210;
wire n_5772;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_6964;
wire n_5801;
wire n_6117;
wire n_4231;
wire n_6202;
wire n_7279;
wire n_3165;
wire n_7670;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_6681;
wire n_5971;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_745;
wire n_2381;
wire n_6661;
wire n_3303;
wire n_1654;
wire n_6640;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_7371;
wire n_6962;
wire n_4101;
wire n_6455;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_7606;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_6963;
wire n_6644;
wire n_4389;
wire n_6896;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_6832;
wire n_1595;
wire n_2161;
wire n_6160;
wire n_7564;
wire n_2404;
wire n_2083;
wire n_6718;
wire n_2503;
wire n_6542;
wire n_1540;
wire n_1936;
wire n_6031;
wire n_5502;
wire n_2027;
wire n_5568;
wire n_2642;
wire n_720;
wire n_2500;
wire n_7653;
wire n_1918;
wire n_5656;
wire n_863;
wire n_6763;
wire n_4831;
wire n_2513;
wire n_5974;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_6280;
wire n_2414;
wire n_6438;
wire n_1402;
wire n_3662;
wire n_6316;
wire n_7383;
wire n_4319;
wire n_5474;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_5413;
wire n_6758;
wire n_2004;
wire n_5412;
wire n_3694;
wire n_2586;
wire n_6069;
wire n_5752;
wire n_6874;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_811;
wire n_6030;
wire n_6077;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_6299;
wire n_4474;
wire n_1089;
wire n_6386;
wire n_5217;
wire n_1004;
wire n_5957;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_7655;
wire n_5490;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_6708;
wire n_7433;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_7347;
wire n_4580;
wire n_6792;
wire n_7633;
wire n_1263;
wire n_6177;
wire n_5912;
wire n_1126;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_6033;
wire n_1859;
wire n_1677;
wire n_5557;
wire n_7397;
wire n_7389;
wire n_5472;
wire n_7602;
wire n_2955;
wire n_4112;
wire n_6002;
wire n_4337;
wire n_5711;
wire n_4138;
wire n_7554;
wire n_5396;
wire n_7693;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_1198;
wire n_6557;
wire n_7300;
wire n_956;
wire n_2134;
wire n_5960;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_7532;
wire n_5143;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_6142;
wire n_6917;
wire n_7510;
wire n_1545;
wire n_2374;
wire n_5859;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_854;
wire n_2396;
wire n_1799;
wire n_4734;
wire n_674;
wire n_1939;
wire n_2486;
wire n_6163;
wire n_4635;
wire n_3501;
wire n_1152;
wire n_7118;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_6285;
wire n_6778;
wire n_6025;
wire n_7257;
wire n_4242;
wire n_6862;
wire n_6319;
wire n_7067;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_7669;
wire n_5268;
wire n_6318;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_6089;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_1261;
wire n_6315;
wire n_938;
wire n_3186;
wire n_4955;
wire n_1154;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_5840;
wire n_2761;
wire n_6343;
wire n_3157;
wire n_709;
wire n_2537;
wire n_2144;
wire n_6049;
wire n_6919;
wire n_7423;
wire n_920;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_6052;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_7069;
wire n_6886;
wire n_1949;
wire n_976;
wire n_1946;
wire n_2936;
wire n_6912;
wire n_5914;
wire n_775;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_6061;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_7252;
wire n_5542;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_7133;
wire n_1850;
wire n_6883;
wire n_5519;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_6009;
wire n_7061;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_7518;
wire n_5586;
wire n_2693;
wire n_4065;
wire n_3798;
wire n_6378;
wire n_5187;
wire n_4944;
wire n_5675;
wire n_926;
wire n_2249;
wire n_2180;
wire n_4135;
wire n_1218;
wire n_2632;
wire n_6601;
wire n_5771;
wire n_7216;
wire n_1547;
wire n_777;
wire n_6407;
wire n_1755;
wire n_6749;
wire n_6839;
wire n_958;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_6051;
wire n_4716;
wire n_4942;
wire n_6217;
wire n_6680;
wire n_5844;
wire n_2432;
wire n_1521;
wire n_6532;
wire n_3405;
wire n_4745;
wire n_6155;
wire n_6446;
wire n_6738;
wire n_6250;
wire n_7458;
wire n_7614;
wire n_2337;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_6736;
wire n_5344;
wire n_923;
wire n_6526;
wire n_4629;
wire n_6339;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_6350;
wire n_7013;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_5662;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_5705;
wire n_4753;
wire n_4552;
wire n_7656;
wire n_3885;
wire n_6845;
wire n_7105;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_1197;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_6829;
wire n_5574;
wire n_5126;
wire n_1039;
wire n_6508;
wire n_2214;
wire n_2055;
wire n_3427;
wire n_4067;
wire n_1403;
wire n_5553;
wire n_4176;
wire n_4042;
wire n_7570;
wire n_4385;
wire n_3320;
wire n_7052;
wire n_5009;
wire n_7262;
wire n_5368;
wire n_2688;
wire n_1202;
wire n_5626;
wire n_6603;
wire n_6114;
wire n_1463;
wire n_6576;
wire n_3651;
wire n_4333;
wire n_7364;
wire n_3359;
wire n_7208;
wire n_6245;
wire n_2865;
wire n_2706;
wire n_5499;
wire n_6703;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_7202;
wire n_4246;
wire n_3580;
wire n_7011;
wire n_2139;
wire n_4609;
wire n_7621;
wire n_5291;
wire n_5876;
wire n_6970;
wire n_5114;
wire n_2674;
wire n_6409;
wire n_6704;
wire n_1565;
wire n_4088;
wire n_6876;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_7028;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_7313;
wire n_6255;
wire n_7320;
wire n_7343;
wire n_1072;
wire n_5288;
wire n_2305;
wire n_5540;
wire n_5699;
wire n_7525;
wire n_2450;
wire n_3447;
wire n_5810;
wire n_3305;
wire n_4148;
wire n_4151;
wire n_1712;
wire n_3528;
wire n_6938;
wire n_4373;
wire n_5762;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_7337;
wire n_6989;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_6427;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_7038;
wire n_4683;
wire n_5366;
wire n_728;
wire n_1162;
wire n_1847;
wire n_2767;
wire n_6360;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_6146;
wire n_887;
wire n_6270;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_5451;
wire n_3923;
wire n_931;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_5901;
wire n_6353;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_3643;
wire n_2825;
wire n_4876;
wire n_6345;
wire n_1997;
wire n_6691;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_7392;
wire n_2215;
wire n_5053;
wire n_1259;
wire n_6239;
wire n_4553;
wire n_706;
wire n_746;
wire n_6803;
wire n_784;
wire n_3978;
wire n_6340;
wire n_7583;
wire n_4809;
wire n_5226;
wire n_1244;
wire n_7657;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_5867;
wire n_6048;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_5590;
wire n_913;
wire n_6773;
wire n_3833;
wire n_5632;
wire n_865;
wire n_697;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_2022;
wire n_6336;
wire n_3814;
wire n_7041;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4911;
wire n_4842;
wire n_4340;
wire n_7370;
wire n_3513;
wire n_3133;
wire n_5660;
wire n_4645;
wire n_1191;
wire n_7557;
wire n_2992;
wire n_6174;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_6023;
wire n_2517;
wire n_6776;
wire n_3128;
wire n_5426;
wire n_6463;
wire n_744;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_6372;
wire n_7176;
wire n_1529;
wire n_2469;
wire n_5778;
wire n_5625;
wire n_6396;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_6669;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_5531;
wire n_3000;
wire n_5429;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1839;
wire n_1837;
wire n_5818;
wire n_5646;
wire n_6940;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_6394;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_7590;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_6995;
wire n_7185;
wire n_1656;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_6254;
wire n_6161;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_7332;
wire n_6660;
wire n_4771;
wire n_5719;
wire n_7225;
wire n_908;
wire n_6128;
wire n_4086;
wire n_2412;
wire n_7037;
wire n_4814;
wire n_724;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_5749;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_7409;
wire n_4692;
wire n_959;
wire n_3031;
wire n_7258;
wire n_7432;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_6334;
wire n_1169;
wire n_2666;
wire n_3385;
wire n_6848;
wire n_2171;
wire n_4708;
wire n_6321;
wire n_2768;
wire n_2314;
wire n_6794;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_1079;
wire n_7197;
wire n_5489;
wire n_1593;
wire n_6400;
wire n_3767;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_6705;
wire n_2162;
wire n_7619;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_750;
wire n_742;
wire n_5436;
wire n_5907;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_6044;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_6495;
wire n_5013;
wire n_2312;
wire n_7403;
wire n_6902;
wire n_6470;
wire n_3015;
wire n_1171;
wire n_1920;
wire n_1065;
wire n_5569;
wire n_5439;
wire n_5619;
wire n_4147;
wire n_2048;
wire n_6481;
wire n_3607;
wire n_4925;
wire n_7548;
wire n_1921;
wire n_1309;
wire n_6534;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_6181;
wire n_3276;
wire n_1177;
wire n_6728;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_5715;
wire n_6133;
wire n_6528;
wire n_7604;
wire n_7407;
wire n_1119;
wire n_1240;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_6670;
wire n_6774;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_6741;
wire n_7424;
wire n_700;
wire n_6038;
wire n_4818;
wire n_4514;
wire n_4800;
wire n_1366;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_6282;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_6700;
wire n_7334;
wire n_1591;
wire n_2033;
wire n_7684;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_5932;
wire n_6178;
wire n_1111;
wire n_2132;
wire n_6234;
wire n_6012;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_1140;
wire n_891;
wire n_3387;
wire n_5186;
wire n_7367;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_6715;
wire n_5828;
wire n_2831;
wire n_7200;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_7582;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_987;
wire n_3037;
wire n_6337;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_6770;
wire n_6743;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_1131;
wire n_6682;
wire n_5054;
wire n_7673;
wire n_5631;
wire n_2467;
wire n_6539;
wire n_1094;
wire n_7243;
wire n_7179;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_6314;
wire n_6617;
wire n_1209;
wire n_3592;
wire n_5694;
wire n_4650;
wire n_4888;
wire n_7274;
wire n_5326;
wire n_1435;
wire n_879;
wire n_3394;
wire n_4874;
wire n_7608;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_6595;
wire n_1645;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_4060;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_6385;
wire n_6289;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_7373;
wire n_3589;
wire n_952;
wire n_2534;
wire n_1229;
wire n_6186;
wire n_4799;
wire n_5153;
wire n_6257;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_6852;
wire n_2789;
wire n_6346;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_5809;
wire n_1897;
wire n_764;
wire n_1424;
wire n_5365;
wire n_2933;
wire n_7587;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_6274;
wire n_7372;
wire n_2328;
wire n_4248;
wire n_5915;
wire n_6818;
wire n_5452;
wire n_7226;
wire n_4754;
wire n_7057;
wire n_7685;
wire n_4554;
wire n_5595;
wire n_6609;
wire n_4845;
wire n_6753;
wire n_6815;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_6764;
wire n_5535;
wire n_1432;
wire n_3875;
wire n_5370;
wire n_6391;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_5594;
wire n_4301;
wire n_841;
wire n_4586;
wire n_1050;
wire n_1954;
wire n_4048;
wire n_6471;
wire n_1844;
wire n_3777;
wire n_6627;
wire n_5761;
wire n_4784;
wire n_7203;
wire n_2999;
wire n_7512;
wire n_1644;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_7215;
wire n_3080;
wire n_6636;
wire n_4199;
wire n_2701;
wire n_5929;
wire n_3362;
wire n_1631;
wire n_5559;
wire n_3105;
wire n_5478;
wire n_7388;
wire n_7694;
wire n_1179;
wire n_6243;
wire n_753;
wire n_6488;
wire n_1048;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_6022;
wire n_6457;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_692;
wire n_820;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_6867;
wire n_3417;
wire n_1143;
wire n_1579;
wire n_5868;
wire n_6230;
wire n_4034;
wire n_6538;
wire n_1688;
wire n_6633;
wire n_6187;
wire n_3327;
wire n_6172;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_7311;
wire n_2755;
wire n_5989;
wire n_3237;
wire n_6574;
wire n_1992;
wire n_6395;
wire n_4402;
wire n_4239;
wire n_6854;
wire n_3400;
wire n_6233;
wire n_4550;
wire n_6456;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_3382;
wire n_7488;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_7198;
wire n_1557;
wire n_4201;
wire n_6784;
wire n_6168;
wire n_896;
wire n_3316;
wire n_6766;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_6330;
wire n_2192;
wire n_5520;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_7249;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_5947;
wire n_7336;
wire n_4416;
wire n_3372;
wire n_7031;
wire n_4539;
wire n_814;
wire n_2707;
wire n_6799;
wire n_5920;
wire n_6672;
wire n_2471;
wire n_1472;
wire n_6149;
wire n_1671;
wire n_7142;
wire n_3230;
wire n_5808;
wire n_3342;
wire n_1062;
wire n_6054;
wire n_7089;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_1204;
wire n_6450;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_7042;
wire n_3780;
wire n_783;
wire n_1928;
wire n_5244;
wire n_6523;
wire n_5382;
wire n_1188;
wire n_6107;
wire n_3957;
wire n_6775;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_6232;
wire n_6445;
wire n_7181;
wire n_6134;
wire n_5384;
wire n_3608;
wire n_6056;
wire n_6932;
wire n_7036;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_5587;
wire n_2619;
wire n_6855;
wire n_2444;
wire n_5789;
wire n_1110;
wire n_3123;
wire n_5787;
wire n_6585;
wire n_6369;
wire n_5056;
wire n_1088;
wire n_5249;
wire n_3393;
wire n_7447;
wire n_866;
wire n_5198;
wire n_5360;
wire n_7455;
wire n_5233;
wire n_4887;
wire n_5829;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_6252;
wire n_5866;
wire n_6493;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_5899;
wire n_7629;
wire n_693;
wire n_4792;
wire n_7104;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_7601;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_6026;
wire n_4290;
wire n_5247;
wire n_5865;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_6544;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_7138;
wire n_7290;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_6679;
wire n_1371;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_5924;
wire n_3182;
wire n_7625;
wire n_5822;
wire n_2564;
wire n_6259;
wire n_4947;
wire n_876;
wire n_7284;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_3958;
wire n_6390;
wire n_3450;
wire n_966;
wire n_4729;
wire n_5786;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_3174;
wire n_982;
wire n_1453;
wire n_2217;
wire n_6630;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_5658;
wire n_3408;
wire n_899;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_6279;
wire n_1514;
wire n_1771;
wire n_1005;
wire n_679;
wire n_710;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_1168;
wire n_6813;
wire n_5564;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_7106;
wire n_6042;
wire n_7644;
wire n_1853;
wire n_1356;
wire n_6057;
wire n_1787;
wire n_4137;
wire n_7529;
wire n_6675;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_6476;
wire n_3972;
wire n_6207;
wire n_5539;
wire n_6268;
wire n_6878;
wire n_6286;
wire n_3308;
wire n_6524;
wire n_791;
wire n_1533;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_6225;
wire n_4322;
wire n_1720;
wire n_7297;
wire n_6291;
wire n_2830;
wire n_5893;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_7199;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_715;
wire n_1480;
wire n_5261;
wire n_6520;
wire n_7648;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_1782;
wire n_2245;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_810;
wire n_2965;
wire n_3635;
wire n_6024;
wire n_5022;
wire n_5005;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_7487;
wire n_2213;
wire n_1170;
wire n_6425;
wire n_5993;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_7638;
wire n_5703;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_855;
wire n_5534;
wire n_6432;
wire n_1461;
wire n_3204;
wire n_7259;
wire n_2136;
wire n_6540;
wire n_6955;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_698;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_7237;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_6388;
wire n_5904;
wire n_4880;
wire n_6760;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_5572;
wire n_5750;
wire n_7063;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_7576;
wire n_1762;
wire n_1013;
wire n_718;
wire n_3023;
wire n_6795;
wire n_5881;
wire n_6664;
wire n_5815;
wire n_6261;
wire n_4193;
wire n_5873;
wire n_4075;
wire n_3104;
wire n_6487;
wire n_4737;
wire n_6729;
wire n_3647;
wire n_5755;
wire n_825;
wire n_2819;
wire n_5949;
wire n_737;
wire n_5195;
wire n_7483;
wire n_3609;
wire n_4136;
wire n_6608;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_7385;
wire n_3720;
wire n_4535;
wire n_7668;
wire n_733;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_6663;
wire n_4794;
wire n_5955;
wire n_7476;
wire n_3959;
wire n_7327;
wire n_5763;
wire n_6656;
wire n_792;
wire n_6843;
wire n_3140;
wire n_5246;
wire n_5964;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_7266;
wire n_5164;
wire n_4196;
wire n_6969;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_5665;
wire n_6485;
wire n_3069;
wire n_5498;
wire n_7100;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5783;
wire n_5183;
wire n_6075;
wire n_7082;
wire n_3084;
wire n_6120;
wire n_1727;
wire n_6659;
wire n_2735;
wire n_6750;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_1046;
wire n_3761;
wire n_7689;
wire n_4889;
wire n_7132;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_5739;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_6003;
wire n_5385;
wire n_4558;
wire n_6478;
wire n_2172;
wire n_6066;
wire n_7034;
wire n_6086;
wire n_4722;
wire n_6650;
wire n_6224;
wire n_1129;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_961;
wire n_2250;
wire n_7084;
wire n_5845;
wire n_7293;
wire n_1225;
wire n_4092;
wire n_5990;
wire n_3908;
wire n_6175;
wire n_6060;
wire n_7253;
wire n_2423;
wire n_3671;
wire n_6891;
wire n_5663;
wire n_994;
wire n_6410;
wire n_3344;
wire n_2194;
wire n_848;
wire n_4465;
wire n_5973;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_1223;
wire n_2680;
wire n_6059;
wire n_5130;
wire n_1567;
wire n_7520;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_6103;
wire n_6809;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_6267;
wire n_1797;
wire n_2957;
wire n_5855;
wire n_2357;
wire n_1250;
wire n_5757;
wire n_6437;
wire n_3309;
wire n_7331;
wire n_6610;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_6957;
wire n_5704;
wire n_7514;
wire n_7163;
wire n_7620;
wire n_2570;
wire n_1086;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_5473;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_5946;
wire n_2744;
wire n_6711;
wire n_4287;
wire n_2397;
wire n_7445;
wire n_2208;
wire n_6847;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_7123;
wire n_6384;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_1113;
wire n_7563;
wire n_6298;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_7361;
wire n_852;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_7322;
wire n_5710;
wire n_7453;
wire n_6067;
wire n_5070;
wire n_6377;
wire n_1337;
wire n_4445;
wire n_699;
wire n_5566;
wire n_5414;
wire n_1627;
wire n_1245;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_6348;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_6129;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_6834;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_6136;
wire n_7261;
wire n_6723;
wire n_5834;
wire n_2823;
wire n_1076;
wire n_1408;
wire n_1761;
wire n_5874;
wire n_730;
wire n_7508;
wire n_7021;
wire n_5270;
wire n_5956;
wire n_795;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_6078;
wire n_7000;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_7130;
wire n_1526;
wire n_5823;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_5465;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_7538;
wire n_712;
wire n_7517;
wire n_1583;
wire n_5853;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_7077;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_6642;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_7346;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_7333;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_7546;
wire n_3853;
wire n_4216;
wire n_5934;
wire n_6942;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_6511;
wire n_3721;
wire n_1254;
wire n_6507;
wire n_1026;
wire n_2026;
wire n_1234;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_1032;
wire n_2614;
wire n_7319;
wire n_2991;
wire n_6497;
wire n_6001;
wire n_6007;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_6606;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_5395;
wire n_2237;
wire n_7078;
wire n_3463;
wire n_7047;
wire n_3699;
wire n_5067;
wire n_7107;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_7469;
wire n_2728;
wire n_3857;

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_578),
.Y(n_661)
);

BUFx2_ASAP7_75t_SL g662 ( 
.A(n_651),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_138),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_48),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_441),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_383),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_477),
.Y(n_667)
);

CKINVDCx16_ASAP7_75t_R g668 ( 
.A(n_411),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_104),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_417),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_384),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_604),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_498),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_371),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_179),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_14),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_47),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_334),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_294),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_519),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_514),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_409),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_287),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_347),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_223),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_173),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_262),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_167),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_475),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_506),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_203),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_620),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_475),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_137),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_189),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_292),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_605),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_187),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_561),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_304),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_353),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_143),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_84),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_9),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_653),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_140),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_299),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_557),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_641),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_186),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_489),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_429),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_103),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_291),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_119),
.Y(n_715)
);

BUFx8_ASAP7_75t_SL g716 ( 
.A(n_360),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_546),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_507),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_655),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_320),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_385),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_264),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_436),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_170),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_85),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_142),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_44),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_78),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_411),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_209),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_291),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_650),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_591),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_490),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_304),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_474),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_358),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_279),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_631),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_351),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_8),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_520),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_31),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_272),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_149),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_229),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_24),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_147),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_292),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_649),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_494),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_133),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_233),
.Y(n_753)
);

CKINVDCx14_ASAP7_75t_R g754 ( 
.A(n_272),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_319),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_332),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_182),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_434),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_469),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_218),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_247),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_41),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_303),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_12),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_234),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_177),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_556),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_155),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_163),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_148),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_517),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_34),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_616),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_562),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_652),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_615),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_581),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_442),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_367),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_579),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_146),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_567),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_316),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_322),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_554),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_466),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_499),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_201),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_22),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_499),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_244),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_215),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_481),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_109),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_103),
.Y(n_795)
);

HB1xp67_ASAP7_75t_SL g796 ( 
.A(n_476),
.Y(n_796)
);

CKINVDCx14_ASAP7_75t_R g797 ( 
.A(n_403),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_1),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_504),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_494),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_596),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_370),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_441),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_522),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_332),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_548),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_242),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_275),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_24),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_301),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_307),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_456),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_552),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_416),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_342),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_1),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_49),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_56),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_223),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_496),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_534),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_151),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_585),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_581),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_454),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_53),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_23),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_65),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_370),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_422),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_287),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_249),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_34),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_514),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_60),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_306),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_359),
.Y(n_837)
);

BUFx10_ASAP7_75t_L g838 ( 
.A(n_328),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_542),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_310),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_439),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_55),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_574),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_140),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_112),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_180),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_549),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_23),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_183),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_216),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_74),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_242),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_13),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_305),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_70),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_342),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_225),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_98),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_423),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_595),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_48),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_561),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_607),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_247),
.Y(n_864)
);

BUFx2_ASAP7_75t_SL g865 ( 
.A(n_124),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_516),
.Y(n_866)
);

BUFx10_ASAP7_75t_L g867 ( 
.A(n_483),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_421),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_617),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_76),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_446),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_451),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_204),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_194),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_205),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_69),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_30),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_390),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_637),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_176),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_439),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_115),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_42),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_11),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_393),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_357),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_602),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_485),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_314),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_572),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_53),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_63),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_288),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_599),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_180),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_469),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_398),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_603),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_461),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_52),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_323),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_183),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_177),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_402),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_536),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_171),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_275),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_158),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_270),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_471),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_125),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_457),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_124),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_550),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_109),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_630),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_393),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_259),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_225),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_535),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_464),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_251),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_445),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_306),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_529),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_407),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_286),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_17),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_557),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_546),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_436),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_403),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_584),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_625),
.Y(n_934)
);

CKINVDCx16_ASAP7_75t_R g935 ( 
.A(n_4),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_47),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_406),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_52),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_606),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_659),
.Y(n_940)
);

BUFx10_ASAP7_75t_L g941 ( 
.A(n_563),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_260),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_3),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_372),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_354),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_467),
.Y(n_946)
);

INVx4_ASAP7_75t_R g947 ( 
.A(n_285),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_645),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_81),
.Y(n_949)
);

CKINVDCx16_ASAP7_75t_R g950 ( 
.A(n_483),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_383),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_3),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_614),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_288),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_160),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_123),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_299),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_432),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_580),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_620),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_613),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_18),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_168),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_627),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_333),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_5),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_642),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_450),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_432),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_639),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_386),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_497),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_380),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_131),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_252),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_255),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_419),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_365),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_482),
.Y(n_979)
);

BUFx10_ASAP7_75t_L g980 ( 
.A(n_385),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_491),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_132),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_321),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_43),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_612),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_523),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_45),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_294),
.Y(n_988)
);

BUFx10_ASAP7_75t_L g989 ( 
.A(n_646),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_331),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_417),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_551),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_10),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_326),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_262),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_75),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_100),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_496),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_228),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_93),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_538),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_171),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_76),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_446),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_307),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_567),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_531),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_597),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_633),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_283),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_67),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_584),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_596),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_372),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_338),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_90),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_464),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_209),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_45),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_25),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_202),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_350),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_365),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_602),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_643),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_107),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_224),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_337),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_229),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_228),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_440),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_465),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_82),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_654),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_333),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_130),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_248),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_219),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_520),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_321),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_324),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_476),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_542),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_606),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_462),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_90),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_558),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_656),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_349),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_481),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_495),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_71),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_310),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_320),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_472),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_7),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_623),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_613),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_256),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_472),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_205),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_16),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_463),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_338),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_564),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_318),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_219),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_57),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_80),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_153),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_309),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_159),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_407),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_164),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_580),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_134),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_528),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_64),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_67),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_85),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_311),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_166),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_590),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_258),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_334),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_145),
.Y(n_1086)
);

CKINVDCx16_ASAP7_75t_R g1087 ( 
.A(n_208),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_516),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_35),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_200),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_239),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_492),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_612),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_538),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_357),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_248),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_421),
.Y(n_1097)
);

BUFx8_ASAP7_75t_SL g1098 ( 
.A(n_438),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_271),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_218),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_15),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_298),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_363),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_46),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_367),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_179),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_638),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_644),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_96),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_250),
.Y(n_1110)
);

BUFx10_ASAP7_75t_L g1111 ( 
.A(n_323),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_215),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_513),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_312),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_284),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_341),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_398),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_54),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_111),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_536),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_583),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_208),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_227),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_470),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_594),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_547),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_470),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_597),
.Y(n_1128)
);

CKINVDCx16_ASAP7_75t_R g1129 ( 
.A(n_232),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_195),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_412),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_13),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_473),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_493),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_386),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_455),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_444),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_381),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_463),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_628),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_255),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_592),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_96),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_505),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_100),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_577),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_376),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_78),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_61),
.Y(n_1149)
);

CKINVDCx14_ASAP7_75t_R g1150 ( 
.A(n_243),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_394),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_251),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_296),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_9),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_373),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_107),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_465),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_426),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_16),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_231),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_122),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_344),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_622),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_197),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_176),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_2),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_541),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_5),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_135),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_314),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_491),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_316),
.Y(n_1172)
);

CKINVDCx16_ASAP7_75t_R g1173 ( 
.A(n_268),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_640),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_589),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_414),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_174),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_252),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_6),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_198),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_374),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_619),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_20),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_489),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_647),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_519),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_113),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_413),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_387),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_501),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_347),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_261),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_409),
.Y(n_1193)
);

BUFx10_ASAP7_75t_L g1194 ( 
.A(n_119),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_582),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_276),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_426),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_543),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_371),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_468),
.Y(n_1200)
);

BUFx2_ASAP7_75t_SL g1201 ( 
.A(n_74),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_530),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_562),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_624),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_305),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_648),
.Y(n_1206)
);

CKINVDCx16_ASAP7_75t_R g1207 ( 
.A(n_268),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_591),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_19),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_705),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_716),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_716),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_739),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_739),
.Y(n_1214)
);

CKINVDCx14_ASAP7_75t_R g1215 ( 
.A(n_754),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_989),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_989),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_750),
.Y(n_1218)
);

CKINVDCx14_ASAP7_75t_R g1219 ( 
.A(n_754),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_750),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1098),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_775),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1098),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_775),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_797),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_797),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_916),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1150),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_989),
.Y(n_1229)
);

NOR2xp67_ASAP7_75t_L g1230 ( 
.A(n_1183),
.B(n_0),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_734),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1150),
.Y(n_1232)
);

INVxp67_ASAP7_75t_L g1233 ( 
.A(n_734),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1183),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_916),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_948),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_948),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1207),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1207),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_668),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_668),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1174),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_703),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1174),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_989),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_663),
.B(n_664),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_682),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_682),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_705),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_970),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1183),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_764),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_719),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_682),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_764),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_935),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1183),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_686),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_686),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_763),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_686),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_935),
.Y(n_1262)
);

BUFx10_ASAP7_75t_L g1263 ( 
.A(n_990),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_950),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_757),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_757),
.Y(n_1266)
);

BUFx10_ASAP7_75t_L g1267 ( 
.A(n_990),
.Y(n_1267)
);

BUFx10_ASAP7_75t_L g1268 ( 
.A(n_1028),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_757),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_831),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_703),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_950),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1028),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_831),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1087),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_831),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1087),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_663),
.B(n_0),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1129),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_843),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_843),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1129),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_843),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_856),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_856),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_856),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_732),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1173),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_879),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_860),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_940),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_740),
.Y(n_1292)
);

CKINVDCx16_ASAP7_75t_R g1293 ( 
.A(n_1173),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_666),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1187),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_667),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_669),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_763),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_967),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_763),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1009),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_763),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_860),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1034),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_860),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_874),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_672),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_740),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1048),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_820),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_874),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_679),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1107),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_684),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_874),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_689),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_945),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_945),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_690),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_945),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1108),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1046),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1046),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_691),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_970),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_664),
.B(n_2),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1046),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_763),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_695),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_763),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_796),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1065),
.Y(n_1332)
);

INVxp33_ASAP7_75t_L g1333 ( 
.A(n_1187),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_696),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1065),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1065),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_970),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_697),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_820),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_701),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_970),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_702),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1067),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1067),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_704),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1067),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_706),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_960),
.Y(n_1348)
);

CKINVDCx16_ASAP7_75t_R g1349 ( 
.A(n_796),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_960),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1025),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1025),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1025),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_707),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_763),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_966),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_710),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_713),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_714),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_773),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_773),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_773),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_966),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_773),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_773),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_717),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_721),
.Y(n_1367)
);

BUFx10_ASAP7_75t_L g1368 ( 
.A(n_773),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1185),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_773),
.Y(n_1370)
);

INVxp67_ASAP7_75t_SL g1371 ( 
.A(n_850),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_722),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_712),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_723),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_725),
.Y(n_1375)
);

BUFx10_ASAP7_75t_L g1376 ( 
.A(n_850),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_850),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_726),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1082),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_850),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_850),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_728),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_727),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_712),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_850),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_850),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_918),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_735),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_918),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_918),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_736),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_918),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_1082),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_918),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_742),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_918),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_970),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_918),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_972),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_972),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_972),
.Y(n_1401)
);

CKINVDCx16_ASAP7_75t_R g1402 ( 
.A(n_712),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_972),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_972),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_972),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_743),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_746),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_972),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_996),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_748),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_996),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_996),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_996),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_749),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_751),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_970),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_996),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_752),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_756),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_996),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_758),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_970),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_759),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_996),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1075),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_760),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1075),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_761),
.Y(n_1428)
);

BUFx10_ASAP7_75t_L g1429 ( 
.A(n_1075),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1075),
.Y(n_1430)
);

CKINVDCx16_ASAP7_75t_R g1431 ( 
.A(n_712),
.Y(n_1431)
);

CKINVDCx16_ASAP7_75t_R g1432 ( 
.A(n_838),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1075),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1075),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1075),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_670),
.Y(n_1436)
);

BUFx5_ASAP7_75t_L g1437 ( 
.A(n_670),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_675),
.Y(n_1438)
);

BUFx2_ASAP7_75t_SL g1439 ( 
.A(n_709),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_762),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_838),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_730),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_765),
.Y(n_1443)
);

CKINVDCx14_ASAP7_75t_R g1444 ( 
.A(n_1139),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_770),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_772),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_774),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_709),
.B(n_1206),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_777),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_665),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_780),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_781),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_675),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1139),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_676),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_782),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_783),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_676),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1197),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_785),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_677),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_677),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_786),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_789),
.Y(n_1464)
);

CKINVDCx16_ASAP7_75t_R g1465 ( 
.A(n_838),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_678),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_678),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_680),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_680),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_681),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_791),
.Y(n_1471)
);

INVxp33_ASAP7_75t_L g1472 ( 
.A(n_1197),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_681),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_794),
.Y(n_1474)
);

CKINVDCx16_ASAP7_75t_R g1475 ( 
.A(n_838),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_687),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1203),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_687),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_692),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_692),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_693),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_795),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_799),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_802),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_867),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_867),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_693),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_694),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_694),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_803),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_805),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_699),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_806),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_699),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_807),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_809),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_700),
.Y(n_1497)
);

CKINVDCx16_ASAP7_75t_R g1498 ( 
.A(n_867),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_737),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_810),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_700),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_708),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_811),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_708),
.Y(n_1504)
);

BUFx10_ASAP7_75t_L g1505 ( 
.A(n_828),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_812),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_711),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1203),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_711),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_813),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_665),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_715),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_715),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_814),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_744),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_815),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_816),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_718),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_718),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_766),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_720),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_720),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_724),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_817),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_771),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_724),
.Y(n_1526)
);

CKINVDCx14_ASAP7_75t_R g1527 ( 
.A(n_867),
.Y(n_1527)
);

CKINVDCx16_ASAP7_75t_R g1528 ( 
.A(n_941),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_793),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_729),
.Y(n_1530)
);

BUFx2_ASAP7_75t_SL g1531 ( 
.A(n_1206),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_821),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_729),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_731),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_941),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_941),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_731),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_865),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_822),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_665),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_733),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_733),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_798),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_738),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_738),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_741),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_826),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_832),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_833),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_741),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_837),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_745),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_745),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_753),
.Y(n_1554)
);

NOR2xp67_ASAP7_75t_L g1555 ( 
.A(n_888),
.B(n_4),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_753),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_685),
.Y(n_1557)
);

CKINVDCx16_ASAP7_75t_R g1558 ( 
.A(n_941),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_839),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_767),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_840),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_842),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_685),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_847),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_767),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_852),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_854),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_685),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_769),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_855),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_824),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_836),
.Y(n_1572)
);

CKINVDCx20_ASAP7_75t_R g1573 ( 
.A(n_862),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_857),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_769),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_858),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_747),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_776),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_776),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_861),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_870),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_863),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_914),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_779),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_871),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_873),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_875),
.Y(n_1587)
);

CKINVDCx16_ASAP7_75t_R g1588 ( 
.A(n_980),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_956),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_779),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_784),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_980),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_784),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_878),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_880),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_882),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_787),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_883),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_747),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_787),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_790),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_980),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_885),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_889),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_747),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_890),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_790),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_891),
.Y(n_1608)
);

NOR2xp67_ASAP7_75t_L g1609 ( 
.A(n_888),
.B(n_6),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_792),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_792),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_800),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_800),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_892),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_895),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_896),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_980),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_897),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_801),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_768),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_901),
.Y(n_1621)
);

CKINVDCx16_ASAP7_75t_R g1622 ( 
.A(n_1111),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_801),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_902),
.Y(n_1624)
);

BUFx10_ASAP7_75t_L g1625 ( 
.A(n_828),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_804),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_971),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_904),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_804),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_1038),
.Y(n_1630)
);

CKINVDCx20_ASAP7_75t_R g1631 ( 
.A(n_1040),
.Y(n_1631)
);

NOR2xp67_ASAP7_75t_L g1632 ( 
.A(n_828),
.B(n_7),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_808),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_808),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_768),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1042),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_906),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_907),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_768),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_818),
.Y(n_1640)
);

BUFx10_ASAP7_75t_L g1641 ( 
.A(n_835),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_908),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_778),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_818),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1069),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_911),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_819),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_919),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_835),
.B(n_10),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_819),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_823),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_823),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_827),
.B(n_8),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_920),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_921),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_925),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_926),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1073),
.Y(n_1658)
);

CKINVDCx20_ASAP7_75t_R g1659 ( 
.A(n_1090),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_927),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_661),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_827),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_830),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_830),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_778),
.Y(n_1665)
);

CKINVDCx16_ASAP7_75t_R g1666 ( 
.A(n_1111),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_834),
.B(n_11),
.Y(n_1667)
);

CKINVDCx16_ASAP7_75t_R g1668 ( 
.A(n_1111),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_778),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_661),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_928),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_834),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_825),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_841),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_929),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_841),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_844),
.Y(n_1677)
);

BUFx5_ASAP7_75t_L g1678 ( 
.A(n_844),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_845),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_930),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_825),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_931),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_932),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_933),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_845),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_846),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_825),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_846),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_848),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_848),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_849),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_849),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_851),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_968),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1253),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1371),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_1210),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1234),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1287),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1234),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1251),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1289),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_1291),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1299),
.Y(n_1704)
);

CKINVDCx20_ASAP7_75t_R g1705 ( 
.A(n_1249),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1251),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1260),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1257),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1258),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1259),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1301),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1261),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1265),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1448),
.B(n_662),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1661),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_1670),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1383),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1304),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1266),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1309),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1269),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1439),
.B(n_662),
.Y(n_1722)
);

INVxp67_ASAP7_75t_SL g1723 ( 
.A(n_1538),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1270),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1274),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1313),
.Y(n_1726)
);

CKINVDCx20_ASAP7_75t_R g1727 ( 
.A(n_1442),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1280),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1281),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1283),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1284),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1285),
.Y(n_1732)
);

INVxp33_ASAP7_75t_SL g1733 ( 
.A(n_1225),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1286),
.Y(n_1734)
);

CKINVDCx20_ASAP7_75t_R g1735 ( 
.A(n_1499),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1290),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1303),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1305),
.Y(n_1738)
);

INVxp67_ASAP7_75t_SL g1739 ( 
.A(n_1248),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1306),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1311),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1315),
.Y(n_1742)
);

CKINVDCx16_ASAP7_75t_R g1743 ( 
.A(n_1331),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1248),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1531),
.B(n_835),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1317),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1318),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1321),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1320),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1322),
.Y(n_1750)
);

INVxp33_ASAP7_75t_SL g1751 ( 
.A(n_1225),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1594),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1323),
.Y(n_1753)
);

NOR2xp67_ASAP7_75t_L g1754 ( 
.A(n_1294),
.B(n_629),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1327),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1369),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1238),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1332),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1349),
.Y(n_1759)
);

CKINVDCx20_ASAP7_75t_R g1760 ( 
.A(n_1515),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1335),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1216),
.B(n_864),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1336),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1216),
.B(n_864),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1215),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1294),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1343),
.Y(n_1767)
);

INVxp67_ASAP7_75t_SL g1768 ( 
.A(n_1254),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1346),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1296),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1213),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1296),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1230),
.B(n_968),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1614),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1214),
.Y(n_1775)
);

CKINVDCx20_ASAP7_75t_R g1776 ( 
.A(n_1520),
.Y(n_1776)
);

CKINVDCx20_ASAP7_75t_R g1777 ( 
.A(n_1529),
.Y(n_1777)
);

INVxp67_ASAP7_75t_SL g1778 ( 
.A(n_1254),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1682),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1218),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1297),
.Y(n_1781)
);

CKINVDCx20_ASAP7_75t_R g1782 ( 
.A(n_1543),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1238),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1220),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1222),
.Y(n_1785)
);

INVxp67_ASAP7_75t_L g1786 ( 
.A(n_1566),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1297),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1307),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1224),
.Y(n_1789)
);

CKINVDCx16_ASAP7_75t_R g1790 ( 
.A(n_1293),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1307),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1226),
.B(n_864),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1227),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1235),
.Y(n_1794)
);

INVxp67_ASAP7_75t_SL g1795 ( 
.A(n_1276),
.Y(n_1795)
);

INVxp67_ASAP7_75t_SL g1796 ( 
.A(n_1276),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1312),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1236),
.Y(n_1798)
);

CKINVDCx20_ASAP7_75t_R g1799 ( 
.A(n_1572),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1237),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1242),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1244),
.Y(n_1802)
);

CKINVDCx16_ASAP7_75t_R g1803 ( 
.A(n_1527),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1246),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1226),
.B(n_1228),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1312),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1246),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1314),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1314),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1316),
.Y(n_1810)
);

CKINVDCx20_ASAP7_75t_R g1811 ( 
.A(n_1573),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1344),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1316),
.Y(n_1813)
);

CKINVDCx20_ASAP7_75t_R g1814 ( 
.A(n_1582),
.Y(n_1814)
);

CKINVDCx16_ASAP7_75t_R g1815 ( 
.A(n_1219),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1239),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1344),
.Y(n_1817)
);

CKINVDCx16_ASAP7_75t_R g1818 ( 
.A(n_1384),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1355),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_1319),
.Y(n_1820)
);

CKINVDCx20_ASAP7_75t_R g1821 ( 
.A(n_1583),
.Y(n_1821)
);

CKINVDCx20_ASAP7_75t_R g1822 ( 
.A(n_1589),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1576),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1319),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1360),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1324),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1228),
.B(n_877),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1324),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1329),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1450),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1329),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1361),
.Y(n_1832)
);

NOR2xp67_ASAP7_75t_L g1833 ( 
.A(n_1334),
.B(n_632),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1260),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1334),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1364),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1338),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1232),
.B(n_877),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1239),
.Y(n_1839)
);

NOR2xp67_ASAP7_75t_L g1840 ( 
.A(n_1338),
.B(n_634),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1232),
.B(n_877),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1377),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1380),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1340),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1381),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1340),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1342),
.Y(n_1847)
);

INVxp33_ASAP7_75t_SL g1848 ( 
.A(n_1211),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1385),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1387),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1587),
.Y(n_1851)
);

INVxp33_ASAP7_75t_SL g1852 ( 
.A(n_1211),
.Y(n_1852)
);

CKINVDCx20_ASAP7_75t_R g1853 ( 
.A(n_1627),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1240),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1390),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1342),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1240),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1298),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1345),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1345),
.Y(n_1860)
);

CKINVDCx20_ASAP7_75t_R g1861 ( 
.A(n_1630),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1392),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_1631),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1347),
.Y(n_1864)
);

INVx3_ASAP7_75t_L g1865 ( 
.A(n_1450),
.Y(n_1865)
);

INVxp67_ASAP7_75t_SL g1866 ( 
.A(n_1441),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1394),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1396),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1347),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1217),
.B(n_1001),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1298),
.Y(n_1871)
);

CKINVDCx20_ASAP7_75t_R g1872 ( 
.A(n_1659),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1398),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1354),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1354),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1357),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1399),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1401),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1403),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1300),
.Y(n_1880)
);

NOR2xp67_ASAP7_75t_L g1881 ( 
.A(n_1357),
.B(n_635),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1404),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1358),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1358),
.Y(n_1884)
);

CKINVDCx20_ASAP7_75t_R g1885 ( 
.A(n_1212),
.Y(n_1885)
);

CKINVDCx20_ASAP7_75t_R g1886 ( 
.A(n_1212),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1405),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_R g1888 ( 
.A(n_1359),
.B(n_1366),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1359),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_1366),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1408),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1221),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1409),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1367),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1587),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1367),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1372),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1372),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1411),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1412),
.Y(n_1900)
);

INVxp67_ASAP7_75t_L g1901 ( 
.A(n_1441),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1374),
.Y(n_1902)
);

INVxp67_ASAP7_75t_L g1903 ( 
.A(n_1485),
.Y(n_1903)
);

NAND2xp33_ASAP7_75t_R g1904 ( 
.A(n_1374),
.B(n_936),
.Y(n_1904)
);

BUFx3_ASAP7_75t_L g1905 ( 
.A(n_1247),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1485),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1375),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1413),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1417),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1420),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1424),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1425),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1427),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1430),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1300),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1375),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1433),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1525),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1217),
.B(n_1001),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1378),
.Y(n_1920)
);

CKINVDCx20_ASAP7_75t_R g1921 ( 
.A(n_1221),
.Y(n_1921)
);

INVxp67_ASAP7_75t_SL g1922 ( 
.A(n_1486),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1223),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1435),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1386),
.Y(n_1925)
);

CKINVDCx20_ASAP7_75t_R g1926 ( 
.A(n_1223),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1386),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1389),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1450),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_1378),
.Y(n_1930)
);

INVxp67_ASAP7_75t_SL g1931 ( 
.A(n_1486),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1389),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1382),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1400),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1382),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1388),
.Y(n_1936)
);

CKINVDCx20_ASAP7_75t_R g1937 ( 
.A(n_1444),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1302),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1388),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1391),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1400),
.Y(n_1941)
);

CKINVDCx20_ASAP7_75t_R g1942 ( 
.A(n_1402),
.Y(n_1942)
);

CKINVDCx20_ASAP7_75t_R g1943 ( 
.A(n_1431),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1436),
.Y(n_1944)
);

BUFx10_ASAP7_75t_L g1945 ( 
.A(n_1391),
.Y(n_1945)
);

INVxp67_ASAP7_75t_L g1946 ( 
.A(n_1536),
.Y(n_1946)
);

CKINVDCx20_ASAP7_75t_R g1947 ( 
.A(n_1432),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1395),
.Y(n_1948)
);

INVxp33_ASAP7_75t_L g1949 ( 
.A(n_1348),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1536),
.Y(n_1950)
);

INVx3_ASAP7_75t_L g1951 ( 
.A(n_1450),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1241),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1229),
.B(n_1001),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1395),
.Y(n_1954)
);

INVxp67_ASAP7_75t_L g1955 ( 
.A(n_1592),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1438),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1453),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1455),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1458),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1461),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1462),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1466),
.Y(n_1962)
);

BUFx10_ASAP7_75t_L g1963 ( 
.A(n_1406),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1467),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1468),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1469),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1406),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1470),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1407),
.Y(n_1969)
);

CKINVDCx20_ASAP7_75t_R g1970 ( 
.A(n_1465),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1241),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1407),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_R g1973 ( 
.A(n_1410),
.B(n_937),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1473),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1302),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1476),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1410),
.Y(n_1977)
);

CKINVDCx20_ASAP7_75t_R g1978 ( 
.A(n_1475),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1478),
.Y(n_1979)
);

INVxp67_ASAP7_75t_SL g1980 ( 
.A(n_1592),
.Y(n_1980)
);

CKINVDCx20_ASAP7_75t_R g1981 ( 
.A(n_1498),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1479),
.Y(n_1982)
);

CKINVDCx20_ASAP7_75t_R g1983 ( 
.A(n_1528),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1480),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1481),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1487),
.Y(n_1986)
);

XNOR2x1_ASAP7_75t_L g1987 ( 
.A(n_1571),
.B(n_671),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_1414),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1229),
.B(n_1037),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_1558),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1488),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1489),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1414),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1415),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1492),
.Y(n_1995)
);

BUFx2_ASAP7_75t_L g1996 ( 
.A(n_1252),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1415),
.Y(n_1997)
);

INVx1_ASAP7_75t_SL g1998 ( 
.A(n_1636),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1494),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1418),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1497),
.Y(n_2001)
);

CKINVDCx20_ASAP7_75t_R g2002 ( 
.A(n_1588),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1501),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1418),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1502),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_1419),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1504),
.Y(n_2007)
);

BUFx3_ASAP7_75t_L g2008 ( 
.A(n_1247),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1507),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1419),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1602),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1421),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1252),
.Y(n_2013)
);

CKINVDCx20_ASAP7_75t_R g2014 ( 
.A(n_1622),
.Y(n_2014)
);

CKINVDCx20_ASAP7_75t_R g2015 ( 
.A(n_1666),
.Y(n_2015)
);

CKINVDCx20_ASAP7_75t_R g2016 ( 
.A(n_1668),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1509),
.Y(n_2017)
);

CKINVDCx16_ASAP7_75t_R g2018 ( 
.A(n_1645),
.Y(n_2018)
);

INVxp67_ASAP7_75t_SL g2019 ( 
.A(n_1602),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1512),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1421),
.Y(n_2021)
);

CKINVDCx20_ASAP7_75t_R g2022 ( 
.A(n_1255),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1245),
.B(n_1037),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1513),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1518),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1519),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1521),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1522),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1523),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1526),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1423),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1530),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1423),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1533),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1534),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1537),
.Y(n_2036)
);

CKINVDCx20_ASAP7_75t_R g2037 ( 
.A(n_1255),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1245),
.B(n_1037),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1541),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1426),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1328),
.Y(n_2041)
);

NOR2xp67_ASAP7_75t_L g2042 ( 
.A(n_1426),
.B(n_636),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1542),
.Y(n_2043)
);

CKINVDCx20_ASAP7_75t_R g2044 ( 
.A(n_1256),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_1428),
.B(n_1052),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1428),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1440),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1440),
.B(n_1052),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1443),
.Y(n_2049)
);

CKINVDCx20_ASAP7_75t_R g2050 ( 
.A(n_1256),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1443),
.Y(n_2051)
);

CKINVDCx20_ASAP7_75t_R g2052 ( 
.A(n_1262),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1544),
.Y(n_2053)
);

CKINVDCx20_ASAP7_75t_R g2054 ( 
.A(n_1262),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1292),
.B(n_1198),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1545),
.Y(n_2056)
);

INVxp67_ASAP7_75t_SL g2057 ( 
.A(n_1617),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1546),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_1445),
.Y(n_2059)
);

INVxp67_ASAP7_75t_L g2060 ( 
.A(n_1617),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1550),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_1308),
.B(n_1339),
.Y(n_2062)
);

CKINVDCx20_ASAP7_75t_R g2063 ( 
.A(n_1264),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_1459),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1445),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1446),
.B(n_1052),
.Y(n_2066)
);

CKINVDCx20_ASAP7_75t_R g2067 ( 
.A(n_1264),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1446),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_1368),
.Y(n_2069)
);

CKINVDCx20_ASAP7_75t_R g2070 ( 
.A(n_1272),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_1447),
.Y(n_2071)
);

CKINVDCx16_ASAP7_75t_R g2072 ( 
.A(n_1658),
.Y(n_2072)
);

CKINVDCx20_ASAP7_75t_R g2073 ( 
.A(n_1272),
.Y(n_2073)
);

CKINVDCx20_ASAP7_75t_R g2074 ( 
.A(n_1275),
.Y(n_2074)
);

CKINVDCx20_ASAP7_75t_R g2075 ( 
.A(n_1275),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1552),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1553),
.Y(n_2077)
);

CKINVDCx20_ASAP7_75t_R g2078 ( 
.A(n_1277),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1554),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_1447),
.Y(n_2080)
);

CKINVDCx20_ASAP7_75t_R g2081 ( 
.A(n_1277),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1556),
.Y(n_2082)
);

CKINVDCx20_ASAP7_75t_R g2083 ( 
.A(n_1279),
.Y(n_2083)
);

CKINVDCx20_ASAP7_75t_R g2084 ( 
.A(n_1279),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1560),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_1449),
.Y(n_2086)
);

INVx1_ASAP7_75t_SL g2087 ( 
.A(n_1282),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1565),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1707),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1925),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1830),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_2062),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1696),
.B(n_1714),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1739),
.B(n_1328),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1830),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1707),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1927),
.Y(n_2097)
);

NAND2xp33_ASAP7_75t_SL g2098 ( 
.A(n_2048),
.B(n_1083),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_1830),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1834),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1904),
.A2(n_1288),
.B1(n_1282),
.B2(n_1449),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_2069),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1709),
.Y(n_2103)
);

AND2x2_ASAP7_75t_R g2104 ( 
.A(n_1987),
.B(n_683),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_1918),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1830),
.Y(n_2106)
);

INVx5_ASAP7_75t_L g2107 ( 
.A(n_1929),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1710),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1744),
.B(n_1330),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_1929),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1905),
.B(n_1540),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1834),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1858),
.Y(n_2113)
);

INVx2_ASAP7_75t_SL g2114 ( 
.A(n_1905),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_L g2115 ( 
.A(n_1929),
.Y(n_2115)
);

BUFx6f_ASAP7_75t_L g2116 ( 
.A(n_1929),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2008),
.B(n_1540),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1928),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1768),
.B(n_1330),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_1778),
.B(n_1557),
.Y(n_2120)
);

OAI21x1_ASAP7_75t_L g2121 ( 
.A1(n_1932),
.A2(n_1365),
.B(n_1362),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1851),
.A2(n_1288),
.B1(n_1452),
.B2(n_1451),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_1795),
.B(n_1557),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1796),
.B(n_1362),
.Y(n_2124)
);

INVx2_ASAP7_75t_SL g2125 ( 
.A(n_2008),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1722),
.B(n_1934),
.Y(n_2126)
);

BUFx3_ASAP7_75t_L g2127 ( 
.A(n_2069),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1941),
.B(n_1365),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_1858),
.Y(n_2129)
);

OAI21x1_ASAP7_75t_L g2130 ( 
.A1(n_2066),
.A2(n_1434),
.B(n_1370),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_1773),
.B(n_1563),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1871),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1745),
.B(n_1370),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1712),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1713),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1711),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_1773),
.B(n_1563),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1870),
.B(n_1434),
.Y(n_2138)
);

BUFx8_ASAP7_75t_SL g2139 ( 
.A(n_1715),
.Y(n_2139)
);

AND2x4_ASAP7_75t_L g2140 ( 
.A(n_1773),
.B(n_1568),
.Y(n_2140)
);

OAI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_1804),
.A2(n_1393),
.B1(n_1356),
.B2(n_1379),
.Y(n_2141)
);

CKINVDCx11_ASAP7_75t_R g2142 ( 
.A(n_1937),
.Y(n_2142)
);

BUFx6f_ASAP7_75t_L g2143 ( 
.A(n_1865),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_1998),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_SL g2145 ( 
.A(n_1803),
.B(n_1363),
.Y(n_2145)
);

OA21x2_ASAP7_75t_L g2146 ( 
.A1(n_1819),
.A2(n_1352),
.B(n_1351),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1989),
.B(n_1451),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1708),
.Y(n_2148)
);

OA21x2_ASAP7_75t_L g2149 ( 
.A1(n_1825),
.A2(n_1353),
.B(n_1568),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1832),
.Y(n_2150)
);

OAI22xp5_ASAP7_75t_SL g2151 ( 
.A1(n_2022),
.A2(n_688),
.B1(n_886),
.B2(n_683),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1836),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1871),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1880),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1842),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1843),
.Y(n_2156)
);

AND2x2_ASAP7_75t_SL g2157 ( 
.A(n_1743),
.B(n_1649),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1880),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1845),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_SL g2160 ( 
.A(n_1945),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1849),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1850),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1915),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_1752),
.B(n_1452),
.Y(n_2164)
);

OAI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_1807),
.A2(n_1477),
.B1(n_1457),
.B2(n_1460),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1855),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2038),
.B(n_1456),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1718),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_1812),
.B(n_1577),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1915),
.Y(n_2170)
);

NAND2xp33_ASAP7_75t_L g2171 ( 
.A(n_1762),
.B(n_1437),
.Y(n_2171)
);

BUFx3_ASAP7_75t_L g2172 ( 
.A(n_1817),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_1951),
.Y(n_2173)
);

CKINVDCx20_ASAP7_75t_R g2174 ( 
.A(n_1715),
.Y(n_2174)
);

CKINVDCx6p67_ASAP7_75t_R g2175 ( 
.A(n_1937),
.Y(n_2175)
);

INVx3_ASAP7_75t_L g2176 ( 
.A(n_1938),
.Y(n_2176)
);

INVx4_ASAP7_75t_L g2177 ( 
.A(n_1951),
.Y(n_2177)
);

OAI22xp5_ASAP7_75t_SL g2178 ( 
.A1(n_2022),
.A2(n_886),
.B1(n_944),
.B2(n_688),
.Y(n_2178)
);

NOR2x1_ASAP7_75t_L g2179 ( 
.A(n_1754),
.B(n_1833),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_1951),
.Y(n_2180)
);

OAI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2045),
.A2(n_1457),
.B1(n_1460),
.B2(n_1456),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_1938),
.Y(n_2182)
);

NAND3xp33_ASAP7_75t_L g2183 ( 
.A(n_1792),
.B(n_1295),
.C(n_1233),
.Y(n_2183)
);

OAI22xp5_ASAP7_75t_SL g2184 ( 
.A1(n_2037),
.A2(n_946),
.B1(n_1137),
.B2(n_944),
.Y(n_2184)
);

HB1xp67_ASAP7_75t_L g2185 ( 
.A(n_2018),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1815),
.B(n_1463),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1719),
.Y(n_2187)
);

BUFx6f_ASAP7_75t_L g2188 ( 
.A(n_1975),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1862),
.Y(n_2189)
);

OAI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_1827),
.A2(n_1463),
.B1(n_1471),
.B2(n_1464),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1867),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1975),
.Y(n_2192)
);

INVx3_ASAP7_75t_L g2193 ( 
.A(n_2041),
.Y(n_2193)
);

HB1xp67_ASAP7_75t_L g2194 ( 
.A(n_2072),
.Y(n_2194)
);

NAND2xp33_ASAP7_75t_L g2195 ( 
.A(n_1764),
.B(n_1437),
.Y(n_2195)
);

OA21x2_ASAP7_75t_L g2196 ( 
.A1(n_1868),
.A2(n_1599),
.B(n_1577),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2041),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1873),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1877),
.Y(n_2199)
);

NAND2xp33_ASAP7_75t_L g2200 ( 
.A(n_1919),
.B(n_1437),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_SL g2201 ( 
.A1(n_2037),
.A2(n_1137),
.B1(n_1141),
.B2(n_946),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1878),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_1879),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1723),
.B(n_1464),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1882),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1887),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1891),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1893),
.Y(n_2208)
);

BUFx6f_ASAP7_75t_L g2209 ( 
.A(n_1899),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_1721),
.B(n_1599),
.Y(n_2210)
);

INVx4_ASAP7_75t_L g2211 ( 
.A(n_1900),
.Y(n_2211)
);

AOI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_1895),
.A2(n_1779),
.B1(n_1774),
.B2(n_1786),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_1908),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1909),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1866),
.B(n_1471),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1922),
.B(n_1474),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1724),
.B(n_1605),
.Y(n_2217)
);

INVx3_ASAP7_75t_L g2218 ( 
.A(n_1910),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_1911),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_2055),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1912),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_SL g2222 ( 
.A1(n_2044),
.A2(n_1151),
.B1(n_1176),
.B2(n_1141),
.Y(n_2222)
);

INVx6_ASAP7_75t_L g2223 ( 
.A(n_1945),
.Y(n_2223)
);

BUFx6f_ASAP7_75t_L g2224 ( 
.A(n_1913),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_1987),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1914),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_1917),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_1720),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1725),
.B(n_1605),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1924),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1698),
.Y(n_2231)
);

AND2x2_ASAP7_75t_SL g2232 ( 
.A(n_1783),
.B(n_1278),
.Y(n_2232)
);

BUFx6f_ASAP7_75t_L g2233 ( 
.A(n_1771),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1931),
.B(n_1474),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1700),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_1973),
.B(n_1482),
.Y(n_2236)
);

INVx3_ASAP7_75t_L g2237 ( 
.A(n_1701),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_1775),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1706),
.Y(n_2239)
);

BUFx6f_ASAP7_75t_L g2240 ( 
.A(n_1780),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1784),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1785),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1789),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1793),
.Y(n_2244)
);

BUFx12f_ASAP7_75t_L g2245 ( 
.A(n_1765),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1794),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1980),
.B(n_1482),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1798),
.Y(n_2248)
);

INVx3_ASAP7_75t_L g2249 ( 
.A(n_1800),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1801),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1802),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1944),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1728),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1729),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_1956),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1957),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1958),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2019),
.B(n_1483),
.Y(n_2258)
);

AOI22xp5_ASAP7_75t_L g2259 ( 
.A1(n_1823),
.A2(n_1484),
.B1(n_1490),
.B2(n_1483),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_1730),
.B(n_1620),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1731),
.Y(n_2261)
);

BUFx6f_ASAP7_75t_L g2262 ( 
.A(n_1959),
.Y(n_2262)
);

OAI21x1_ASAP7_75t_L g2263 ( 
.A1(n_1953),
.A2(n_1687),
.B(n_1681),
.Y(n_2263)
);

BUFx2_ASAP7_75t_L g2264 ( 
.A(n_2064),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1960),
.Y(n_2265)
);

INVx3_ASAP7_75t_L g2266 ( 
.A(n_1961),
.Y(n_2266)
);

BUFx6f_ASAP7_75t_L g2267 ( 
.A(n_1962),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_1964),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1732),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1734),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_1965),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1966),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_1736),
.B(n_1620),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1737),
.Y(n_2274)
);

BUFx6f_ASAP7_75t_L g2275 ( 
.A(n_1968),
.Y(n_2275)
);

OA21x2_ASAP7_75t_L g2276 ( 
.A1(n_1738),
.A2(n_1639),
.B(n_1635),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1740),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2057),
.B(n_1484),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1741),
.Y(n_2279)
);

INVx6_ASAP7_75t_L g2280 ( 
.A(n_1945),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_1838),
.B(n_1490),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_1974),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1742),
.Y(n_2283)
);

NAND2xp33_ASAP7_75t_L g2284 ( 
.A(n_2023),
.B(n_1437),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_1976),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1746),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1979),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_1841),
.A2(n_1805),
.B1(n_1751),
.B2(n_1733),
.Y(n_2288)
);

OAI22xp5_ASAP7_75t_SL g2289 ( 
.A1(n_2044),
.A2(n_1176),
.B1(n_1186),
.B2(n_1151),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_1726),
.Y(n_2290)
);

BUFx3_ASAP7_75t_L g2291 ( 
.A(n_1747),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_1749),
.B(n_1635),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_1901),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1903),
.B(n_1491),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1906),
.B(n_1491),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1750),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_1982),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_1984),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1985),
.Y(n_2299)
);

INVx5_ASAP7_75t_L g2300 ( 
.A(n_1963),
.Y(n_2300)
);

AND2x6_ASAP7_75t_L g2301 ( 
.A(n_1753),
.B(n_968),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1755),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1758),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_1761),
.B(n_1639),
.Y(n_2304)
);

BUFx6f_ASAP7_75t_L g2305 ( 
.A(n_1986),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1991),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1763),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_1946),
.B(n_1493),
.Y(n_2308)
);

OAI21x1_ASAP7_75t_L g2309 ( 
.A1(n_1767),
.A2(n_1694),
.B(n_1665),
.Y(n_2309)
);

INVx6_ASAP7_75t_L g2310 ( 
.A(n_1963),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_1992),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_1995),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_1950),
.B(n_1493),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1769),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_1955),
.B(n_1495),
.Y(n_2315)
);

XNOR2x2_ASAP7_75t_L g2316 ( 
.A(n_2087),
.B(n_671),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1999),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2001),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_L g2319 ( 
.A(n_2003),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2005),
.B(n_1643),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2007),
.Y(n_2321)
);

OAI22xp5_ASAP7_75t_SL g2322 ( 
.A1(n_2050),
.A2(n_1196),
.B1(n_1204),
.B2(n_1186),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_1840),
.B(n_1881),
.Y(n_2323)
);

INVx3_ASAP7_75t_L g2324 ( 
.A(n_2009),
.Y(n_2324)
);

INVxp67_ASAP7_75t_L g2325 ( 
.A(n_1816),
.Y(n_2325)
);

OAI21x1_ASAP7_75t_L g2326 ( 
.A1(n_2017),
.A2(n_1694),
.B(n_1665),
.Y(n_2326)
);

BUFx6f_ASAP7_75t_L g2327 ( 
.A(n_2020),
.Y(n_2327)
);

INVxp67_ASAP7_75t_L g2328 ( 
.A(n_1839),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_2011),
.B(n_1495),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2024),
.Y(n_2330)
);

OA21x2_ASAP7_75t_L g2331 ( 
.A1(n_2025),
.A2(n_1669),
.B(n_1643),
.Y(n_2331)
);

AND2x4_ASAP7_75t_L g2332 ( 
.A(n_2042),
.B(n_1669),
.Y(n_2332)
);

BUFx12f_ASAP7_75t_L g2333 ( 
.A(n_1765),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2026),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2027),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_2028),
.B(n_1673),
.Y(n_2336)
);

OAI22xp5_ASAP7_75t_L g2337 ( 
.A1(n_1733),
.A2(n_1500),
.B1(n_1503),
.B2(n_1496),
.Y(n_2337)
);

INVx4_ASAP7_75t_L g2338 ( 
.A(n_2029),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2060),
.B(n_1496),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2030),
.B(n_1500),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2032),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_2034),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2035),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_2036),
.B(n_1673),
.Y(n_2344)
);

INVx4_ASAP7_75t_L g2345 ( 
.A(n_2039),
.Y(n_2345)
);

HB1xp67_ASAP7_75t_L g2346 ( 
.A(n_1757),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2043),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2053),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2056),
.Y(n_2349)
);

INVx6_ASAP7_75t_L g2350 ( 
.A(n_1963),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2058),
.B(n_1503),
.Y(n_2351)
);

AOI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_1751),
.A2(n_1510),
.B1(n_1514),
.B2(n_1506),
.Y(n_2352)
);

INVx4_ASAP7_75t_L g2353 ( 
.A(n_2061),
.Y(n_2353)
);

OAI21x1_ASAP7_75t_L g2354 ( 
.A1(n_2076),
.A2(n_1687),
.B(n_1681),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2077),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2079),
.B(n_1506),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2082),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2085),
.Y(n_2358)
);

BUFx8_ASAP7_75t_L g2359 ( 
.A(n_1857),
.Y(n_2359)
);

AOI22xp5_ASAP7_75t_L g2360 ( 
.A1(n_1854),
.A2(n_1514),
.B1(n_1516),
.B2(n_1510),
.Y(n_2360)
);

BUFx2_ASAP7_75t_L g2361 ( 
.A(n_1888),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2088),
.B(n_1505),
.Y(n_2362)
);

INVx3_ASAP7_75t_L g2363 ( 
.A(n_1790),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_1952),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1971),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2013),
.Y(n_2366)
);

OA21x2_ASAP7_75t_L g2367 ( 
.A1(n_1996),
.A2(n_1632),
.B(n_1575),
.Y(n_2367)
);

AND2x4_ASAP7_75t_L g2368 ( 
.A(n_1766),
.B(n_1569),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_1770),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1772),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_1781),
.Y(n_2371)
);

INVx3_ASAP7_75t_L g2372 ( 
.A(n_1787),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_1788),
.B(n_1516),
.Y(n_2373)
);

BUFx6f_ASAP7_75t_L g2374 ( 
.A(n_1791),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_1797),
.Y(n_2375)
);

OAI21x1_ASAP7_75t_L g2376 ( 
.A1(n_1949),
.A2(n_1326),
.B(n_1278),
.Y(n_2376)
);

CKINVDCx6p67_ASAP7_75t_R g2377 ( 
.A(n_1818),
.Y(n_2377)
);

OAI22xp5_ASAP7_75t_SL g2378 ( 
.A1(n_2050),
.A2(n_1204),
.B1(n_1209),
.B2(n_1196),
.Y(n_2378)
);

INVx6_ASAP7_75t_L g2379 ( 
.A(n_1848),
.Y(n_2379)
);

BUFx8_ASAP7_75t_L g2380 ( 
.A(n_1848),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_1806),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_1808),
.Y(n_2382)
);

OAI21x1_ASAP7_75t_L g2383 ( 
.A1(n_1809),
.A2(n_1653),
.B(n_1326),
.Y(n_2383)
);

BUFx2_ASAP7_75t_L g2384 ( 
.A(n_1759),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1810),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_1813),
.B(n_1517),
.Y(n_2386)
);

HB1xp67_ASAP7_75t_L g2387 ( 
.A(n_1759),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1820),
.Y(n_2388)
);

OA21x2_ASAP7_75t_L g2389 ( 
.A1(n_2068),
.A2(n_1579),
.B(n_1578),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_1824),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_1826),
.Y(n_2391)
);

INVx3_ASAP7_75t_L g2392 ( 
.A(n_1828),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_1829),
.B(n_1517),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_1831),
.B(n_1524),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1835),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_1837),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_1844),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_1846),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1847),
.Y(n_2399)
);

INVx4_ASAP7_75t_L g2400 ( 
.A(n_1856),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_1859),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_1860),
.Y(n_2402)
);

INVx5_ASAP7_75t_L g2403 ( 
.A(n_1864),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_1869),
.Y(n_2404)
);

INVxp33_ASAP7_75t_L g2405 ( 
.A(n_1716),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_1874),
.B(n_1505),
.Y(n_2406)
);

HB1xp67_ASAP7_75t_L g2407 ( 
.A(n_1875),
.Y(n_2407)
);

OA21x2_ASAP7_75t_L g2408 ( 
.A1(n_2068),
.A2(n_1590),
.B(n_1584),
.Y(n_2408)
);

CKINVDCx5p33_ASAP7_75t_R g2409 ( 
.A(n_1748),
.Y(n_2409)
);

AOI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_1876),
.A2(n_1532),
.B1(n_1539),
.B2(n_1524),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_1883),
.B(n_1505),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_1884),
.Y(n_2412)
);

CKINVDCx20_ASAP7_75t_R g2413 ( 
.A(n_1716),
.Y(n_2413)
);

AND2x2_ASAP7_75t_SL g2414 ( 
.A(n_2086),
.B(n_1653),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_1889),
.B(n_1532),
.Y(n_2415)
);

INVx3_ASAP7_75t_L g2416 ( 
.A(n_1890),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_1894),
.B(n_1625),
.Y(n_2417)
);

BUFx12f_ASAP7_75t_L g2418 ( 
.A(n_1892),
.Y(n_2418)
);

NAND2xp33_ASAP7_75t_L g2419 ( 
.A(n_2071),
.B(n_1437),
.Y(n_2419)
);

AND2x2_ASAP7_75t_SL g2420 ( 
.A(n_2071),
.B(n_1667),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1896),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_1897),
.B(n_1539),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_1898),
.Y(n_2423)
);

OAI21x1_ASAP7_75t_L g2424 ( 
.A1(n_1902),
.A2(n_1667),
.B(n_1175),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_1907),
.Y(n_2425)
);

OAI21x1_ASAP7_75t_L g2426 ( 
.A1(n_1916),
.A2(n_1175),
.B(n_1123),
.Y(n_2426)
);

BUFx3_ASAP7_75t_L g2427 ( 
.A(n_1920),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_1930),
.Y(n_2428)
);

BUFx6f_ASAP7_75t_L g2429 ( 
.A(n_1933),
.Y(n_2429)
);

NOR2x1_ASAP7_75t_L g2430 ( 
.A(n_2052),
.B(n_1555),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_1935),
.B(n_1547),
.Y(n_2431)
);

BUFx2_ASAP7_75t_L g2432 ( 
.A(n_2052),
.Y(n_2432)
);

INVx6_ASAP7_75t_L g2433 ( 
.A(n_1852),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_1936),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_1939),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_1940),
.B(n_1547),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_1948),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_1954),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_1967),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_1969),
.B(n_1548),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_1972),
.B(n_1548),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_1977),
.B(n_1549),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_1988),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_1993),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_1994),
.Y(n_2445)
);

INVx3_ASAP7_75t_L g2446 ( 
.A(n_1997),
.Y(n_2446)
);

AND2x4_ASAP7_75t_L g2447 ( 
.A(n_2000),
.B(n_1591),
.Y(n_2447)
);

INVx3_ASAP7_75t_L g2448 ( 
.A(n_2004),
.Y(n_2448)
);

HB1xp67_ASAP7_75t_L g2449 ( 
.A(n_2006),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2010),
.Y(n_2450)
);

AOI22x1_ASAP7_75t_SL g2451 ( 
.A1(n_1697),
.A2(n_1209),
.B1(n_674),
.B2(n_698),
.Y(n_2451)
);

AOI22xp5_ASAP7_75t_L g2452 ( 
.A1(n_2012),
.A2(n_1551),
.B1(n_1559),
.B2(n_1549),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2021),
.B(n_1551),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2031),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2033),
.B(n_1625),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2040),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2046),
.Y(n_2457)
);

AND2x4_ASAP7_75t_L g2458 ( 
.A(n_2047),
.B(n_1593),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2049),
.Y(n_2459)
);

NAND2xp33_ASAP7_75t_L g2460 ( 
.A(n_2080),
.B(n_1437),
.Y(n_2460)
);

INVx2_ASAP7_75t_SL g2461 ( 
.A(n_2051),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2059),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_2065),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2080),
.Y(n_2464)
);

BUFx3_ASAP7_75t_L g2465 ( 
.A(n_2086),
.Y(n_2465)
);

HB1xp67_ASAP7_75t_L g2466 ( 
.A(n_1695),
.Y(n_2466)
);

BUFx2_ASAP7_75t_L g2467 ( 
.A(n_2054),
.Y(n_2467)
);

BUFx3_ASAP7_75t_L g2468 ( 
.A(n_1717),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_1892),
.Y(n_2469)
);

BUFx6f_ASAP7_75t_L g2470 ( 
.A(n_1695),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_1699),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_1852),
.Y(n_2472)
);

BUFx6f_ASAP7_75t_L g2473 ( 
.A(n_1699),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2054),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_1702),
.B(n_1625),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_1702),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_1703),
.Y(n_2477)
);

INVx5_ASAP7_75t_L g2478 ( 
.A(n_1703),
.Y(n_2478)
);

BUFx12f_ASAP7_75t_L g2479 ( 
.A(n_1704),
.Y(n_2479)
);

HB1xp67_ASAP7_75t_L g2480 ( 
.A(n_1704),
.Y(n_2480)
);

BUFx6f_ASAP7_75t_L g2481 ( 
.A(n_1756),
.Y(n_2481)
);

INVx3_ASAP7_75t_L g2482 ( 
.A(n_1756),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2063),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2063),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2067),
.Y(n_2485)
);

AOI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2067),
.A2(n_1561),
.B1(n_1562),
.B2(n_1559),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2070),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2070),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2073),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2074),
.Y(n_2490)
);

INVx3_ASAP7_75t_L g2491 ( 
.A(n_2074),
.Y(n_2491)
);

AOI22x1_ASAP7_75t_SL g2492 ( 
.A1(n_1697),
.A2(n_674),
.B1(n_698),
.B2(n_673),
.Y(n_2492)
);

AOI22xp5_ASAP7_75t_L g2493 ( 
.A1(n_2075),
.A2(n_1562),
.B1(n_1564),
.B2(n_1561),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2075),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2078),
.Y(n_2495)
);

BUFx6f_ASAP7_75t_L g2496 ( 
.A(n_2078),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2081),
.Y(n_2497)
);

INVx3_ASAP7_75t_L g2498 ( 
.A(n_2081),
.Y(n_2498)
);

OAI22x1_ASAP7_75t_R g2499 ( 
.A1(n_1885),
.A2(n_1567),
.B1(n_1570),
.B2(n_1564),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2083),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2083),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2084),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2084),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_1942),
.B(n_1567),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_1717),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_1727),
.Y(n_2506)
);

AND2x4_ASAP7_75t_L g2507 ( 
.A(n_1942),
.B(n_1597),
.Y(n_2507)
);

BUFx6f_ASAP7_75t_L g2508 ( 
.A(n_1943),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_1943),
.B(n_1641),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_1947),
.B(n_1641),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_1947),
.Y(n_2511)
);

INVxp67_ASAP7_75t_L g2512 ( 
.A(n_1970),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_1970),
.B(n_1570),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2016),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2016),
.Y(n_2515)
);

INVxp67_ASAP7_75t_L g2516 ( 
.A(n_1978),
.Y(n_2516)
);

OAI21x1_ASAP7_75t_L g2517 ( 
.A1(n_1978),
.A2(n_1175),
.B(n_1123),
.Y(n_2517)
);

INVx4_ASAP7_75t_L g2518 ( 
.A(n_1981),
.Y(n_2518)
);

AND2x4_ASAP7_75t_L g2519 ( 
.A(n_1981),
.B(n_1600),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_1983),
.B(n_1601),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_1983),
.Y(n_2521)
);

OAI22xp5_ASAP7_75t_L g2522 ( 
.A1(n_1990),
.A2(n_1574),
.B1(n_1581),
.B2(n_1580),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_1990),
.Y(n_2523)
);

OAI22xp5_ASAP7_75t_SL g2524 ( 
.A1(n_2002),
.A2(n_755),
.B1(n_788),
.B2(n_673),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2002),
.Y(n_2525)
);

AOI22xp5_ASAP7_75t_SL g2526 ( 
.A1(n_2014),
.A2(n_1472),
.B1(n_1333),
.B2(n_899),
.Y(n_2526)
);

AND2x6_ASAP7_75t_L g2527 ( 
.A(n_2014),
.B(n_1123),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2015),
.B(n_1574),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2015),
.B(n_1641),
.Y(n_2529)
);

BUFx2_ASAP7_75t_L g2530 ( 
.A(n_1727),
.Y(n_2530)
);

INVx3_ASAP7_75t_L g2531 ( 
.A(n_2326),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2169),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2326),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2354),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2354),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2331),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2196),
.Y(n_2537)
);

AND2x2_ASAP7_75t_SL g2538 ( 
.A(n_2414),
.B(n_2420),
.Y(n_2538)
);

BUFx6f_ASAP7_75t_L g2539 ( 
.A(n_2331),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2196),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2196),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2196),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2331),
.Y(n_2543)
);

BUFx6f_ASAP7_75t_L g2544 ( 
.A(n_2331),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2169),
.Y(n_2545)
);

OR2x6_ASAP7_75t_L g2546 ( 
.A(n_2517),
.B(n_865),
.Y(n_2546)
);

OAI21x1_ASAP7_75t_L g2547 ( 
.A1(n_2130),
.A2(n_2263),
.B(n_2121),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2276),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2276),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2111),
.B(n_1373),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2323),
.B(n_1580),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2137),
.Y(n_2552)
);

OAI21x1_ASAP7_75t_L g2553 ( 
.A1(n_2130),
.A2(n_1610),
.B(n_1607),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2137),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2276),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2131),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2309),
.Y(n_2557)
);

INVx3_ASAP7_75t_L g2558 ( 
.A(n_2309),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2276),
.Y(n_2559)
);

BUFx6f_ASAP7_75t_L g2560 ( 
.A(n_2121),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2149),
.Y(n_2561)
);

AOI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_2419),
.A2(n_1585),
.B1(n_1586),
.B2(n_1581),
.Y(n_2562)
);

BUFx8_ASAP7_75t_L g2563 ( 
.A(n_2160),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2149),
.Y(n_2564)
);

NAND2xp33_ASAP7_75t_SL g2565 ( 
.A(n_2406),
.B(n_1585),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2149),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2149),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2089),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2368),
.B(n_1586),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2089),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_2172),
.B(n_1611),
.Y(n_2571)
);

BUFx2_ASAP7_75t_L g2572 ( 
.A(n_2105),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2096),
.Y(n_2573)
);

OA21x2_ASAP7_75t_L g2574 ( 
.A1(n_2263),
.A2(n_1613),
.B(n_1612),
.Y(n_2574)
);

INVx1_ASAP7_75t_SL g2575 ( 
.A(n_2105),
.Y(n_2575)
);

BUFx6f_ASAP7_75t_L g2576 ( 
.A(n_2173),
.Y(n_2576)
);

HB1xp67_ASAP7_75t_L g2577 ( 
.A(n_2144),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_2368),
.B(n_1595),
.Y(n_2578)
);

AND2x4_ASAP7_75t_L g2579 ( 
.A(n_2172),
.B(n_1619),
.Y(n_2579)
);

AND2x6_ASAP7_75t_L g2580 ( 
.A(n_2323),
.B(n_851),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2096),
.Y(n_2581)
);

BUFx2_ASAP7_75t_L g2582 ( 
.A(n_2092),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2100),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_2092),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2100),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2112),
.Y(n_2586)
);

BUFx6f_ASAP7_75t_L g2587 ( 
.A(n_2173),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2112),
.Y(n_2588)
);

AND2x4_ASAP7_75t_L g2589 ( 
.A(n_2120),
.B(n_1623),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2113),
.Y(n_2590)
);

INVx3_ASAP7_75t_L g2591 ( 
.A(n_2146),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2113),
.Y(n_2592)
);

HB1xp67_ASAP7_75t_L g2593 ( 
.A(n_2185),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2132),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_2281),
.B(n_1595),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2132),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2131),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2131),
.Y(n_2598)
);

BUFx6f_ASAP7_75t_L g2599 ( 
.A(n_2233),
.Y(n_2599)
);

INVx3_ASAP7_75t_L g2600 ( 
.A(n_2146),
.Y(n_2600)
);

NAND2xp33_ASAP7_75t_L g2601 ( 
.A(n_2301),
.B(n_1437),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2111),
.B(n_2117),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2153),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2117),
.B(n_2114),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2114),
.B(n_1373),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2153),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2154),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2154),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2323),
.B(n_1596),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2158),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2158),
.Y(n_2611)
);

BUFx8_ASAP7_75t_L g2612 ( 
.A(n_2160),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_2147),
.B(n_1596),
.Y(n_2613)
);

INVx3_ASAP7_75t_L g2614 ( 
.A(n_2146),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2163),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2163),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2170),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2133),
.B(n_1598),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2170),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2192),
.Y(n_2620)
);

NAND3xp33_ASAP7_75t_L g2621 ( 
.A(n_2183),
.B(n_1603),
.C(n_1598),
.Y(n_2621)
);

BUFx6f_ASAP7_75t_L g2622 ( 
.A(n_2233),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2194),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2192),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2125),
.B(n_1535),
.Y(n_2625)
);

NOR2xp33_ASAP7_75t_L g2626 ( 
.A(n_2167),
.B(n_2204),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2197),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_SL g2628 ( 
.A(n_2368),
.B(n_1603),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2197),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2146),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2140),
.Y(n_2631)
);

NAND3xp33_ASAP7_75t_L g2632 ( 
.A(n_2313),
.B(n_1606),
.C(n_1604),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2235),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2140),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_2447),
.B(n_1604),
.Y(n_2635)
);

INVxp67_ASAP7_75t_L g2636 ( 
.A(n_2220),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2235),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2235),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2140),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2181),
.B(n_1606),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2125),
.B(n_1535),
.Y(n_2641)
);

AND2x6_ASAP7_75t_L g2642 ( 
.A(n_2179),
.B(n_853),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2237),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2231),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2231),
.Y(n_2645)
);

AND2x2_ASAP7_75t_SL g2646 ( 
.A(n_2414),
.B(n_1310),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2239),
.Y(n_2647)
);

INVxp67_ASAP7_75t_L g2648 ( 
.A(n_2264),
.Y(n_2648)
);

INVx3_ASAP7_75t_L g2649 ( 
.A(n_2177),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2237),
.Y(n_2650)
);

OAI21x1_ASAP7_75t_L g2651 ( 
.A1(n_2426),
.A2(n_1629),
.B(n_1626),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2239),
.Y(n_2652)
);

NAND2xp33_ASAP7_75t_L g2653 ( 
.A(n_2301),
.B(n_1437),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2237),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2376),
.B(n_1310),
.Y(n_2655)
);

AND2x4_ASAP7_75t_L g2656 ( 
.A(n_2120),
.B(n_1633),
.Y(n_2656)
);

OR2x6_ASAP7_75t_L g2657 ( 
.A(n_2517),
.B(n_1201),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2128),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2129),
.Y(n_2659)
);

BUFx6f_ASAP7_75t_L g2660 ( 
.A(n_2233),
.Y(n_2660)
);

HB1xp67_ASAP7_75t_L g2661 ( 
.A(n_2507),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2090),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2376),
.B(n_1454),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2090),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2093),
.B(n_1608),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2097),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2097),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2129),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2129),
.Y(n_2669)
);

INVx3_ASAP7_75t_L g2670 ( 
.A(n_2177),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2118),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2118),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2176),
.Y(n_2673)
);

HB1xp67_ASAP7_75t_L g2674 ( 
.A(n_2507),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2150),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2176),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2150),
.Y(n_2677)
);

NOR2xp33_ASAP7_75t_L g2678 ( 
.A(n_2190),
.B(n_1608),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2362),
.B(n_1454),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2176),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2193),
.Y(n_2681)
);

INVxp67_ASAP7_75t_L g2682 ( 
.A(n_2264),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2193),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2152),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2152),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2155),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2155),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2193),
.Y(n_2688)
);

AOI22xp5_ASAP7_75t_L g2689 ( 
.A1(n_2419),
.A2(n_2460),
.B1(n_2389),
.B2(n_2408),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2205),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2120),
.B(n_1615),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2156),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2156),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2205),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2362),
.B(n_1508),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2159),
.Y(n_2696)
);

BUFx2_ASAP7_75t_L g2697 ( 
.A(n_2507),
.Y(n_2697)
);

OAI21x1_ASAP7_75t_L g2698 ( 
.A1(n_2426),
.A2(n_2424),
.B(n_2218),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2123),
.B(n_1615),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2389),
.B(n_1508),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2159),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2123),
.B(n_1616),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2161),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2161),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2206),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2206),
.Y(n_2706)
);

NAND2xp33_ASAP7_75t_SL g2707 ( 
.A(n_2406),
.B(n_1616),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2162),
.Y(n_2708)
);

INVx3_ASAP7_75t_L g2709 ( 
.A(n_2177),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2207),
.Y(n_2710)
);

OA21x2_ASAP7_75t_L g2711 ( 
.A1(n_2138),
.A2(n_1640),
.B(n_1634),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2123),
.B(n_1618),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2162),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2207),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_SL g2715 ( 
.A(n_2447),
.B(n_1618),
.Y(n_2715)
);

BUFx6f_ASAP7_75t_L g2716 ( 
.A(n_2233),
.Y(n_2716)
);

NAND2xp33_ASAP7_75t_SL g2717 ( 
.A(n_2411),
.B(n_1621),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2320),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2320),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2094),
.B(n_1621),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2241),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2241),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2243),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2243),
.Y(n_2724)
);

NOR2xp33_ASAP7_75t_L g2725 ( 
.A(n_2373),
.B(n_1624),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2214),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2214),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2248),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2230),
.Y(n_2729)
);

AND2x6_ASAP7_75t_L g2730 ( 
.A(n_2102),
.B(n_853),
.Y(n_2730)
);

BUFx3_ASAP7_75t_L g2731 ( 
.A(n_2102),
.Y(n_2731)
);

HB1xp67_ASAP7_75t_L g2732 ( 
.A(n_2519),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2248),
.Y(n_2733)
);

OA21x2_ASAP7_75t_L g2734 ( 
.A1(n_2109),
.A2(n_2124),
.B(n_2119),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2249),
.B(n_1624),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2389),
.B(n_1243),
.Y(n_2736)
);

AND2x4_ASAP7_75t_L g2737 ( 
.A(n_2250),
.B(n_1644),
.Y(n_2737)
);

OA21x2_ASAP7_75t_L g2738 ( 
.A1(n_2126),
.A2(n_1650),
.B(n_1647),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2230),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2249),
.B(n_1628),
.Y(n_2740)
);

BUFx6f_ASAP7_75t_L g2741 ( 
.A(n_2233),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2250),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2166),
.Y(n_2743)
);

OAI21x1_ASAP7_75t_L g2744 ( 
.A1(n_2424),
.A2(n_1652),
.B(n_1651),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2251),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2166),
.Y(n_2746)
);

AND2x4_ASAP7_75t_L g2747 ( 
.A(n_2251),
.B(n_1662),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2317),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2189),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2317),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2318),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2318),
.B(n_1663),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2519),
.Y(n_2753)
);

NAND2xp33_ASAP7_75t_SL g2754 ( 
.A(n_2411),
.B(n_1628),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2321),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2189),
.Y(n_2756)
);

OAI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2215),
.A2(n_1637),
.B1(n_1642),
.B2(n_1638),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2389),
.B(n_1271),
.Y(n_2758)
);

BUFx2_ASAP7_75t_L g2759 ( 
.A(n_2519),
.Y(n_2759)
);

BUFx2_ASAP7_75t_L g2760 ( 
.A(n_2520),
.Y(n_2760)
);

INVx3_ASAP7_75t_L g2761 ( 
.A(n_2143),
.Y(n_2761)
);

OR2x2_ASAP7_75t_L g2762 ( 
.A(n_2225),
.B(n_1350),
.Y(n_2762)
);

INVx3_ASAP7_75t_L g2763 ( 
.A(n_2143),
.Y(n_2763)
);

BUFx2_ASAP7_75t_L g2764 ( 
.A(n_2520),
.Y(n_2764)
);

BUFx6f_ASAP7_75t_L g2765 ( 
.A(n_2238),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2191),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2191),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2198),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2143),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2255),
.B(n_1637),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2321),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2198),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2255),
.B(n_1638),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2408),
.B(n_1263),
.Y(n_2774)
);

INVx3_ASAP7_75t_L g2775 ( 
.A(n_2143),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2330),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2330),
.Y(n_2777)
);

HB1xp67_ASAP7_75t_L g2778 ( 
.A(n_2520),
.Y(n_2778)
);

OAI22xp5_ASAP7_75t_SL g2779 ( 
.A1(n_2151),
.A2(n_1872),
.B1(n_1735),
.B2(n_1776),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2148),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2148),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_2447),
.B(n_1642),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2199),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2199),
.Y(n_2784)
);

BUFx6f_ASAP7_75t_L g2785 ( 
.A(n_2238),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2202),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2202),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2208),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2208),
.Y(n_2789)
);

BUFx6f_ASAP7_75t_L g2790 ( 
.A(n_2238),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2221),
.Y(n_2791)
);

INVx3_ASAP7_75t_L g2792 ( 
.A(n_2143),
.Y(n_2792)
);

HB1xp67_ASAP7_75t_L g2793 ( 
.A(n_2408),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2221),
.Y(n_2794)
);

CKINVDCx20_ASAP7_75t_R g2795 ( 
.A(n_2174),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2273),
.Y(n_2796)
);

BUFx6f_ASAP7_75t_L g2797 ( 
.A(n_2238),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2244),
.Y(n_2798)
);

BUFx6f_ASAP7_75t_L g2799 ( 
.A(n_2238),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_SL g2800 ( 
.A(n_2458),
.B(n_2300),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2244),
.Y(n_2801)
);

BUFx2_ASAP7_75t_L g2802 ( 
.A(n_2527),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2246),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2273),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2246),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2252),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2273),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2408),
.B(n_1263),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2336),
.Y(n_2809)
);

XNOR2xp5_ASAP7_75t_L g2810 ( 
.A(n_2178),
.B(n_1735),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2336),
.Y(n_2811)
);

OAI22xp5_ASAP7_75t_SL g2812 ( 
.A1(n_2184),
.A2(n_2222),
.B1(n_2289),
.B2(n_2201),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2252),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2420),
.B(n_1263),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2256),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2256),
.Y(n_2816)
);

AND2x4_ASAP7_75t_L g2817 ( 
.A(n_2291),
.B(n_1664),
.Y(n_2817)
);

AND2x4_ASAP7_75t_L g2818 ( 
.A(n_2291),
.B(n_1672),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2253),
.Y(n_2819)
);

BUFx6f_ASAP7_75t_L g2820 ( 
.A(n_2240),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2253),
.Y(n_2821)
);

AND2x4_ASAP7_75t_L g2822 ( 
.A(n_2335),
.B(n_1674),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2254),
.Y(n_2823)
);

CKINVDCx16_ASAP7_75t_R g2824 ( 
.A(n_2174),
.Y(n_2824)
);

BUFx6f_ASAP7_75t_L g2825 ( 
.A(n_2240),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2257),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2257),
.Y(n_2827)
);

AND2x4_ASAP7_75t_L g2828 ( 
.A(n_2341),
.B(n_1676),
.Y(n_2828)
);

HB1xp67_ASAP7_75t_L g2829 ( 
.A(n_2458),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2254),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2261),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2261),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2286),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2286),
.Y(n_2834)
);

AND2x4_ASAP7_75t_L g2835 ( 
.A(n_2348),
.B(n_2355),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2336),
.Y(n_2836)
);

CKINVDCx20_ASAP7_75t_R g2837 ( 
.A(n_2413),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2344),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_2139),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2307),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2307),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2314),
.Y(n_2842)
);

OA21x2_ASAP7_75t_L g2843 ( 
.A1(n_2314),
.A2(n_1679),
.B(n_1677),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2265),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2266),
.B(n_1646),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2265),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2344),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2282),
.B(n_1646),
.Y(n_2848)
);

BUFx2_ASAP7_75t_L g2849 ( 
.A(n_2527),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2268),
.Y(n_2850)
);

OAI22xp5_ASAP7_75t_SL g2851 ( 
.A1(n_2322),
.A2(n_1822),
.B1(n_1853),
.B2(n_1821),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2344),
.Y(n_2852)
);

BUFx2_ASAP7_75t_L g2853 ( 
.A(n_2527),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2210),
.Y(n_2854)
);

BUFx6f_ASAP7_75t_L g2855 ( 
.A(n_2240),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_SL g2856 ( 
.A(n_2458),
.B(n_1648),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2268),
.Y(n_2857)
);

HB1xp67_ASAP7_75t_L g2858 ( 
.A(n_2293),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2210),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2272),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2272),
.Y(n_2861)
);

BUFx3_ASAP7_75t_L g2862 ( 
.A(n_2127),
.Y(n_2862)
);

BUFx6f_ASAP7_75t_L g2863 ( 
.A(n_2240),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2217),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2287),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2282),
.B(n_1648),
.Y(n_2866)
);

OAI21x1_ASAP7_75t_L g2867 ( 
.A1(n_2203),
.A2(n_1686),
.B(n_1685),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2217),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2287),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2229),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2298),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2282),
.B(n_1654),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2298),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2232),
.B(n_1267),
.Y(n_2874)
);

BUFx2_ASAP7_75t_L g2875 ( 
.A(n_2527),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2229),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2299),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2299),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_SL g2879 ( 
.A(n_2300),
.B(n_1654),
.Y(n_2879)
);

OAI21x1_ASAP7_75t_L g2880 ( 
.A1(n_2203),
.A2(n_1689),
.B(n_1688),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2306),
.Y(n_2881)
);

BUFx2_ASAP7_75t_L g2882 ( 
.A(n_2527),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2311),
.B(n_1655),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2306),
.Y(n_2884)
);

OAI22xp5_ASAP7_75t_L g2885 ( 
.A1(n_2216),
.A2(n_2247),
.B1(n_2258),
.B2(n_2234),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2312),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2312),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2334),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2334),
.Y(n_2889)
);

AND2x2_ASAP7_75t_L g2890 ( 
.A(n_2232),
.B(n_1267),
.Y(n_2890)
);

AOI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2460),
.A2(n_1655),
.B1(n_1657),
.B2(n_1656),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2343),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2260),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2311),
.B(n_1656),
.Y(n_2894)
);

HB1xp67_ASAP7_75t_L g2895 ( 
.A(n_2367),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2260),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2343),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2347),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2311),
.B(n_1657),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2347),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2349),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2292),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2349),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2357),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2292),
.Y(n_2905)
);

BUFx3_ASAP7_75t_L g2906 ( 
.A(n_2127),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2357),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_L g2908 ( 
.A(n_2240),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_2367),
.B(n_1267),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2304),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2304),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2203),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2218),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2182),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2218),
.Y(n_2915)
);

OAI21x1_ASAP7_75t_L g2916 ( 
.A1(n_2091),
.A2(n_1691),
.B(n_1690),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2324),
.Y(n_2917)
);

OA21x2_ASAP7_75t_L g2918 ( 
.A1(n_2358),
.A2(n_2108),
.B(n_2103),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2182),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2324),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2182),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2324),
.Y(n_2922)
);

CKINVDCx5p33_ASAP7_75t_R g2923 ( 
.A(n_2139),
.Y(n_2923)
);

BUFx8_ASAP7_75t_L g2924 ( 
.A(n_2160),
.Y(n_2924)
);

INVx3_ASAP7_75t_L g2925 ( 
.A(n_2180),
.Y(n_2925)
);

NAND2xp33_ASAP7_75t_SL g2926 ( 
.A(n_2417),
.B(n_1660),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2134),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2135),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2187),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2269),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2270),
.Y(n_2931)
);

NOR2xp33_ASAP7_75t_L g2932 ( 
.A(n_2386),
.B(n_1660),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2182),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2274),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2182),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2277),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2279),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2283),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2296),
.Y(n_2939)
);

BUFx6f_ASAP7_75t_L g2940 ( 
.A(n_2242),
.Y(n_2940)
);

AOI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2157),
.A2(n_1671),
.B1(n_1680),
.B2(n_1675),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2302),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2303),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2180),
.Y(n_2944)
);

BUFx6f_ASAP7_75t_L g2945 ( 
.A(n_2242),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_2300),
.B(n_1671),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2188),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2188),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2188),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2188),
.Y(n_2950)
);

INVx3_ASAP7_75t_L g2951 ( 
.A(n_2188),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2209),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2209),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2091),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2209),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2209),
.Y(n_2956)
);

INVx3_ASAP7_75t_L g2957 ( 
.A(n_2091),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2209),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2213),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_SL g2960 ( 
.A(n_2300),
.B(n_1675),
.Y(n_2960)
);

AND2x4_ASAP7_75t_L g2961 ( 
.A(n_2338),
.B(n_1692),
.Y(n_2961)
);

NAND2xp33_ASAP7_75t_SL g2962 ( 
.A(n_2417),
.B(n_1680),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2211),
.B(n_1683),
.Y(n_2963)
);

BUFx6f_ASAP7_75t_L g2964 ( 
.A(n_2242),
.Y(n_2964)
);

NOR2x1_ASAP7_75t_L g2965 ( 
.A(n_2361),
.B(n_1609),
.Y(n_2965)
);

BUFx6f_ASAP7_75t_L g2966 ( 
.A(n_2242),
.Y(n_2966)
);

BUFx6f_ASAP7_75t_L g2967 ( 
.A(n_2242),
.Y(n_2967)
);

INVx6_ASAP7_75t_L g2968 ( 
.A(n_2338),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2338),
.Y(n_2969)
);

BUFx6f_ASAP7_75t_L g2970 ( 
.A(n_2262),
.Y(n_2970)
);

OA21x2_ASAP7_75t_L g2971 ( 
.A1(n_2383),
.A2(n_1693),
.B(n_866),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2626),
.B(n_2367),
.Y(n_2972)
);

BUFx6f_ASAP7_75t_L g2973 ( 
.A(n_2539),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2631),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2631),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2561),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2634),
.Y(n_2977)
);

AND2x2_ASAP7_75t_SL g2978 ( 
.A(n_2538),
.B(n_2157),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2602),
.B(n_2367),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_SL g2980 ( 
.A(n_2538),
.B(n_2300),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2560),
.Y(n_2981)
);

INVx5_ASAP7_75t_L g2982 ( 
.A(n_2539),
.Y(n_2982)
);

AND2x4_ASAP7_75t_L g2983 ( 
.A(n_2604),
.B(n_2403),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2583),
.Y(n_2984)
);

INVx3_ASAP7_75t_L g2985 ( 
.A(n_2560),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2658),
.B(n_2315),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2634),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2583),
.Y(n_2988)
);

BUFx3_ASAP7_75t_L g2989 ( 
.A(n_2572),
.Y(n_2989)
);

INVxp67_ASAP7_75t_L g2990 ( 
.A(n_2572),
.Y(n_2990)
);

AOI22xp33_ASAP7_75t_L g2991 ( 
.A1(n_2793),
.A2(n_2301),
.B1(n_2211),
.B2(n_2267),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2561),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2564),
.Y(n_2993)
);

AND2x2_ASAP7_75t_SL g2994 ( 
.A(n_2646),
.B(n_2470),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2658),
.B(n_2329),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2854),
.B(n_2455),
.Y(n_2996)
);

OR2x6_ASAP7_75t_L g2997 ( 
.A(n_2802),
.B(n_2849),
.Y(n_2997)
);

INVx1_ASAP7_75t_SL g2998 ( 
.A(n_2575),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2564),
.Y(n_2999)
);

XOR2xp5_ASAP7_75t_L g3000 ( 
.A(n_2810),
.B(n_1760),
.Y(n_3000)
);

INVx4_ASAP7_75t_L g3001 ( 
.A(n_2599),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2639),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2639),
.Y(n_3003)
);

NAND2xp33_ASAP7_75t_SL g3004 ( 
.A(n_2802),
.B(n_2374),
.Y(n_3004)
);

INVx3_ASAP7_75t_L g3005 ( 
.A(n_2560),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2854),
.B(n_2345),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2859),
.B(n_2345),
.Y(n_3007)
);

AOI22xp33_ASAP7_75t_L g3008 ( 
.A1(n_2700),
.A2(n_2301),
.B1(n_2211),
.B2(n_2267),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_SL g3009 ( 
.A(n_2735),
.B(n_2403),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2566),
.Y(n_3010)
);

NOR2x1p5_ASAP7_75t_L g3011 ( 
.A(n_2551),
.B(n_2377),
.Y(n_3011)
);

AOI22xp5_ASAP7_75t_L g3012 ( 
.A1(n_2885),
.A2(n_2164),
.B1(n_2353),
.B2(n_2345),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2566),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2556),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2567),
.Y(n_3015)
);

BUFx6f_ASAP7_75t_L g3016 ( 
.A(n_2539),
.Y(n_3016)
);

AND2x4_ASAP7_75t_L g3017 ( 
.A(n_2731),
.B(n_2403),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2859),
.B(n_2353),
.Y(n_3018)
);

BUFx3_ASAP7_75t_L g3019 ( 
.A(n_2731),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_L g3020 ( 
.A(n_2595),
.B(n_2415),
.Y(n_3020)
);

INVx4_ASAP7_75t_L g3021 ( 
.A(n_2599),
.Y(n_3021)
);

OR2x2_ASAP7_75t_L g3022 ( 
.A(n_2762),
.B(n_2165),
.Y(n_3022)
);

AOI22xp33_ASAP7_75t_L g3023 ( 
.A1(n_2700),
.A2(n_2301),
.B1(n_2267),
.B2(n_2271),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2864),
.B(n_2353),
.Y(n_3024)
);

AND2x2_ASAP7_75t_SL g3025 ( 
.A(n_2646),
.B(n_2470),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2597),
.Y(n_3026)
);

INVx1_ASAP7_75t_SL g3027 ( 
.A(n_2582),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2598),
.Y(n_3028)
);

AOI22xp33_ASAP7_75t_L g3029 ( 
.A1(n_2736),
.A2(n_2301),
.B1(n_2267),
.B2(n_2271),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2796),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2567),
.Y(n_3031)
);

INVx2_ASAP7_75t_SL g3032 ( 
.A(n_2582),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2796),
.Y(n_3033)
);

INVx3_ASAP7_75t_L g3034 ( 
.A(n_2560),
.Y(n_3034)
);

NOR2xp33_ASAP7_75t_L g3035 ( 
.A(n_2613),
.B(n_2393),
.Y(n_3035)
);

NOR2xp33_ASAP7_75t_L g3036 ( 
.A(n_2665),
.B(n_2725),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2568),
.Y(n_3037)
);

NAND3xp33_ASAP7_75t_L g3038 ( 
.A(n_2640),
.B(n_2259),
.C(n_2410),
.Y(n_3038)
);

INVx2_ASAP7_75t_L g3039 ( 
.A(n_2568),
.Y(n_3039)
);

OAI22xp33_ASAP7_75t_L g3040 ( 
.A1(n_2675),
.A2(n_2464),
.B1(n_2280),
.B2(n_2310),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2585),
.Y(n_3041)
);

INVx3_ASAP7_75t_L g3042 ( 
.A(n_2560),
.Y(n_3042)
);

OR2x2_ASAP7_75t_L g3043 ( 
.A(n_2762),
.B(n_2528),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2570),
.Y(n_3044)
);

AOI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_2736),
.A2(n_2267),
.B1(n_2271),
.B2(n_2262),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2864),
.B(n_2262),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2868),
.B(n_2262),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2570),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2585),
.Y(n_3049)
);

INVx2_ASAP7_75t_SL g3050 ( 
.A(n_2605),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2804),
.Y(n_3051)
);

NOR2xp33_ASAP7_75t_L g3052 ( 
.A(n_2932),
.B(n_2394),
.Y(n_3052)
);

AND3x2_ASAP7_75t_L g3053 ( 
.A(n_2678),
.B(n_2361),
.C(n_2145),
.Y(n_3053)
);

AND3x2_ASAP7_75t_L g3054 ( 
.A(n_2829),
.B(n_2467),
.C(n_2432),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2586),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2586),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2573),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2868),
.B(n_2455),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2588),
.Y(n_3059)
);

BUFx6f_ASAP7_75t_SL g3060 ( 
.A(n_2862),
.Y(n_3060)
);

OR2x6_ASAP7_75t_L g3061 ( 
.A(n_2849),
.B(n_2853),
.Y(n_3061)
);

NAND3xp33_ASAP7_75t_L g3062 ( 
.A(n_2562),
.B(n_2452),
.C(n_2122),
.Y(n_3062)
);

AND2x2_ASAP7_75t_L g3063 ( 
.A(n_2870),
.B(n_2464),
.Y(n_3063)
);

OAI22xp33_ASAP7_75t_SL g3064 ( 
.A1(n_2691),
.A2(n_2280),
.B1(n_2310),
.B2(n_2223),
.Y(n_3064)
);

INVx1_ASAP7_75t_SL g3065 ( 
.A(n_2577),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_2870),
.B(n_2876),
.Y(n_3066)
);

OA22x2_ASAP7_75t_L g3067 ( 
.A1(n_2812),
.A2(n_2383),
.B1(n_2378),
.B2(n_2524),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2648),
.B(n_2422),
.Y(n_3068)
);

INVx1_ASAP7_75t_SL g3069 ( 
.A(n_2584),
.Y(n_3069)
);

AOI22xp33_ASAP7_75t_L g3070 ( 
.A1(n_2758),
.A2(n_2271),
.B1(n_2275),
.B2(n_2262),
.Y(n_3070)
);

BUFx6f_ASAP7_75t_L g3071 ( 
.A(n_2539),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2573),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2581),
.Y(n_3073)
);

INVx5_ASAP7_75t_L g3074 ( 
.A(n_2539),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2581),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_L g3076 ( 
.A(n_2682),
.B(n_2431),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2588),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2590),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_2636),
.B(n_2436),
.Y(n_3079)
);

AND2x4_ASAP7_75t_L g3080 ( 
.A(n_2862),
.B(n_2403),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2876),
.B(n_2271),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2594),
.Y(n_3082)
);

INVx1_ASAP7_75t_SL g3083 ( 
.A(n_2593),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2594),
.Y(n_3084)
);

BUFx6f_ASAP7_75t_L g3085 ( 
.A(n_2544),
.Y(n_3085)
);

BUFx8_ASAP7_75t_SL g3086 ( 
.A(n_2795),
.Y(n_3086)
);

INVx1_ASAP7_75t_SL g3087 ( 
.A(n_2623),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2804),
.Y(n_3088)
);

INVx3_ASAP7_75t_L g3089 ( 
.A(n_2957),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2893),
.B(n_2896),
.Y(n_3090)
);

AOI22xp33_ASAP7_75t_L g3091 ( 
.A1(n_2758),
.A2(n_2655),
.B1(n_2663),
.B2(n_2893),
.Y(n_3091)
);

AND2x6_ASAP7_75t_L g3092 ( 
.A(n_2537),
.B(n_2374),
.Y(n_3092)
);

OR2x6_ASAP7_75t_L g3093 ( 
.A(n_2853),
.B(n_2223),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2896),
.B(n_2275),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2590),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2902),
.B(n_2275),
.Y(n_3096)
);

NOR2xp33_ASAP7_75t_L g3097 ( 
.A(n_2618),
.B(n_2440),
.Y(n_3097)
);

CKINVDCx11_ASAP7_75t_R g3098 ( 
.A(n_2795),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2592),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2807),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2809),
.Y(n_3101)
);

AOI22xp33_ASAP7_75t_L g3102 ( 
.A1(n_2655),
.A2(n_2285),
.B1(n_2297),
.B2(n_2275),
.Y(n_3102)
);

INVx2_ASAP7_75t_SL g3103 ( 
.A(n_2605),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2809),
.Y(n_3104)
);

INVx3_ASAP7_75t_L g3105 ( 
.A(n_2957),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2592),
.Y(n_3106)
);

AND2x4_ASAP7_75t_L g3107 ( 
.A(n_2906),
.B(n_2403),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2902),
.B(n_2905),
.Y(n_3108)
);

NOR2xp33_ASAP7_75t_L g3109 ( 
.A(n_2720),
.B(n_2441),
.Y(n_3109)
);

BUFx6f_ASAP7_75t_L g3110 ( 
.A(n_2544),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2596),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2596),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2811),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_2663),
.A2(n_2285),
.B1(n_2297),
.B2(n_2275),
.Y(n_3114)
);

OR2x2_ASAP7_75t_L g3115 ( 
.A(n_2679),
.B(n_2474),
.Y(n_3115)
);

CKINVDCx5p33_ASAP7_75t_R g3116 ( 
.A(n_2839),
.Y(n_3116)
);

INVx2_ASAP7_75t_SL g3117 ( 
.A(n_2625),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2811),
.Y(n_3118)
);

NOR2xp33_ASAP7_75t_SL g3119 ( 
.A(n_2839),
.B(n_2136),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2836),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_SL g3121 ( 
.A(n_2740),
.B(n_2374),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2836),
.Y(n_3122)
);

NOR2xp33_ASAP7_75t_L g3123 ( 
.A(n_2632),
.B(n_2442),
.Y(n_3123)
);

INVx2_ASAP7_75t_SL g3124 ( 
.A(n_2625),
.Y(n_3124)
);

OAI21xp33_ASAP7_75t_SL g3125 ( 
.A1(n_2689),
.A2(n_2677),
.B(n_2675),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2838),
.Y(n_3126)
);

AOI22xp5_ASAP7_75t_L g3127 ( 
.A1(n_2969),
.A2(n_2288),
.B1(n_2278),
.B2(n_2340),
.Y(n_3127)
);

INVx3_ASAP7_75t_L g3128 ( 
.A(n_2957),
.Y(n_3128)
);

BUFx3_ASAP7_75t_L g3129 ( 
.A(n_2906),
.Y(n_3129)
);

BUFx3_ASAP7_75t_L g3130 ( 
.A(n_2697),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_2544),
.Y(n_3131)
);

AND2x2_ASAP7_75t_L g3132 ( 
.A(n_2905),
.B(n_2372),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2607),
.Y(n_3133)
);

BUFx3_ASAP7_75t_L g3134 ( 
.A(n_2697),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2607),
.Y(n_3135)
);

BUFx3_ASAP7_75t_L g3136 ( 
.A(n_2759),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2620),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2677),
.B(n_2285),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2603),
.Y(n_3139)
);

NOR2xp33_ASAP7_75t_L g3140 ( 
.A(n_2757),
.B(n_2453),
.Y(n_3140)
);

INVx5_ASAP7_75t_L g3141 ( 
.A(n_2544),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2684),
.B(n_2285),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2620),
.Y(n_3143)
);

AOI22xp33_ASAP7_75t_L g3144 ( 
.A1(n_2580),
.A2(n_2297),
.B1(n_2305),
.B2(n_2285),
.Y(n_3144)
);

CKINVDCx20_ASAP7_75t_R g3145 ( 
.A(n_2837),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2684),
.B(n_2297),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2627),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2603),
.Y(n_3148)
);

INVx4_ASAP7_75t_L g3149 ( 
.A(n_2599),
.Y(n_3149)
);

INVx2_ASAP7_75t_SL g3150 ( 
.A(n_2641),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2627),
.Y(n_3151)
);

OR2x6_ASAP7_75t_L g3152 ( 
.A(n_2875),
.B(n_2223),
.Y(n_3152)
);

INVx3_ASAP7_75t_L g3153 ( 
.A(n_2544),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_SL g3154 ( 
.A(n_2770),
.B(n_2381),
.Y(n_3154)
);

INVxp67_ASAP7_75t_SL g3155 ( 
.A(n_2649),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2537),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2540),
.Y(n_3157)
);

AOI22xp33_ASAP7_75t_L g3158 ( 
.A1(n_2580),
.A2(n_2305),
.B1(n_2319),
.B2(n_2297),
.Y(n_3158)
);

NOR2xp33_ASAP7_75t_L g3159 ( 
.A(n_2858),
.B(n_2372),
.Y(n_3159)
);

NAND3xp33_ASAP7_75t_L g3160 ( 
.A(n_2891),
.B(n_2352),
.C(n_2360),
.Y(n_3160)
);

AND2x2_ASAP7_75t_L g3161 ( 
.A(n_2550),
.B(n_2372),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2606),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2550),
.B(n_2392),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2540),
.Y(n_3164)
);

AOI22xp5_ASAP7_75t_L g3165 ( 
.A1(n_2552),
.A2(n_2554),
.B1(n_2911),
.B2(n_2910),
.Y(n_3165)
);

INVx3_ASAP7_75t_L g3166 ( 
.A(n_2649),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2541),
.Y(n_3167)
);

AO22x2_ASAP7_75t_L g3168 ( 
.A1(n_2774),
.A2(n_2451),
.B1(n_2492),
.B2(n_2104),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2838),
.Y(n_3169)
);

INVx3_ASAP7_75t_L g3170 ( 
.A(n_2649),
.Y(n_3170)
);

OA22x2_ASAP7_75t_L g3171 ( 
.A1(n_2941),
.A2(n_2493),
.B1(n_2486),
.B2(n_2212),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2847),
.Y(n_3172)
);

OAI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_2968),
.A2(n_2223),
.B1(n_2310),
.B2(n_2280),
.Y(n_3173)
);

NOR2xp33_ASAP7_75t_L g3174 ( 
.A(n_2814),
.B(n_2392),
.Y(n_3174)
);

INVx4_ASAP7_75t_L g3175 ( 
.A(n_2599),
.Y(n_3175)
);

CKINVDCx5p33_ASAP7_75t_R g3176 ( 
.A(n_2923),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_SL g3177 ( 
.A(n_2773),
.B(n_2381),
.Y(n_3177)
);

INVx3_ASAP7_75t_L g3178 ( 
.A(n_2670),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2847),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2852),
.Y(n_3180)
);

BUFx3_ASAP7_75t_L g3181 ( 
.A(n_2759),
.Y(n_3181)
);

INVx4_ASAP7_75t_L g3182 ( 
.A(n_2599),
.Y(n_3182)
);

NOR2xp33_ASAP7_75t_L g3183 ( 
.A(n_2814),
.B(n_2392),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2852),
.Y(n_3184)
);

NOR2xp33_ASAP7_75t_L g3185 ( 
.A(n_2874),
.B(n_2416),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2541),
.Y(n_3186)
);

NOR2xp33_ASAP7_75t_L g3187 ( 
.A(n_2874),
.B(n_2416),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2654),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2685),
.B(n_2305),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2542),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2542),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2548),
.Y(n_3192)
);

NAND3xp33_ASAP7_75t_L g3193 ( 
.A(n_2909),
.B(n_2101),
.C(n_2337),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2548),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2606),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2549),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2685),
.B(n_2305),
.Y(n_3197)
);

INVx3_ASAP7_75t_L g3198 ( 
.A(n_2670),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2608),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2686),
.B(n_2305),
.Y(n_3200)
);

INVx3_ASAP7_75t_L g3201 ( 
.A(n_2670),
.Y(n_3201)
);

BUFx4f_ASAP7_75t_L g3202 ( 
.A(n_2730),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_L g3203 ( 
.A(n_2890),
.B(n_2416),
.Y(n_3203)
);

INVx3_ASAP7_75t_L g3204 ( 
.A(n_2709),
.Y(n_3204)
);

CKINVDCx16_ASAP7_75t_R g3205 ( 
.A(n_2824),
.Y(n_3205)
);

AOI22xp33_ASAP7_75t_L g3206 ( 
.A1(n_2580),
.A2(n_2911),
.B1(n_2910),
.B2(n_2808),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2608),
.Y(n_3207)
);

AND2x2_ASAP7_75t_SL g3208 ( 
.A(n_2875),
.B(n_2470),
.Y(n_3208)
);

BUFx8_ASAP7_75t_SL g3209 ( 
.A(n_2837),
.Y(n_3209)
);

INVx2_ASAP7_75t_L g3210 ( 
.A(n_2549),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2686),
.B(n_2319),
.Y(n_3211)
);

INVx3_ASAP7_75t_L g3212 ( 
.A(n_2709),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2555),
.Y(n_3213)
);

BUFx8_ASAP7_75t_SL g3214 ( 
.A(n_2923),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2555),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_SL g3216 ( 
.A(n_2563),
.B(n_2136),
.Y(n_3216)
);

CKINVDCx5p33_ASAP7_75t_R g3217 ( 
.A(n_2563),
.Y(n_3217)
);

AND3x1_ASAP7_75t_L g3218 ( 
.A(n_2890),
.B(n_2515),
.C(n_2514),
.Y(n_3218)
);

INVxp33_ASAP7_75t_L g3219 ( 
.A(n_2679),
.Y(n_3219)
);

AND2x4_ASAP7_75t_L g3220 ( 
.A(n_2835),
.B(n_2478),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2687),
.B(n_2319),
.Y(n_3221)
);

BUFx6f_ASAP7_75t_L g3222 ( 
.A(n_2622),
.Y(n_3222)
);

INVx4_ASAP7_75t_L g3223 ( 
.A(n_2622),
.Y(n_3223)
);

AND2x2_ASAP7_75t_L g3224 ( 
.A(n_2695),
.B(n_2446),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2559),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2687),
.B(n_2319),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_2559),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_SL g3228 ( 
.A(n_2845),
.B(n_2381),
.Y(n_3228)
);

BUFx6f_ASAP7_75t_L g3229 ( 
.A(n_2622),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2692),
.B(n_2319),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2610),
.Y(n_3231)
);

AOI22xp33_ASAP7_75t_L g3232 ( 
.A1(n_2580),
.A2(n_2342),
.B1(n_2327),
.B2(n_2098),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2692),
.B(n_2327),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_2693),
.B(n_2327),
.Y(n_3234)
);

OR2x2_ASAP7_75t_L g3235 ( 
.A(n_2695),
.B(n_2474),
.Y(n_3235)
);

INVxp33_ASAP7_75t_L g3236 ( 
.A(n_2661),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2654),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2693),
.B(n_2696),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2610),
.Y(n_3239)
);

NOR2x1p5_ASAP7_75t_L g3240 ( 
.A(n_2609),
.B(n_2377),
.Y(n_3240)
);

AOI22xp33_ASAP7_75t_L g3241 ( 
.A1(n_2580),
.A2(n_2342),
.B1(n_2327),
.B2(n_2098),
.Y(n_3241)
);

CKINVDCx20_ASAP7_75t_R g3242 ( 
.A(n_2779),
.Y(n_3242)
);

INVx6_ASAP7_75t_L g3243 ( 
.A(n_2576),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2912),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_2611),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_SL g3246 ( 
.A(n_2848),
.B(n_2402),
.Y(n_3246)
);

INVx1_ASAP7_75t_SL g3247 ( 
.A(n_2641),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2912),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2913),
.Y(n_3249)
);

BUFx6f_ASAP7_75t_L g3250 ( 
.A(n_2622),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2913),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_SL g3252 ( 
.A(n_2866),
.B(n_2402),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_SL g3253 ( 
.A(n_2872),
.B(n_2402),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_2611),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_2718),
.B(n_2446),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_SL g3256 ( 
.A(n_2883),
.B(n_2402),
.Y(n_3256)
);

AOI22xp33_ASAP7_75t_L g3257 ( 
.A1(n_2580),
.A2(n_2808),
.B1(n_2774),
.B2(n_2746),
.Y(n_3257)
);

INVx4_ASAP7_75t_L g3258 ( 
.A(n_2622),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2915),
.Y(n_3259)
);

AOI22xp33_ASAP7_75t_L g3260 ( 
.A1(n_2743),
.A2(n_2749),
.B1(n_2756),
.B2(n_2746),
.Y(n_3260)
);

BUFx6f_ASAP7_75t_L g3261 ( 
.A(n_2660),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_2615),
.Y(n_3262)
);

OR2x6_ASAP7_75t_L g3263 ( 
.A(n_2882),
.B(n_2280),
.Y(n_3263)
);

XNOR2xp5_ASAP7_75t_L g3264 ( 
.A(n_2810),
.B(n_1760),
.Y(n_3264)
);

NOR2xp33_ASAP7_75t_L g3265 ( 
.A(n_2963),
.B(n_2446),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_2615),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_2696),
.B(n_2327),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2701),
.B(n_2342),
.Y(n_3268)
);

BUFx3_ASAP7_75t_L g3269 ( 
.A(n_2760),
.Y(n_3269)
);

AO22x2_ASAP7_75t_L g3270 ( 
.A1(n_2909),
.A2(n_2451),
.B1(n_2492),
.B2(n_1083),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_2835),
.B(n_2478),
.Y(n_3271)
);

NOR3xp33_ASAP7_75t_L g3272 ( 
.A(n_2851),
.B(n_2522),
.C(n_2513),
.Y(n_3272)
);

CKINVDCx20_ASAP7_75t_R g3273 ( 
.A(n_2563),
.Y(n_3273)
);

AND3x1_ASAP7_75t_L g3274 ( 
.A(n_2674),
.B(n_2515),
.C(n_2514),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2915),
.Y(n_3275)
);

AND2x6_ASAP7_75t_L g3276 ( 
.A(n_2630),
.B(n_2402),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2917),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2616),
.Y(n_3278)
);

BUFx6f_ASAP7_75t_L g3279 ( 
.A(n_2660),
.Y(n_3279)
);

OR2x6_ASAP7_75t_L g3280 ( 
.A(n_2882),
.B(n_2310),
.Y(n_3280)
);

INVxp33_ASAP7_75t_L g3281 ( 
.A(n_2732),
.Y(n_3281)
);

BUFx3_ASAP7_75t_L g3282 ( 
.A(n_2760),
.Y(n_3282)
);

INVxp67_ASAP7_75t_SL g3283 ( 
.A(n_2709),
.Y(n_3283)
);

BUFx3_ASAP7_75t_L g3284 ( 
.A(n_2764),
.Y(n_3284)
);

AOI22xp33_ASAP7_75t_L g3285 ( 
.A1(n_2743),
.A2(n_2342),
.B1(n_2195),
.B2(n_2200),
.Y(n_3285)
);

BUFx10_ASAP7_75t_L g3286 ( 
.A(n_2730),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_L g3287 ( 
.A(n_2894),
.B(n_2448),
.Y(n_3287)
);

INVx2_ASAP7_75t_SL g3288 ( 
.A(n_2589),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2616),
.Y(n_3289)
);

BUFx10_ASAP7_75t_L g3290 ( 
.A(n_2730),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2917),
.Y(n_3291)
);

NOR2xp33_ASAP7_75t_L g3292 ( 
.A(n_2899),
.B(n_2448),
.Y(n_3292)
);

HB1xp67_ASAP7_75t_L g3293 ( 
.A(n_2753),
.Y(n_3293)
);

INVx4_ASAP7_75t_L g3294 ( 
.A(n_2660),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2701),
.B(n_2342),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2617),
.Y(n_3296)
);

INVx3_ASAP7_75t_L g3297 ( 
.A(n_2633),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_2617),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_2703),
.B(n_2332),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2619),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_2619),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_SL g3302 ( 
.A(n_2961),
.B(n_2425),
.Y(n_3302)
);

BUFx3_ASAP7_75t_L g3303 ( 
.A(n_2764),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_L g3304 ( 
.A1(n_2749),
.A2(n_2195),
.B1(n_2200),
.B2(n_2171),
.Y(n_3304)
);

NOR2xp33_ASAP7_75t_L g3305 ( 
.A(n_2699),
.B(n_2448),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_2624),
.Y(n_3306)
);

OAI22xp5_ASAP7_75t_L g3307 ( 
.A1(n_2968),
.A2(n_2350),
.B1(n_2375),
.B2(n_2371),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_2703),
.B(n_2332),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_2624),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_2629),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_2629),
.Y(n_3311)
);

AOI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_2756),
.A2(n_2284),
.B1(n_2171),
.B2(n_2527),
.Y(n_3312)
);

INVx5_ASAP7_75t_L g3313 ( 
.A(n_2660),
.Y(n_3313)
);

BUFx2_ASAP7_75t_L g3314 ( 
.A(n_2778),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2633),
.Y(n_3315)
);

INVx3_ASAP7_75t_L g3316 ( 
.A(n_2637),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2637),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_2536),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_SL g3319 ( 
.A(n_2961),
.B(n_2425),
.Y(n_3319)
);

INVx3_ASAP7_75t_L g3320 ( 
.A(n_2638),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_2536),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_2543),
.Y(n_3322)
);

NOR2x1p5_ASAP7_75t_L g3323 ( 
.A(n_2702),
.B(n_2363),
.Y(n_3323)
);

AND2x6_ASAP7_75t_L g3324 ( 
.A(n_2630),
.B(n_2543),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2704),
.B(n_2332),
.Y(n_3325)
);

BUFx2_ASAP7_75t_L g3326 ( 
.A(n_2546),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2638),
.Y(n_3327)
);

BUFx3_ASAP7_75t_L g3328 ( 
.A(n_2576),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_2643),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_2643),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_2650),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_2650),
.Y(n_3332)
);

INVx3_ASAP7_75t_L g3333 ( 
.A(n_2761),
.Y(n_3333)
);

OR2x2_ASAP7_75t_L g3334 ( 
.A(n_2712),
.B(n_2485),
.Y(n_3334)
);

INVx2_ASAP7_75t_SL g3335 ( 
.A(n_2589),
.Y(n_3335)
);

CKINVDCx16_ASAP7_75t_R g3336 ( 
.A(n_2565),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_2690),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_SL g3338 ( 
.A(n_2961),
.B(n_2425),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_2690),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2644),
.Y(n_3340)
);

BUFx4f_ASAP7_75t_L g3341 ( 
.A(n_2730),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_2704),
.B(n_2351),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_2644),
.Y(n_3343)
);

INVx5_ASAP7_75t_L g3344 ( 
.A(n_2660),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_2694),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_2968),
.A2(n_2350),
.B1(n_2375),
.B2(n_2371),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_2772),
.A2(n_2284),
.B1(n_2219),
.B2(n_2224),
.Y(n_3347)
);

NOR2xp33_ASAP7_75t_L g3348 ( 
.A(n_2621),
.B(n_2463),
.Y(n_3348)
);

AOI22xp33_ASAP7_75t_L g3349 ( 
.A1(n_2772),
.A2(n_2219),
.B1(n_2224),
.B2(n_2213),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_2708),
.B(n_2356),
.Y(n_3350)
);

OR2x2_ASAP7_75t_L g3351 ( 
.A(n_2719),
.B(n_2485),
.Y(n_3351)
);

INVx2_ASAP7_75t_SL g3352 ( 
.A(n_2589),
.Y(n_3352)
);

NOR2xp33_ASAP7_75t_L g3353 ( 
.A(n_2569),
.B(n_2463),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2645),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_2645),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2647),
.Y(n_3356)
);

AND2x4_ASAP7_75t_L g3357 ( 
.A(n_2835),
.B(n_2478),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_2647),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_2920),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_SL g3360 ( 
.A(n_2656),
.B(n_2425),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_2694),
.Y(n_3361)
);

AND2x6_ASAP7_75t_L g3362 ( 
.A(n_2591),
.B(n_2425),
.Y(n_3362)
);

NOR2xp33_ASAP7_75t_L g3363 ( 
.A(n_2578),
.B(n_2463),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_SL g3364 ( 
.A(n_2656),
.B(n_2429),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2920),
.Y(n_3365)
);

BUFx6f_ASAP7_75t_L g3366 ( 
.A(n_2716),
.Y(n_3366)
);

BUFx6f_ASAP7_75t_L g3367 ( 
.A(n_2716),
.Y(n_3367)
);

AOI22xp33_ASAP7_75t_L g3368 ( 
.A1(n_2784),
.A2(n_2224),
.B1(n_2226),
.B2(n_2219),
.Y(n_3368)
);

INVx2_ASAP7_75t_SL g3369 ( 
.A(n_2656),
.Y(n_3369)
);

AND2x6_ASAP7_75t_L g3370 ( 
.A(n_2591),
.B(n_2429),
.Y(n_3370)
);

OR2x2_ASAP7_75t_L g3371 ( 
.A(n_2532),
.B(n_2497),
.Y(n_3371)
);

AND2x6_ASAP7_75t_L g3372 ( 
.A(n_2591),
.B(n_2429),
.Y(n_3372)
);

AOI22xp5_ASAP7_75t_L g3373 ( 
.A1(n_2545),
.A2(n_2391),
.B1(n_2396),
.B2(n_2388),
.Y(n_3373)
);

BUFx6f_ASAP7_75t_L g3374 ( 
.A(n_2716),
.Y(n_3374)
);

HB1xp67_ASAP7_75t_L g3375 ( 
.A(n_2817),
.Y(n_3375)
);

HB1xp67_ASAP7_75t_L g3376 ( 
.A(n_2817),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_SL g3377 ( 
.A(n_2817),
.B(n_2429),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_2922),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_2922),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_2705),
.Y(n_3380)
);

BUFx6f_ASAP7_75t_L g3381 ( 
.A(n_2716),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_L g3382 ( 
.A(n_2628),
.B(n_2325),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_2708),
.B(n_2294),
.Y(n_3383)
);

OAI22xp33_ASAP7_75t_L g3384 ( 
.A1(n_2713),
.A2(n_2350),
.B1(n_2391),
.B2(n_2388),
.Y(n_3384)
);

INVx2_ASAP7_75t_L g3385 ( 
.A(n_2705),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_2706),
.Y(n_3386)
);

NAND2x1p5_ASAP7_75t_L g3387 ( 
.A(n_2867),
.B(n_2478),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_2706),
.Y(n_3388)
);

INVx4_ASAP7_75t_L g3389 ( 
.A(n_2716),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_2710),
.Y(n_3390)
);

NAND2xp33_ASAP7_75t_L g3391 ( 
.A(n_2741),
.B(n_2429),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_2652),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_2713),
.B(n_2295),
.Y(n_3393)
);

NAND3xp33_ASAP7_75t_L g3394 ( 
.A(n_2965),
.B(n_1684),
.C(n_1683),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_2652),
.Y(n_3395)
);

AND2x4_ASAP7_75t_L g3396 ( 
.A(n_2927),
.B(n_2478),
.Y(n_3396)
);

NOR2x1p5_ASAP7_75t_L g3397 ( 
.A(n_2721),
.B(n_2363),
.Y(n_3397)
);

NAND2xp33_ASAP7_75t_L g3398 ( 
.A(n_2741),
.B(n_2462),
.Y(n_3398)
);

OR2x2_ASAP7_75t_L g3399 ( 
.A(n_2635),
.B(n_2497),
.Y(n_3399)
);

BUFx2_ASAP7_75t_L g3400 ( 
.A(n_2546),
.Y(n_3400)
);

AND3x2_ASAP7_75t_L g3401 ( 
.A(n_2895),
.B(n_2467),
.C(n_2432),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_2710),
.Y(n_3402)
);

NAND2xp33_ASAP7_75t_L g3403 ( 
.A(n_2741),
.B(n_2462),
.Y(n_3403)
);

HB1xp67_ASAP7_75t_L g3404 ( 
.A(n_2818),
.Y(n_3404)
);

NAND2xp33_ASAP7_75t_SL g3405 ( 
.A(n_2800),
.B(n_2462),
.Y(n_3405)
);

BUFx3_ASAP7_75t_L g3406 ( 
.A(n_2576),
.Y(n_3406)
);

INVx3_ASAP7_75t_L g3407 ( 
.A(n_2761),
.Y(n_3407)
);

BUFx6f_ASAP7_75t_SL g3408 ( 
.A(n_2642),
.Y(n_3408)
);

NOR2xp33_ASAP7_75t_L g3409 ( 
.A(n_2715),
.B(n_2328),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2784),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_SL g3411 ( 
.A(n_2818),
.B(n_2462),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_2714),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_2766),
.B(n_2308),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_2766),
.B(n_2767),
.Y(n_3414)
);

INVx2_ASAP7_75t_SL g3415 ( 
.A(n_2571),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_2767),
.B(n_2339),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_SL g3417 ( 
.A(n_2818),
.B(n_2462),
.Y(n_3417)
);

XOR2xp5_ASAP7_75t_L g3418 ( 
.A(n_2782),
.B(n_1776),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_2714),
.Y(n_3419)
);

INVx2_ASAP7_75t_SL g3420 ( 
.A(n_2571),
.Y(n_3420)
);

BUFx6f_ASAP7_75t_L g3421 ( 
.A(n_2741),
.Y(n_3421)
);

INVxp67_ASAP7_75t_SL g3422 ( 
.A(n_2741),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_2768),
.B(n_2396),
.Y(n_3423)
);

AOI22xp33_ASAP7_75t_L g3424 ( 
.A1(n_2786),
.A2(n_2224),
.B1(n_2226),
.B2(n_2219),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_SL g3425 ( 
.A(n_2786),
.B(n_2397),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_2726),
.Y(n_3426)
);

INVx1_ASAP7_75t_SL g3427 ( 
.A(n_2707),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_2726),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_2787),
.B(n_2397),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_2727),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_2727),
.Y(n_3431)
);

NAND3xp33_ASAP7_75t_L g3432 ( 
.A(n_2927),
.B(n_1684),
.C(n_2365),
.Y(n_3432)
);

INVx4_ASAP7_75t_L g3433 ( 
.A(n_2765),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_2729),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_2729),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_2739),
.Y(n_3436)
);

INVx3_ASAP7_75t_L g3437 ( 
.A(n_2761),
.Y(n_3437)
);

INVxp33_ASAP7_75t_L g3438 ( 
.A(n_2856),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_2739),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_2533),
.Y(n_3440)
);

INVx3_ASAP7_75t_L g3441 ( 
.A(n_2763),
.Y(n_3441)
);

NAND2xp33_ASAP7_75t_L g3442 ( 
.A(n_2765),
.B(n_2461),
.Y(n_3442)
);

BUFx6f_ASAP7_75t_L g3443 ( 
.A(n_3222),
.Y(n_3443)
);

NOR2x1p5_ASAP7_75t_L g3444 ( 
.A(n_3038),
.B(n_2363),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_3219),
.B(n_2398),
.Y(n_3445)
);

NOR3xp33_ASAP7_75t_L g3446 ( 
.A(n_3020),
.B(n_2504),
.C(n_2476),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3331),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3331),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3231),
.Y(n_3449)
);

NAND2xp33_ASAP7_75t_L g3450 ( 
.A(n_3276),
.B(n_2470),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3231),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3036),
.B(n_2768),
.Y(n_3452)
);

INVx2_ASAP7_75t_L g3453 ( 
.A(n_3239),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3035),
.B(n_2783),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_2984),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_SL g3456 ( 
.A(n_2994),
.B(n_2470),
.Y(n_3456)
);

INVx2_ASAP7_75t_L g3457 ( 
.A(n_3239),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3109),
.B(n_3052),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_2984),
.Y(n_3459)
);

INVxp33_ASAP7_75t_L g3460 ( 
.A(n_3043),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3245),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3097),
.B(n_2783),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3245),
.Y(n_3463)
);

INVx3_ASAP7_75t_L g3464 ( 
.A(n_3243),
.Y(n_3464)
);

BUFx6f_ASAP7_75t_SL g3465 ( 
.A(n_2989),
.Y(n_3465)
);

AND2x6_ASAP7_75t_SL g3466 ( 
.A(n_3382),
.B(n_2483),
.Y(n_3466)
);

CKINVDCx5p33_ASAP7_75t_R g3467 ( 
.A(n_3086),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_2986),
.B(n_2788),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_SL g3469 ( 
.A(n_2994),
.B(n_2471),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_2995),
.B(n_2788),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_2988),
.Y(n_3471)
);

AND2x2_ASAP7_75t_L g3472 ( 
.A(n_3219),
.B(n_2398),
.Y(n_3472)
);

BUFx6f_ASAP7_75t_SL g3473 ( 
.A(n_2989),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_SL g3474 ( 
.A(n_3025),
.B(n_2471),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_3287),
.B(n_2791),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3292),
.B(n_2789),
.Y(n_3476)
);

NOR2xp33_ASAP7_75t_L g3477 ( 
.A(n_3043),
.B(n_2461),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3063),
.B(n_2789),
.Y(n_3478)
);

NOR3xp33_ASAP7_75t_L g3479 ( 
.A(n_3160),
.B(n_2476),
.C(n_2482),
.Y(n_3479)
);

OR2x2_ASAP7_75t_L g3480 ( 
.A(n_3115),
.B(n_2530),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_3247),
.B(n_2400),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3224),
.B(n_2401),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_3254),
.Y(n_3483)
);

NOR2xp33_ASAP7_75t_L g3484 ( 
.A(n_3022),
.B(n_2400),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_2988),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_SL g3486 ( 
.A(n_3025),
.B(n_2471),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3063),
.B(n_2794),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3265),
.B(n_3161),
.Y(n_3488)
);

NAND2xp33_ASAP7_75t_L g3489 ( 
.A(n_3276),
.B(n_2471),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3161),
.B(n_3163),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3254),
.Y(n_3491)
);

INVxp33_ASAP7_75t_L g3492 ( 
.A(n_3086),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3041),
.Y(n_3493)
);

NOR2xp33_ASAP7_75t_L g3494 ( 
.A(n_3022),
.B(n_3079),
.Y(n_3494)
);

NOR3xp33_ASAP7_75t_L g3495 ( 
.A(n_3062),
.B(n_2482),
.C(n_2494),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3041),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3049),
.Y(n_3497)
);

AND2x2_ASAP7_75t_L g3498 ( 
.A(n_3224),
.B(n_2401),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3163),
.B(n_2794),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3342),
.B(n_2662),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_SL g3501 ( 
.A(n_3185),
.B(n_2471),
.Y(n_3501)
);

NOR2xp67_ASAP7_75t_SL g3502 ( 
.A(n_2982),
.B(n_2350),
.Y(n_3502)
);

BUFx6f_ASAP7_75t_L g3503 ( 
.A(n_3222),
.Y(n_3503)
);

NOR2xp33_ASAP7_75t_L g3504 ( 
.A(n_3068),
.B(n_2400),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3350),
.B(n_2662),
.Y(n_3505)
);

NOR2xp33_ASAP7_75t_L g3506 ( 
.A(n_3076),
.B(n_3140),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3262),
.Y(n_3507)
);

BUFx6f_ASAP7_75t_L g3508 ( 
.A(n_3222),
.Y(n_3508)
);

NAND2xp33_ASAP7_75t_L g3509 ( 
.A(n_3276),
.B(n_2473),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3132),
.B(n_2664),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_2996),
.B(n_2404),
.Y(n_3511)
);

INVx2_ASAP7_75t_L g3512 ( 
.A(n_3262),
.Y(n_3512)
);

NAND2xp33_ASAP7_75t_L g3513 ( 
.A(n_3276),
.B(n_2473),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3266),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3266),
.Y(n_3515)
);

AOI221xp5_ASAP7_75t_L g3516 ( 
.A1(n_3193),
.A2(n_3272),
.B1(n_3123),
.B2(n_868),
.C(n_869),
.Y(n_3516)
);

AND2x2_ASAP7_75t_L g3517 ( 
.A(n_2996),
.B(n_3058),
.Y(n_3517)
);

BUFx5_ASAP7_75t_L g3518 ( 
.A(n_3324),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_3334),
.B(n_2465),
.Y(n_3519)
);

OA21x2_ASAP7_75t_L g3520 ( 
.A1(n_3440),
.A2(n_2547),
.B(n_2553),
.Y(n_3520)
);

NOR2xp33_ASAP7_75t_SL g3521 ( 
.A(n_3119),
.B(n_2168),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3058),
.B(n_2404),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3049),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_3132),
.B(n_2664),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3055),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3305),
.B(n_2666),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_SL g3527 ( 
.A(n_3187),
.B(n_2473),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3055),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3278),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3056),
.Y(n_3530)
);

INVxp67_ASAP7_75t_L g3531 ( 
.A(n_3115),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_SL g3532 ( 
.A(n_3203),
.B(n_2473),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3383),
.B(n_2666),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3056),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_SL g3535 ( 
.A(n_3174),
.B(n_3183),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3278),
.Y(n_3536)
);

INVx2_ASAP7_75t_SL g3537 ( 
.A(n_3032),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3289),
.Y(n_3538)
);

AND2x2_ASAP7_75t_L g3539 ( 
.A(n_3235),
.B(n_2412),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_SL g3540 ( 
.A(n_3288),
.B(n_2473),
.Y(n_3540)
);

INVxp33_ASAP7_75t_L g3541 ( 
.A(n_3209),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3059),
.Y(n_3542)
);

BUFx6f_ASAP7_75t_SL g3543 ( 
.A(n_3032),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3059),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3393),
.B(n_2667),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3289),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3413),
.B(n_2667),
.Y(n_3547)
);

NOR2xp67_ASAP7_75t_L g3548 ( 
.A(n_3394),
.B(n_2482),
.Y(n_3548)
);

NAND2xp33_ASAP7_75t_L g3549 ( 
.A(n_3276),
.B(n_2477),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3077),
.Y(n_3550)
);

INVx1_ASAP7_75t_SL g3551 ( 
.A(n_2998),
.Y(n_3551)
);

NOR2xp33_ASAP7_75t_L g3552 ( 
.A(n_3334),
.B(n_2465),
.Y(n_3552)
);

NOR3xp33_ASAP7_75t_L g3553 ( 
.A(n_3432),
.B(n_2484),
.C(n_2483),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3416),
.B(n_2671),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3066),
.B(n_2671),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3298),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3077),
.Y(n_3557)
);

INVx2_ASAP7_75t_L g3558 ( 
.A(n_3298),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3301),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3066),
.B(n_2672),
.Y(n_3560)
);

INVxp67_ASAP7_75t_L g3561 ( 
.A(n_3235),
.Y(n_3561)
);

INVxp67_ASAP7_75t_L g3562 ( 
.A(n_3293),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_3301),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_2990),
.B(n_2407),
.Y(n_3564)
);

NOR2xp33_ASAP7_75t_L g3565 ( 
.A(n_3027),
.B(n_2423),
.Y(n_3565)
);

NAND2xp33_ASAP7_75t_L g3566 ( 
.A(n_3276),
.B(n_2477),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3050),
.B(n_2672),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3050),
.B(n_2722),
.Y(n_3568)
);

NAND2xp33_ASAP7_75t_L g3569 ( 
.A(n_3092),
.B(n_2477),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3103),
.B(n_2723),
.Y(n_3570)
);

OR2x2_ASAP7_75t_SL g3571 ( 
.A(n_3336),
.B(n_2477),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3082),
.Y(n_3572)
);

BUFx5_ASAP7_75t_L g3573 ( 
.A(n_3324),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_L g3574 ( 
.A(n_3423),
.B(n_2438),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3306),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3255),
.B(n_2412),
.Y(n_3576)
);

NOR2xp33_ASAP7_75t_L g3577 ( 
.A(n_2978),
.B(n_2449),
.Y(n_3577)
);

NOR3xp33_ASAP7_75t_L g3578 ( 
.A(n_3409),
.B(n_2488),
.C(n_2484),
.Y(n_3578)
);

INVx2_ASAP7_75t_SL g3579 ( 
.A(n_3065),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3306),
.Y(n_3580)
);

NOR2xp33_ASAP7_75t_L g3581 ( 
.A(n_2978),
.B(n_2434),
.Y(n_3581)
);

NOR2xp33_ASAP7_75t_L g3582 ( 
.A(n_3103),
.B(n_2434),
.Y(n_3582)
);

NOR2xp33_ASAP7_75t_L g3583 ( 
.A(n_3117),
.B(n_2456),
.Y(n_3583)
);

AND3x4_ASAP7_75t_L g3584 ( 
.A(n_3130),
.B(n_2468),
.C(n_2500),
.Y(n_3584)
);

INVx2_ASAP7_75t_SL g3585 ( 
.A(n_3083),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3117),
.B(n_2724),
.Y(n_3586)
);

OR2x2_ASAP7_75t_L g3587 ( 
.A(n_3069),
.B(n_2530),
.Y(n_3587)
);

INVxp33_ASAP7_75t_L g3588 ( 
.A(n_3209),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_L g3589 ( 
.A(n_3124),
.B(n_2456),
.Y(n_3589)
);

INVx2_ASAP7_75t_SL g3590 ( 
.A(n_3087),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3082),
.Y(n_3591)
);

INVx2_ASAP7_75t_SL g3592 ( 
.A(n_3351),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3084),
.Y(n_3593)
);

NOR2xp33_ASAP7_75t_L g3594 ( 
.A(n_3124),
.B(n_2459),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3150),
.B(n_2728),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3150),
.B(n_3127),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3084),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3255),
.B(n_2733),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3139),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3139),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3148),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3148),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3090),
.B(n_2742),
.Y(n_3603)
);

AOI221xp5_ASAP7_75t_L g3604 ( 
.A1(n_3218),
.A2(n_868),
.B1(n_869),
.B2(n_866),
.C(n_859),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3108),
.B(n_2745),
.Y(n_3605)
);

INVx8_ASAP7_75t_L g3606 ( 
.A(n_3060),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3238),
.B(n_2748),
.Y(n_3607)
);

INVx5_ASAP7_75t_L g3608 ( 
.A(n_2973),
.Y(n_3608)
);

INVxp67_ASAP7_75t_SL g3609 ( 
.A(n_2973),
.Y(n_3609)
);

BUFx6f_ASAP7_75t_L g3610 ( 
.A(n_3222),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3414),
.B(n_2750),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3162),
.Y(n_3612)
);

BUFx2_ASAP7_75t_L g3613 ( 
.A(n_3130),
.Y(n_3613)
);

INVxp67_ASAP7_75t_SL g3614 ( 
.A(n_2973),
.Y(n_3614)
);

NOR3xp33_ASAP7_75t_L g3615 ( 
.A(n_3353),
.B(n_2489),
.C(n_2488),
.Y(n_3615)
);

BUFx6f_ASAP7_75t_SL g3616 ( 
.A(n_3019),
.Y(n_3616)
);

NAND3xp33_ASAP7_75t_L g3617 ( 
.A(n_3159),
.B(n_2505),
.C(n_2480),
.Y(n_3617)
);

INVx2_ASAP7_75t_L g3618 ( 
.A(n_3037),
.Y(n_3618)
);

NAND3xp33_ASAP7_75t_L g3619 ( 
.A(n_3373),
.B(n_2505),
.C(n_2466),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_3037),
.Y(n_3620)
);

INVx6_ASAP7_75t_L g3621 ( 
.A(n_3017),
.Y(n_3621)
);

HB1xp67_ASAP7_75t_L g3622 ( 
.A(n_3314),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_2972),
.B(n_2751),
.Y(n_3623)
);

AOI22xp5_ASAP7_75t_L g3624 ( 
.A1(n_3363),
.A2(n_2717),
.B1(n_2926),
.B2(n_2754),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3039),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3165),
.B(n_2755),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3288),
.B(n_2771),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3039),
.Y(n_3628)
);

OR2x6_ASAP7_75t_L g3629 ( 
.A(n_3093),
.B(n_2477),
.Y(n_3629)
);

BUFx5_ASAP7_75t_L g3630 ( 
.A(n_3324),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3044),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3335),
.B(n_2776),
.Y(n_3632)
);

NOR2xp33_ASAP7_75t_L g3633 ( 
.A(n_3438),
.B(n_3236),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3335),
.B(n_2777),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3162),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3352),
.B(n_3369),
.Y(n_3636)
);

OR2x2_ASAP7_75t_SL g3637 ( 
.A(n_3205),
.B(n_2481),
.Y(n_3637)
);

INVx2_ASAP7_75t_SL g3638 ( 
.A(n_3351),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_SL g3639 ( 
.A(n_3352),
.B(n_2481),
.Y(n_3639)
);

INVx2_ASAP7_75t_L g3640 ( 
.A(n_3044),
.Y(n_3640)
);

INVxp67_ASAP7_75t_L g3641 ( 
.A(n_3314),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3369),
.B(n_2780),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_SL g3643 ( 
.A(n_3220),
.B(n_2481),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3048),
.Y(n_3644)
);

BUFx5_ASAP7_75t_L g3645 ( 
.A(n_3324),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3195),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3048),
.Y(n_3647)
);

AND2x2_ASAP7_75t_L g3648 ( 
.A(n_3134),
.B(n_2459),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3195),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3415),
.B(n_2781),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_L g3651 ( 
.A(n_3438),
.B(n_2369),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3057),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3199),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_SL g3654 ( 
.A(n_3220),
.B(n_2481),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3199),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3057),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3072),
.Y(n_3657)
);

NOR2xp33_ASAP7_75t_L g3658 ( 
.A(n_3236),
.B(n_2369),
.Y(n_3658)
);

NOR2xp33_ASAP7_75t_L g3659 ( 
.A(n_3281),
.B(n_3399),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3207),
.Y(n_3660)
);

NOR2xp67_ASAP7_75t_L g3661 ( 
.A(n_3116),
.B(n_2168),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3415),
.B(n_2819),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3420),
.B(n_2821),
.Y(n_3663)
);

NOR2xp33_ASAP7_75t_L g3664 ( 
.A(n_3281),
.B(n_2370),
.Y(n_3664)
);

NAND3xp33_ASAP7_75t_L g3665 ( 
.A(n_3348),
.B(n_2364),
.C(n_2346),
.Y(n_3665)
);

NAND3xp33_ASAP7_75t_L g3666 ( 
.A(n_3399),
.B(n_2290),
.C(n_2228),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3207),
.Y(n_3667)
);

INVxp67_ASAP7_75t_L g3668 ( 
.A(n_3375),
.Y(n_3668)
);

NOR3xp33_ASAP7_75t_L g3669 ( 
.A(n_3360),
.B(n_2490),
.C(n_2489),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3296),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3296),
.Y(n_3671)
);

BUFx5_ASAP7_75t_L g3672 ( 
.A(n_3324),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3300),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3420),
.B(n_2823),
.Y(n_3674)
);

NOR3xp33_ASAP7_75t_L g3675 ( 
.A(n_3364),
.B(n_2495),
.C(n_2490),
.Y(n_3675)
);

BUFx3_ASAP7_75t_L g3676 ( 
.A(n_3145),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_SL g3677 ( 
.A(n_3220),
.B(n_2481),
.Y(n_3677)
);

NOR3xp33_ASAP7_75t_L g3678 ( 
.A(n_3377),
.B(n_2502),
.C(n_2495),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3014),
.B(n_3026),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3300),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3028),
.B(n_2830),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3309),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3155),
.B(n_2831),
.Y(n_3683)
);

NOR3xp33_ASAP7_75t_L g3684 ( 
.A(n_3411),
.B(n_2502),
.C(n_2501),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_SL g3685 ( 
.A(n_3271),
.B(n_2427),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3283),
.B(n_2832),
.Y(n_3686)
);

OR2x2_ASAP7_75t_L g3687 ( 
.A(n_3371),
.B(n_2506),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3309),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3073),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_2974),
.B(n_2833),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_2975),
.B(n_2834),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_2977),
.B(n_2840),
.Y(n_3692)
);

INVx2_ASAP7_75t_SL g3693 ( 
.A(n_3371),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3310),
.Y(n_3694)
);

NOR2xp33_ASAP7_75t_L g3695 ( 
.A(n_3134),
.B(n_2370),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_2987),
.B(n_2841),
.Y(n_3696)
);

INVxp67_ASAP7_75t_SL g3697 ( 
.A(n_2973),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_SL g3698 ( 
.A(n_3271),
.B(n_2427),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3002),
.B(n_2842),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3003),
.B(n_2928),
.Y(n_3700)
);

NOR2xp33_ASAP7_75t_L g3701 ( 
.A(n_3136),
.B(n_2382),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3310),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3311),
.Y(n_3703)
);

BUFx2_ASAP7_75t_R g3704 ( 
.A(n_3214),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_SL g3705 ( 
.A(n_3271),
.B(n_2445),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3006),
.B(n_2928),
.Y(n_3706)
);

NOR2xp33_ASAP7_75t_L g3707 ( 
.A(n_3136),
.B(n_2382),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3073),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3007),
.B(n_3018),
.Y(n_3709)
);

BUFx6f_ASAP7_75t_L g3710 ( 
.A(n_3222),
.Y(n_3710)
);

AND2x2_ASAP7_75t_L g3711 ( 
.A(n_3181),
.B(n_2475),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3024),
.B(n_2929),
.Y(n_3712)
);

INVxp67_ASAP7_75t_L g3713 ( 
.A(n_3376),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_SL g3714 ( 
.A(n_3357),
.B(n_2445),
.Y(n_3714)
);

NOR2xp33_ASAP7_75t_L g3715 ( 
.A(n_3181),
.B(n_2385),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3208),
.B(n_2929),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3075),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_SL g3718 ( 
.A(n_3357),
.B(n_2385),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3208),
.B(n_2930),
.Y(n_3719)
);

AND2x2_ASAP7_75t_L g3720 ( 
.A(n_3269),
.B(n_2475),
.Y(n_3720)
);

INVx1_ASAP7_75t_SL g3721 ( 
.A(n_3145),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3012),
.B(n_2930),
.Y(n_3722)
);

INVx8_ASAP7_75t_L g3723 ( 
.A(n_3060),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3075),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_SL g3725 ( 
.A(n_3357),
.B(n_2390),
.Y(n_3725)
);

NOR2xp33_ASAP7_75t_SL g3726 ( 
.A(n_3116),
.B(n_2228),
.Y(n_3726)
);

INVx1_ASAP7_75t_SL g3727 ( 
.A(n_3098),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3078),
.Y(n_3728)
);

NOR2xp33_ASAP7_75t_L g3729 ( 
.A(n_3269),
.B(n_2390),
.Y(n_3729)
);

INVxp33_ASAP7_75t_L g3730 ( 
.A(n_3418),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3078),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3311),
.Y(n_3732)
);

INVx2_ASAP7_75t_L g3733 ( 
.A(n_3095),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3340),
.Y(n_3734)
);

NAND2xp33_ASAP7_75t_L g3735 ( 
.A(n_3092),
.B(n_2730),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3410),
.B(n_2931),
.Y(n_3736)
);

INVx3_ASAP7_75t_L g3737 ( 
.A(n_3243),
.Y(n_3737)
);

NOR2xp33_ASAP7_75t_L g3738 ( 
.A(n_3282),
.B(n_2395),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3340),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3095),
.Y(n_3740)
);

NOR2xp33_ASAP7_75t_L g3741 ( 
.A(n_3282),
.B(n_2395),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3343),
.Y(n_3742)
);

BUFx6f_ASAP7_75t_L g3743 ( 
.A(n_3229),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3099),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_SL g3745 ( 
.A(n_2983),
.B(n_2399),
.Y(n_3745)
);

OA21x2_ASAP7_75t_L g3746 ( 
.A1(n_3440),
.A2(n_2547),
.B(n_2553),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3343),
.Y(n_3747)
);

NOR2xp33_ASAP7_75t_L g3748 ( 
.A(n_3284),
.B(n_2399),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3354),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3099),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_2983),
.B(n_2934),
.Y(n_3751)
);

NOR2xp33_ASAP7_75t_L g3752 ( 
.A(n_3284),
.B(n_2435),
.Y(n_3752)
);

INVx3_ASAP7_75t_L g3753 ( 
.A(n_3243),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_2983),
.B(n_2934),
.Y(n_3754)
);

NOR2xp33_ASAP7_75t_L g3755 ( 
.A(n_3303),
.B(n_2435),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3260),
.B(n_2936),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3354),
.B(n_2936),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3106),
.Y(n_3758)
);

AO221x1_ASAP7_75t_L g3759 ( 
.A1(n_3040),
.A2(n_2487),
.B1(n_2496),
.B2(n_2498),
.C(n_2491),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3355),
.B(n_2937),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3355),
.B(n_2937),
.Y(n_3761)
);

INVx2_ASAP7_75t_SL g3762 ( 
.A(n_3397),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3356),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3356),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3358),
.B(n_2938),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3358),
.Y(n_3766)
);

BUFx5_ASAP7_75t_L g3767 ( 
.A(n_3324),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3030),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_2979),
.B(n_2938),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3106),
.Y(n_3770)
);

AOI22xp5_ASAP7_75t_L g3771 ( 
.A1(n_3171),
.A2(n_3404),
.B1(n_3319),
.B2(n_3338),
.Y(n_3771)
);

NOR2xp33_ASAP7_75t_L g3772 ( 
.A(n_3303),
.B(n_2437),
.Y(n_3772)
);

BUFx6f_ASAP7_75t_L g3773 ( 
.A(n_3229),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3392),
.B(n_2939),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3395),
.B(n_2939),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_SL g3776 ( 
.A(n_3307),
.B(n_2437),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3033),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_3111),
.Y(n_3778)
);

NOR2xp33_ASAP7_75t_L g3779 ( 
.A(n_3425),
.B(n_2439),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3019),
.B(n_2430),
.Y(n_3780)
);

INVxp67_ASAP7_75t_L g3781 ( 
.A(n_3274),
.Y(n_3781)
);

INVxp67_ASAP7_75t_SL g3782 ( 
.A(n_2973),
.Y(n_3782)
);

NOR2xp67_ASAP7_75t_L g3783 ( 
.A(n_3176),
.B(n_2290),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3429),
.B(n_2942),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3346),
.B(n_2982),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_SL g3786 ( 
.A(n_2982),
.B(n_2439),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3051),
.Y(n_3787)
);

NOR2xp33_ASAP7_75t_L g3788 ( 
.A(n_3171),
.B(n_2457),
.Y(n_3788)
);

BUFx6f_ASAP7_75t_L g3789 ( 
.A(n_3229),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3121),
.B(n_2942),
.Y(n_3790)
);

BUFx3_ASAP7_75t_L g3791 ( 
.A(n_3129),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3088),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3111),
.Y(n_3793)
);

NAND2x1_ASAP7_75t_L g3794 ( 
.A(n_3001),
.B(n_2968),
.Y(n_3794)
);

NOR2xp33_ASAP7_75t_L g3795 ( 
.A(n_3171),
.B(n_2457),
.Y(n_3795)
);

A2O1A1Ixp33_ASAP7_75t_L g3796 ( 
.A1(n_3125),
.A2(n_2943),
.B(n_2698),
.C(n_2962),
.Y(n_3796)
);

NOR2xp33_ASAP7_75t_L g3797 ( 
.A(n_3427),
.B(n_2472),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3112),
.Y(n_3798)
);

INVxp67_ASAP7_75t_L g3799 ( 
.A(n_3417),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_L g3800 ( 
.A(n_3154),
.B(n_2472),
.Y(n_3800)
);

NOR2xp67_ASAP7_75t_SL g3801 ( 
.A(n_2982),
.B(n_2379),
.Y(n_3801)
);

HB1xp67_ASAP7_75t_L g3802 ( 
.A(n_2997),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_SL g3803 ( 
.A(n_2982),
.B(n_2421),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_SL g3804 ( 
.A(n_3074),
.B(n_2428),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3177),
.B(n_2737),
.Y(n_3805)
);

NOR2xp33_ASAP7_75t_L g3806 ( 
.A(n_3228),
.B(n_2365),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3246),
.B(n_2747),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3252),
.B(n_2747),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3112),
.Y(n_3809)
);

BUFx6f_ASAP7_75t_L g3810 ( 
.A(n_3229),
.Y(n_3810)
);

AND2x2_ASAP7_75t_SL g3811 ( 
.A(n_3202),
.B(n_2971),
.Y(n_3811)
);

NOR2xp33_ASAP7_75t_SL g3812 ( 
.A(n_3176),
.B(n_2409),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3100),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3253),
.B(n_2752),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_SL g3815 ( 
.A(n_3074),
.B(n_2443),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3133),
.Y(n_3816)
);

AOI22xp5_ASAP7_75t_L g3817 ( 
.A1(n_3302),
.A2(n_2946),
.B1(n_2960),
.B2(n_2879),
.Y(n_3817)
);

NOR2xp33_ASAP7_75t_L g3818 ( 
.A(n_3256),
.B(n_2366),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3101),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_SL g3820 ( 
.A(n_3074),
.B(n_2444),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_SL g3821 ( 
.A(n_3074),
.B(n_2450),
.Y(n_3821)
);

INVx3_ASAP7_75t_L g3822 ( 
.A(n_3243),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3104),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3091),
.B(n_2752),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_SL g3825 ( 
.A(n_3074),
.B(n_3141),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_SL g3826 ( 
.A(n_3141),
.B(n_2454),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3133),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3113),
.Y(n_3828)
);

NOR2xp33_ASAP7_75t_L g3829 ( 
.A(n_3053),
.B(n_2366),
.Y(n_3829)
);

NOR2xp67_ASAP7_75t_L g3830 ( 
.A(n_3217),
.B(n_2409),
.Y(n_3830)
);

BUFx3_ASAP7_75t_L g3831 ( 
.A(n_3129),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3323),
.B(n_2571),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3384),
.B(n_2752),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3118),
.Y(n_3834)
);

NOR2xp67_ASAP7_75t_L g3835 ( 
.A(n_3217),
.B(n_2479),
.Y(n_3835)
);

INVx4_ASAP7_75t_L g3836 ( 
.A(n_3229),
.Y(n_3836)
);

BUFx6f_ASAP7_75t_L g3837 ( 
.A(n_3250),
.Y(n_3837)
);

NAND2x1p5_ASAP7_75t_L g3838 ( 
.A(n_3608),
.B(n_3141),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_SL g3839 ( 
.A(n_3506),
.B(n_2508),
.Y(n_3839)
);

NAND2xp33_ASAP7_75t_L g3840 ( 
.A(n_3458),
.B(n_3092),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3455),
.Y(n_3841)
);

AND2x6_ASAP7_75t_SL g3842 ( 
.A(n_3565),
.B(n_2511),
.Y(n_3842)
);

INVx8_ASAP7_75t_L g3843 ( 
.A(n_3606),
.Y(n_3843)
);

AND2x2_ASAP7_75t_SL g3844 ( 
.A(n_3506),
.B(n_3216),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3462),
.B(n_2976),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3449),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3459),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3494),
.B(n_2976),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3451),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3453),
.Y(n_3850)
);

BUFx12f_ASAP7_75t_L g3851 ( 
.A(n_3579),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3471),
.Y(n_3852)
);

NAND2x1p5_ASAP7_75t_L g3853 ( 
.A(n_3608),
.B(n_3141),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3457),
.Y(n_3854)
);

NOR2xp33_ASAP7_75t_L g3855 ( 
.A(n_3494),
.B(n_3504),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3454),
.B(n_2992),
.Y(n_3856)
);

NOR2xp33_ASAP7_75t_L g3857 ( 
.A(n_3504),
.B(n_3484),
.Y(n_3857)
);

BUFx3_ASAP7_75t_L g3858 ( 
.A(n_3606),
.Y(n_3858)
);

NOR2x1p5_ASAP7_75t_L g3859 ( 
.A(n_3666),
.B(n_2175),
.Y(n_3859)
);

BUFx3_ASAP7_75t_L g3860 ( 
.A(n_3606),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3452),
.B(n_2992),
.Y(n_3861)
);

OAI22xp5_ASAP7_75t_L g3862 ( 
.A1(n_3533),
.A2(n_3206),
.B1(n_3152),
.B2(n_3093),
.Y(n_3862)
);

AOI22xp33_ASAP7_75t_L g3863 ( 
.A1(n_3516),
.A2(n_3067),
.B1(n_3168),
.B2(n_3326),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3461),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3468),
.B(n_2993),
.Y(n_3865)
);

NOR3xp33_ASAP7_75t_L g3866 ( 
.A(n_3484),
.B(n_2236),
.C(n_2512),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3485),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3463),
.Y(n_3868)
);

AND2x4_ASAP7_75t_L g3869 ( 
.A(n_3762),
.B(n_3017),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3493),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3521),
.B(n_2508),
.Y(n_3871)
);

OR2x6_ASAP7_75t_L g3872 ( 
.A(n_3723),
.B(n_3093),
.Y(n_3872)
);

NOR2xp33_ASAP7_75t_L g3873 ( 
.A(n_3574),
.B(n_2405),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3483),
.Y(n_3874)
);

BUFx3_ASAP7_75t_L g3875 ( 
.A(n_3723),
.Y(n_3875)
);

INVx2_ASAP7_75t_SL g3876 ( 
.A(n_3585),
.Y(n_3876)
);

INVxp67_ASAP7_75t_L g3877 ( 
.A(n_3587),
.Y(n_3877)
);

OR2x2_ASAP7_75t_L g3878 ( 
.A(n_3480),
.B(n_2468),
.Y(n_3878)
);

NOR2xp33_ASAP7_75t_L g3879 ( 
.A(n_3574),
.B(n_1777),
.Y(n_3879)
);

NOR2xp33_ASAP7_75t_L g3880 ( 
.A(n_3460),
.B(n_1777),
.Y(n_3880)
);

NOR2xp33_ASAP7_75t_L g3881 ( 
.A(n_3581),
.B(n_3577),
.Y(n_3881)
);

AO22x1_ASAP7_75t_L g3882 ( 
.A1(n_3481),
.A2(n_2359),
.B1(n_2924),
.B2(n_2612),
.Y(n_3882)
);

INVx2_ASAP7_75t_L g3883 ( 
.A(n_3491),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_SL g3884 ( 
.A(n_3477),
.B(n_2508),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3539),
.B(n_3168),
.Y(n_3885)
);

AOI22xp5_ASAP7_75t_L g3886 ( 
.A1(n_3577),
.A2(n_3418),
.B1(n_2525),
.B2(n_2523),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3470),
.B(n_2993),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3496),
.Y(n_3888)
);

NOR2xp33_ASAP7_75t_L g3889 ( 
.A(n_3581),
.B(n_1782),
.Y(n_3889)
);

NOR2xp33_ASAP7_75t_SL g3890 ( 
.A(n_3704),
.B(n_2479),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3507),
.Y(n_3891)
);

INVx2_ASAP7_75t_SL g3892 ( 
.A(n_3590),
.Y(n_3892)
);

BUFx2_ASAP7_75t_L g3893 ( 
.A(n_3613),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_L g3894 ( 
.A(n_3500),
.B(n_3505),
.Y(n_3894)
);

OAI22xp5_ASAP7_75t_SL g3895 ( 
.A1(n_3730),
.A2(n_3242),
.B1(n_3000),
.B2(n_2413),
.Y(n_3895)
);

AOI22xp33_ASAP7_75t_L g3896 ( 
.A1(n_3516),
.A2(n_3067),
.B1(n_3168),
.B2(n_3326),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_3517),
.B(n_2579),
.Y(n_3897)
);

A2O1A1Ixp33_ASAP7_75t_L g3898 ( 
.A1(n_3788),
.A2(n_3795),
.B(n_3800),
.C(n_3779),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_3545),
.B(n_2579),
.Y(n_3899)
);

AOI22xp33_ASAP7_75t_L g3900 ( 
.A1(n_3446),
.A2(n_3067),
.B1(n_3168),
.B2(n_3400),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3547),
.B(n_2579),
.Y(n_3901)
);

AOI22xp5_ASAP7_75t_L g3902 ( 
.A1(n_3565),
.A2(n_2525),
.B1(n_2523),
.B2(n_2511),
.Y(n_3902)
);

AND2x4_ASAP7_75t_L g3903 ( 
.A(n_3791),
.B(n_3017),
.Y(n_3903)
);

AOI22xp5_ASAP7_75t_L g3904 ( 
.A1(n_3726),
.A2(n_1782),
.B1(n_1811),
.B2(n_1799),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3497),
.Y(n_3905)
);

OR2x6_ASAP7_75t_L g3906 ( 
.A(n_3723),
.B(n_3093),
.Y(n_3906)
);

O2A1O1Ixp33_ASAP7_75t_L g3907 ( 
.A1(n_3446),
.A2(n_2469),
.B(n_2501),
.C(n_2500),
.Y(n_3907)
);

INVx2_ASAP7_75t_SL g3908 ( 
.A(n_3831),
.Y(n_3908)
);

INVx2_ASAP7_75t_SL g3909 ( 
.A(n_3551),
.Y(n_3909)
);

NOR2xp33_ASAP7_75t_L g3910 ( 
.A(n_3477),
.B(n_1799),
.Y(n_3910)
);

AOI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3812),
.A2(n_1811),
.B1(n_1821),
.B2(n_1814),
.Y(n_3911)
);

NAND3xp33_ASAP7_75t_L g3912 ( 
.A(n_3495),
.B(n_3479),
.C(n_3615),
.Y(n_3912)
);

CKINVDCx5p33_ASAP7_75t_R g3913 ( 
.A(n_3467),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3512),
.Y(n_3914)
);

INVx2_ASAP7_75t_L g3915 ( 
.A(n_3514),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3511),
.B(n_3270),
.Y(n_3916)
);

OAI22xp33_ASAP7_75t_L g3917 ( 
.A1(n_3687),
.A2(n_2496),
.B1(n_2487),
.B2(n_2508),
.Y(n_3917)
);

INVx2_ASAP7_75t_L g3918 ( 
.A(n_3515),
.Y(n_3918)
);

AOI22xp33_ASAP7_75t_L g3919 ( 
.A1(n_3788),
.A2(n_3400),
.B1(n_2730),
.B2(n_3396),
.Y(n_3919)
);

O2A1O1Ixp5_ASAP7_75t_L g3920 ( 
.A1(n_3535),
.A2(n_3776),
.B(n_3501),
.C(n_3532),
.Y(n_3920)
);

INVx3_ASAP7_75t_L g3921 ( 
.A(n_3621),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3529),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3554),
.B(n_2822),
.Y(n_3923)
);

O2A1O1Ixp33_ASAP7_75t_L g3924 ( 
.A1(n_3479),
.A2(n_2469),
.B(n_2503),
.C(n_2521),
.Y(n_3924)
);

NOR2xp33_ASAP7_75t_L g3925 ( 
.A(n_3797),
.B(n_1814),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_SL g3926 ( 
.A(n_3481),
.B(n_2508),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3523),
.Y(n_3927)
);

INVx4_ASAP7_75t_L g3928 ( 
.A(n_3608),
.Y(n_3928)
);

A2O1A1Ixp33_ASAP7_75t_L g3929 ( 
.A1(n_3795),
.A2(n_3004),
.B(n_3405),
.C(n_3341),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_3536),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3482),
.B(n_2822),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_3538),
.Y(n_3932)
);

NAND2x1p5_ASAP7_75t_L g3933 ( 
.A(n_3608),
.B(n_3141),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3546),
.Y(n_3934)
);

AOI22xp33_ASAP7_75t_L g3935 ( 
.A1(n_3495),
.A2(n_3396),
.B1(n_2657),
.B2(n_2546),
.Y(n_3935)
);

INVx2_ASAP7_75t_SL g3936 ( 
.A(n_3537),
.Y(n_3936)
);

OAI22xp5_ASAP7_75t_SL g3937 ( 
.A1(n_3584),
.A2(n_3242),
.B1(n_3000),
.B2(n_1705),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_SL g3938 ( 
.A(n_3651),
.B(n_2487),
.Y(n_3938)
);

AOI22xp33_ASAP7_75t_L g3939 ( 
.A1(n_3615),
.A2(n_3396),
.B1(n_2657),
.B2(n_2546),
.Y(n_3939)
);

INVx2_ASAP7_75t_SL g3940 ( 
.A(n_3676),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_SL g3941 ( 
.A(n_3651),
.B(n_2487),
.Y(n_3941)
);

INVx2_ASAP7_75t_L g3942 ( 
.A(n_3556),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3558),
.Y(n_3943)
);

OAI22xp5_ASAP7_75t_SL g3944 ( 
.A1(n_3584),
.A2(n_1705),
.B1(n_1853),
.B2(n_1822),
.Y(n_3944)
);

A2O1A1Ixp33_ASAP7_75t_L g3945 ( 
.A1(n_3800),
.A2(n_3004),
.B(n_3405),
.C(n_3341),
.Y(n_3945)
);

AND2x4_ASAP7_75t_L g3946 ( 
.A(n_3648),
.B(n_3080),
.Y(n_3946)
);

INVx2_ASAP7_75t_L g3947 ( 
.A(n_3559),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3490),
.B(n_2999),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3555),
.B(n_3010),
.Y(n_3949)
);

AOI22xp33_ASAP7_75t_L g3950 ( 
.A1(n_3444),
.A2(n_2657),
.B1(n_3060),
.B2(n_2828),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3560),
.B(n_3010),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3525),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3607),
.B(n_3013),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_SL g3954 ( 
.A(n_3564),
.B(n_2487),
.Y(n_3954)
);

AOI22xp5_ASAP7_75t_L g3955 ( 
.A1(n_3711),
.A2(n_1863),
.B1(n_1872),
.B2(n_1861),
.Y(n_3955)
);

OR2x6_ASAP7_75t_L g3956 ( 
.A(n_3629),
.B(n_3152),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3563),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3611),
.B(n_3013),
.Y(n_3958)
);

AND2x2_ASAP7_75t_L g3959 ( 
.A(n_3522),
.B(n_3270),
.Y(n_3959)
);

AND2x6_ASAP7_75t_SL g3960 ( 
.A(n_3564),
.B(n_2509),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3488),
.B(n_3603),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3528),
.Y(n_3962)
);

AOI22xp5_ASAP7_75t_L g3963 ( 
.A1(n_3720),
.A2(n_1863),
.B1(n_1861),
.B2(n_2503),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3605),
.B(n_3015),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3510),
.B(n_3015),
.Y(n_3965)
);

AOI22xp33_ASAP7_75t_L g3966 ( 
.A1(n_3659),
.A2(n_2657),
.B1(n_2828),
.B2(n_2822),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3575),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_3524),
.B(n_3031),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3580),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3530),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3534),
.Y(n_3971)
);

NOR2x2_ASAP7_75t_L g3972 ( 
.A(n_3629),
.B(n_2499),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3478),
.B(n_3031),
.Y(n_3973)
);

OAI22xp5_ASAP7_75t_L g3974 ( 
.A1(n_3629),
.A2(n_3263),
.B1(n_3280),
.B2(n_3152),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3542),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3487),
.B(n_3156),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3498),
.B(n_3270),
.Y(n_3977)
);

NOR2xp33_ASAP7_75t_L g3978 ( 
.A(n_3519),
.B(n_2516),
.Y(n_3978)
);

NOR2xp33_ASAP7_75t_L g3979 ( 
.A(n_3552),
.B(n_2518),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3526),
.B(n_3164),
.Y(n_3980)
);

INVxp67_ASAP7_75t_L g3981 ( 
.A(n_3622),
.Y(n_3981)
);

NOR2xp33_ASAP7_75t_L g3982 ( 
.A(n_3552),
.B(n_2518),
.Y(n_3982)
);

BUFx3_ASAP7_75t_L g3983 ( 
.A(n_3622),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3475),
.B(n_3499),
.Y(n_3984)
);

AND2x2_ASAP7_75t_L g3985 ( 
.A(n_3576),
.B(n_3270),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3618),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_SL g3987 ( 
.A(n_3633),
.B(n_2496),
.Y(n_3987)
);

NOR2xp33_ASAP7_75t_L g3988 ( 
.A(n_3665),
.B(n_2518),
.Y(n_3988)
);

INVx1_ASAP7_75t_SL g3989 ( 
.A(n_3721),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3769),
.B(n_3191),
.Y(n_3990)
);

NOR2xp33_ASAP7_75t_L g3991 ( 
.A(n_3562),
.B(n_3264),
.Y(n_3991)
);

AND2x2_ASAP7_75t_L g3992 ( 
.A(n_3659),
.B(n_3531),
.Y(n_3992)
);

NOR3xp33_ASAP7_75t_L g3993 ( 
.A(n_3619),
.B(n_2186),
.C(n_2491),
.Y(n_3993)
);

AND2x2_ASAP7_75t_L g3994 ( 
.A(n_3531),
.B(n_2384),
.Y(n_3994)
);

INVx2_ASAP7_75t_L g3995 ( 
.A(n_3620),
.Y(n_3995)
);

INVx2_ASAP7_75t_L g3996 ( 
.A(n_3625),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3544),
.Y(n_3997)
);

AOI22xp33_ASAP7_75t_L g3998 ( 
.A1(n_3553),
.A2(n_2828),
.B1(n_2642),
.B2(n_3120),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3550),
.Y(n_3999)
);

OAI22xp5_ASAP7_75t_L g4000 ( 
.A1(n_3757),
.A2(n_3263),
.B1(n_3280),
.B2(n_3152),
.Y(n_4000)
);

INVx8_ASAP7_75t_L g4001 ( 
.A(n_3465),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3596),
.B(n_3156),
.Y(n_4002)
);

AOI22xp33_ASAP7_75t_L g4003 ( 
.A1(n_3553),
.A2(n_2642),
.B1(n_3126),
.B2(n_3122),
.Y(n_4003)
);

CKINVDCx5p33_ASAP7_75t_R g4004 ( 
.A(n_3465),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_SL g4005 ( 
.A(n_3633),
.B(n_3658),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3561),
.B(n_3445),
.Y(n_4006)
);

AO22x1_ASAP7_75t_L g4007 ( 
.A1(n_3695),
.A2(n_2359),
.B1(n_2924),
.B2(n_2612),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_SL g4008 ( 
.A(n_3658),
.B(n_2496),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3561),
.B(n_3080),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3472),
.B(n_3080),
.Y(n_4010)
);

INVx2_ASAP7_75t_SL g4011 ( 
.A(n_3592),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3598),
.B(n_3107),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_SL g4013 ( 
.A(n_3664),
.B(n_2496),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3557),
.Y(n_4014)
);

NOR2xp33_ASAP7_75t_L g4015 ( 
.A(n_3562),
.B(n_3695),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3638),
.B(n_3107),
.Y(n_4016)
);

NOR2xp33_ASAP7_75t_L g4017 ( 
.A(n_3701),
.B(n_3264),
.Y(n_4017)
);

NOR2xp33_ASAP7_75t_L g4018 ( 
.A(n_3701),
.B(n_2379),
.Y(n_4018)
);

AOI22xp5_ASAP7_75t_L g4019 ( 
.A1(n_3707),
.A2(n_2510),
.B1(n_2529),
.B2(n_2509),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_SL g4020 ( 
.A(n_3664),
.B(n_3107),
.Y(n_4020)
);

AND2x4_ASAP7_75t_L g4021 ( 
.A(n_3832),
.B(n_3011),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3693),
.B(n_3169),
.Y(n_4022)
);

BUFx3_ASAP7_75t_L g4023 ( 
.A(n_3637),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3716),
.B(n_3213),
.Y(n_4024)
);

NOR2xp33_ASAP7_75t_L g4025 ( 
.A(n_3707),
.B(n_2379),
.Y(n_4025)
);

BUFx3_ASAP7_75t_L g4026 ( 
.A(n_3780),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3572),
.Y(n_4027)
);

AND2x4_ASAP7_75t_L g4028 ( 
.A(n_3802),
.B(n_3240),
.Y(n_4028)
);

AND2x4_ASAP7_75t_L g4029 ( 
.A(n_3802),
.B(n_3668),
.Y(n_4029)
);

AOI22xp33_ASAP7_75t_L g4030 ( 
.A1(n_3578),
.A2(n_2642),
.B1(n_3179),
.B2(n_3172),
.Y(n_4030)
);

INVx2_ASAP7_75t_L g4031 ( 
.A(n_3628),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3719),
.B(n_3180),
.Y(n_4032)
);

INVx1_ASAP7_75t_SL g4033 ( 
.A(n_3727),
.Y(n_4033)
);

AOI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3715),
.A2(n_2529),
.B1(n_2510),
.B2(n_2384),
.Y(n_4034)
);

BUFx3_ASAP7_75t_L g4035 ( 
.A(n_3621),
.Y(n_4035)
);

AND2x4_ASAP7_75t_L g4036 ( 
.A(n_3668),
.B(n_3328),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3591),
.Y(n_4037)
);

BUFx6f_ASAP7_75t_L g4038 ( 
.A(n_3503),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3715),
.B(n_3729),
.Y(n_4039)
);

OR2x6_ASAP7_75t_L g4040 ( 
.A(n_3621),
.B(n_3263),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3582),
.B(n_3184),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3631),
.Y(n_4042)
);

INVx2_ASAP7_75t_L g4043 ( 
.A(n_3640),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_3582),
.B(n_3299),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3583),
.B(n_3308),
.Y(n_4045)
);

AND3x1_ASAP7_75t_L g4046 ( 
.A(n_3578),
.B(n_2498),
.C(n_2491),
.Y(n_4046)
);

BUFx6f_ASAP7_75t_L g4047 ( 
.A(n_3503),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3583),
.B(n_3325),
.Y(n_4048)
);

AOI22xp33_ASAP7_75t_L g4049 ( 
.A1(n_3684),
.A2(n_2642),
.B1(n_2980),
.B2(n_2316),
.Y(n_4049)
);

NOR2xp33_ASAP7_75t_L g4050 ( 
.A(n_3729),
.B(n_2379),
.Y(n_4050)
);

NOR2xp33_ASAP7_75t_L g4051 ( 
.A(n_3738),
.B(n_2433),
.Y(n_4051)
);

OAI22xp5_ASAP7_75t_L g4052 ( 
.A1(n_3760),
.A2(n_3263),
.B1(n_3280),
.B2(n_3257),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_SL g4053 ( 
.A(n_3738),
.B(n_2498),
.Y(n_4053)
);

AND2x6_ASAP7_75t_SL g4054 ( 
.A(n_3829),
.B(n_2142),
.Y(n_4054)
);

INVx2_ASAP7_75t_L g4055 ( 
.A(n_3644),
.Y(n_4055)
);

NOR2xp33_ASAP7_75t_L g4056 ( 
.A(n_3741),
.B(n_2433),
.Y(n_4056)
);

BUFx6f_ASAP7_75t_L g4057 ( 
.A(n_3503),
.Y(n_4057)
);

NOR2xp33_ASAP7_75t_L g4058 ( 
.A(n_3741),
.B(n_2433),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3589),
.B(n_3046),
.Y(n_4059)
);

NAND2x1_ASAP7_75t_L g4060 ( 
.A(n_3502),
.B(n_3001),
.Y(n_4060)
);

CKINVDCx5p33_ASAP7_75t_R g4061 ( 
.A(n_3473),
.Y(n_4061)
);

AND2x6_ASAP7_75t_SL g4062 ( 
.A(n_3829),
.B(n_3214),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3589),
.B(n_3594),
.Y(n_4063)
);

BUFx6f_ASAP7_75t_L g4064 ( 
.A(n_3508),
.Y(n_4064)
);

NOR2xp33_ASAP7_75t_L g4065 ( 
.A(n_3748),
.B(n_2433),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_SL g4066 ( 
.A(n_3748),
.B(n_2359),
.Y(n_4066)
);

AND2x4_ASAP7_75t_SL g4067 ( 
.A(n_3464),
.B(n_3280),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3593),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3706),
.B(n_3047),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_3752),
.B(n_2387),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3712),
.B(n_3167),
.Y(n_4071)
);

AND2x6_ASAP7_75t_SL g4072 ( 
.A(n_3755),
.B(n_3772),
.Y(n_4072)
);

AOI21xp5_ASAP7_75t_L g4073 ( 
.A1(n_3450),
.A2(n_3398),
.B(n_3391),
.Y(n_4073)
);

AOI22xp5_ASAP7_75t_L g4074 ( 
.A1(n_3755),
.A2(n_2418),
.B1(n_2175),
.B2(n_2141),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3623),
.B(n_3192),
.Y(n_4075)
);

AND2x2_ASAP7_75t_L g4076 ( 
.A(n_3772),
.B(n_2526),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_SL g4077 ( 
.A(n_3661),
.B(n_3173),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3597),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_3684),
.A2(n_2642),
.B1(n_2316),
.B2(n_2997),
.Y(n_4079)
);

AOI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_3783),
.A2(n_2418),
.B1(n_2380),
.B2(n_2333),
.Y(n_4080)
);

NAND2x1_ASAP7_75t_L g4081 ( 
.A(n_3801),
.B(n_3001),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3599),
.B(n_3167),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_3600),
.B(n_3191),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3601),
.B(n_3192),
.Y(n_4084)
);

INVxp33_ASAP7_75t_L g4085 ( 
.A(n_3830),
.Y(n_4085)
);

NOR2xp33_ASAP7_75t_L g4086 ( 
.A(n_3641),
.B(n_1886),
.Y(n_4086)
);

AOI22xp5_ASAP7_75t_L g4087 ( 
.A1(n_3617),
.A2(n_2380),
.B1(n_2333),
.B2(n_2245),
.Y(n_4087)
);

HB1xp67_ASAP7_75t_L g4088 ( 
.A(n_3641),
.Y(n_4088)
);

NOR2xp33_ASAP7_75t_L g4089 ( 
.A(n_3781),
.B(n_1886),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3602),
.B(n_3157),
.Y(n_4090)
);

AOI21xp5_ASAP7_75t_L g4091 ( 
.A1(n_3489),
.A2(n_3398),
.B(n_3391),
.Y(n_4091)
);

BUFx3_ASAP7_75t_L g4092 ( 
.A(n_3571),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_SL g4093 ( 
.A(n_3624),
.B(n_2612),
.Y(n_4093)
);

INVx2_ASAP7_75t_L g4094 ( 
.A(n_3647),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3612),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_SL g4096 ( 
.A(n_3751),
.B(n_2924),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3635),
.B(n_3157),
.Y(n_4097)
);

OAI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3761),
.A2(n_2997),
.B1(n_3061),
.B2(n_3202),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_3713),
.B(n_2918),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3646),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3649),
.Y(n_4101)
);

NAND3xp33_ASAP7_75t_SL g4102 ( 
.A(n_3669),
.B(n_1923),
.C(n_1921),
.Y(n_4102)
);

BUFx6f_ASAP7_75t_L g4103 ( 
.A(n_3508),
.Y(n_4103)
);

BUFx3_ASAP7_75t_L g4104 ( 
.A(n_3464),
.Y(n_4104)
);

AOI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_3456),
.A2(n_2380),
.B1(n_2245),
.B2(n_1923),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_3653),
.B(n_3194),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_3655),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_3660),
.B(n_3194),
.Y(n_4108)
);

INVx2_ASAP7_75t_L g4109 ( 
.A(n_3652),
.Y(n_4109)
);

AOI22xp33_ASAP7_75t_L g4110 ( 
.A1(n_3669),
.A2(n_2997),
.B1(n_3061),
.B2(n_2971),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_3667),
.B(n_3164),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3670),
.B(n_3213),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_3656),
.Y(n_4113)
);

INVx2_ASAP7_75t_L g4114 ( 
.A(n_3657),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3671),
.B(n_3215),
.Y(n_4115)
);

NAND3xp33_ASAP7_75t_L g4116 ( 
.A(n_3675),
.B(n_3401),
.C(n_3054),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3673),
.Y(n_4117)
);

O2A1O1Ixp5_ASAP7_75t_L g4118 ( 
.A1(n_3527),
.A2(n_3009),
.B(n_3341),
.C(n_3202),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_3680),
.B(n_3186),
.Y(n_4119)
);

NOR2xp67_ASAP7_75t_SL g4120 ( 
.A(n_3443),
.B(n_3313),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3682),
.B(n_3186),
.Y(n_4121)
);

AND2x4_ASAP7_75t_L g4122 ( 
.A(n_3713),
.B(n_3328),
.Y(n_4122)
);

NOR2xp33_ASAP7_75t_L g4123 ( 
.A(n_3781),
.B(n_1921),
.Y(n_4123)
);

INVx2_ASAP7_75t_SL g4124 ( 
.A(n_3685),
.Y(n_4124)
);

AOI22xp33_ASAP7_75t_L g4125 ( 
.A1(n_3675),
.A2(n_3061),
.B1(n_2971),
.B2(n_2846),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3688),
.Y(n_4126)
);

INVx2_ASAP7_75t_SL g4127 ( 
.A(n_3698),
.Y(n_4127)
);

AOI22xp33_ASAP7_75t_L g4128 ( 
.A1(n_3678),
.A2(n_3824),
.B1(n_3474),
.B2(n_3486),
.Y(n_4128)
);

INVxp67_ASAP7_75t_L g4129 ( 
.A(n_3473),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_L g4130 ( 
.A(n_3694),
.B(n_3190),
.Y(n_4130)
);

AND2x6_ASAP7_75t_SL g4131 ( 
.A(n_3806),
.B(n_3098),
.Y(n_4131)
);

AOI21xp5_ASAP7_75t_L g4132 ( 
.A1(n_3509),
.A2(n_3403),
.B(n_3344),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_3702),
.B(n_3196),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3703),
.B(n_3196),
.Y(n_4134)
);

AND2x6_ASAP7_75t_SL g4135 ( 
.A(n_3806),
.B(n_3273),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3732),
.B(n_3215),
.Y(n_4136)
);

AND2x6_ASAP7_75t_SL g4137 ( 
.A(n_3818),
.B(n_3273),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3734),
.B(n_3190),
.Y(n_4138)
);

AOI22xp33_ASAP7_75t_L g4139 ( 
.A1(n_3678),
.A2(n_3061),
.B1(n_2971),
.B2(n_2850),
.Y(n_4139)
);

NOR2x2_ASAP7_75t_L g4140 ( 
.A(n_3689),
.B(n_3318),
.Y(n_4140)
);

NOR2xp33_ASAP7_75t_L g4141 ( 
.A(n_3466),
.B(n_1926),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3739),
.B(n_3227),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3742),
.B(n_3227),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_3747),
.B(n_3210),
.Y(n_4144)
);

AND2x4_ASAP7_75t_L g4145 ( 
.A(n_3705),
.B(n_3406),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_3818),
.B(n_3081),
.Y(n_4146)
);

CKINVDCx5p33_ASAP7_75t_R g4147 ( 
.A(n_3616),
.Y(n_4147)
);

NOR2xp33_ASAP7_75t_L g4148 ( 
.A(n_3568),
.B(n_1926),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3749),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3763),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_SL g4151 ( 
.A(n_3754),
.B(n_3064),
.Y(n_4151)
);

NOR2xp33_ASAP7_75t_L g4152 ( 
.A(n_3570),
.B(n_2844),
.Y(n_4152)
);

OAI21xp5_ASAP7_75t_L g4153 ( 
.A1(n_3833),
.A2(n_3096),
.B(n_3094),
.Y(n_4153)
);

OAI21xp5_ASAP7_75t_L g4154 ( 
.A1(n_3722),
.A2(n_3312),
.B(n_3008),
.Y(n_4154)
);

INVx2_ASAP7_75t_SL g4155 ( 
.A(n_3714),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_3626),
.B(n_2798),
.Y(n_4156)
);

NAND2x1p5_ASAP7_75t_L g4157 ( 
.A(n_3794),
.B(n_3016),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3476),
.B(n_2798),
.Y(n_4158)
);

AOI22xp5_ASAP7_75t_L g4159 ( 
.A1(n_3469),
.A2(n_3403),
.B1(n_3442),
.B2(n_3408),
.Y(n_4159)
);

AND2x2_ASAP7_75t_SL g4160 ( 
.A(n_3513),
.B(n_3442),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_3700),
.B(n_2801),
.Y(n_4161)
);

INVx2_ASAP7_75t_SL g4162 ( 
.A(n_3737),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_3586),
.B(n_2918),
.Y(n_4163)
);

AND2x6_ASAP7_75t_SL g4164 ( 
.A(n_3492),
.B(n_859),
.Y(n_4164)
);

AOI22xp33_ASAP7_75t_L g4165 ( 
.A1(n_3759),
.A2(n_2860),
.B1(n_2861),
.B2(n_2857),
.Y(n_4165)
);

OR2x6_ASAP7_75t_L g4166 ( 
.A(n_3835),
.B(n_3643),
.Y(n_4166)
);

OR2x2_ASAP7_75t_L g4167 ( 
.A(n_3679),
.B(n_2918),
.Y(n_4167)
);

OAI22xp5_ASAP7_75t_L g4168 ( 
.A1(n_3765),
.A2(n_2991),
.B1(n_3070),
.B2(n_3045),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_3764),
.Y(n_4169)
);

NOR2xp33_ASAP7_75t_L g4170 ( 
.A(n_3595),
.B(n_2865),
.Y(n_4170)
);

AOI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_3549),
.A2(n_3344),
.B(n_3313),
.Y(n_4171)
);

OAI22xp5_ASAP7_75t_SL g4172 ( 
.A1(n_3541),
.A2(n_1273),
.B1(n_1231),
.B2(n_1049),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_SL g4173 ( 
.A(n_3548),
.B(n_3771),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_3766),
.B(n_3210),
.Y(n_4174)
);

OR2x2_ASAP7_75t_L g4175 ( 
.A(n_3567),
.B(n_2918),
.Y(n_4175)
);

NOR2xp33_ASAP7_75t_SL g4176 ( 
.A(n_3616),
.B(n_3588),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_SL g4177 ( 
.A(n_3681),
.B(n_3627),
.Y(n_4177)
);

INVx2_ASAP7_75t_L g4178 ( 
.A(n_3708),
.Y(n_4178)
);

BUFx10_ASAP7_75t_L g4179 ( 
.A(n_3543),
.Y(n_4179)
);

NOR3xp33_ASAP7_75t_L g4180 ( 
.A(n_3745),
.B(n_2871),
.C(n_2869),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3717),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_3774),
.B(n_2801),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3724),
.Y(n_4183)
);

AOI22xp5_ASAP7_75t_L g4184 ( 
.A1(n_3718),
.A2(n_3408),
.B1(n_3370),
.B2(n_3372),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_3775),
.B(n_2803),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3728),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_SL g4187 ( 
.A(n_3632),
.B(n_3016),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3756),
.B(n_3225),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_3690),
.B(n_2803),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_3731),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_3691),
.B(n_2805),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_SL g4192 ( 
.A(n_3634),
.B(n_3016),
.Y(n_4192)
);

NOR2xp33_ASAP7_75t_L g4193 ( 
.A(n_3799),
.B(n_2873),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_3733),
.Y(n_4194)
);

OAI22xp5_ASAP7_75t_L g4195 ( 
.A1(n_3692),
.A2(n_3023),
.B1(n_3114),
.B2(n_3102),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_3740),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3709),
.B(n_3225),
.Y(n_4197)
);

NAND3xp33_ASAP7_75t_SL g4198 ( 
.A(n_3604),
.B(n_3241),
.C(n_3232),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_3744),
.Y(n_4199)
);

NOR2xp33_ASAP7_75t_SL g4200 ( 
.A(n_3543),
.B(n_3408),
.Y(n_4200)
);

INVx2_ASAP7_75t_SL g4201 ( 
.A(n_3737),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_3736),
.B(n_3318),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_SL g4203 ( 
.A(n_3642),
.B(n_3016),
.Y(n_4203)
);

OAI22xp33_ASAP7_75t_L g4204 ( 
.A1(n_3696),
.A2(n_3142),
.B1(n_3146),
.B2(n_3138),
.Y(n_4204)
);

CKINVDCx5p33_ASAP7_75t_R g4205 ( 
.A(n_3753),
.Y(n_4205)
);

OAI22xp33_ASAP7_75t_L g4206 ( 
.A1(n_3699),
.A2(n_3197),
.B1(n_3200),
.B2(n_3189),
.Y(n_4206)
);

AOI22xp5_ASAP7_75t_L g4207 ( 
.A1(n_3725),
.A2(n_3370),
.B1(n_3372),
.B2(n_3362),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_3750),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_3855),
.B(n_4039),
.Y(n_4209)
);

AOI21xp5_ASAP7_75t_L g4210 ( 
.A1(n_4073),
.A2(n_3569),
.B(n_3566),
.Y(n_4210)
);

AND2x2_ASAP7_75t_L g4211 ( 
.A(n_3992),
.B(n_3604),
.Y(n_4211)
);

AOI21xp5_ASAP7_75t_L g4212 ( 
.A1(n_4091),
.A2(n_3735),
.B(n_3785),
.Y(n_4212)
);

NOR2xp33_ASAP7_75t_SL g4213 ( 
.A(n_3857),
.B(n_3092),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_3881),
.B(n_3784),
.Y(n_4214)
);

INVx2_ASAP7_75t_L g4215 ( 
.A(n_3846),
.Y(n_4215)
);

AOI21xp5_ASAP7_75t_L g4216 ( 
.A1(n_4132),
.A2(n_3614),
.B(n_3609),
.Y(n_4216)
);

AOI21xp5_ASAP7_75t_L g4217 ( 
.A1(n_4154),
.A2(n_3614),
.B(n_3609),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_3894),
.B(n_3650),
.Y(n_4218)
);

INVx5_ASAP7_75t_L g4219 ( 
.A(n_4040),
.Y(n_4219)
);

BUFx6f_ASAP7_75t_L g4220 ( 
.A(n_4001),
.Y(n_4220)
);

OAI21xp5_ASAP7_75t_L g4221 ( 
.A1(n_3912),
.A2(n_3796),
.B(n_2698),
.Y(n_4221)
);

INVx3_ASAP7_75t_L g4222 ( 
.A(n_4040),
.Y(n_4222)
);

AOI21x1_ASAP7_75t_L g4223 ( 
.A1(n_4173),
.A2(n_3639),
.B(n_3540),
.Y(n_4223)
);

OAI21xp5_ASAP7_75t_L g4224 ( 
.A1(n_3898),
.A2(n_2651),
.B(n_2744),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3841),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_SL g4226 ( 
.A(n_3925),
.B(n_3817),
.Y(n_4226)
);

INVx6_ASAP7_75t_L g4227 ( 
.A(n_3851),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_SL g4228 ( 
.A(n_3979),
.B(n_3662),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3847),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_3894),
.B(n_4063),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_4070),
.B(n_3663),
.Y(n_4231)
);

AOI22xp5_ASAP7_75t_L g4232 ( 
.A1(n_3879),
.A2(n_3654),
.B1(n_3677),
.B2(n_3805),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3852),
.Y(n_4233)
);

NAND2x1p5_ASAP7_75t_L g4234 ( 
.A(n_4120),
.B(n_3928),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_3982),
.B(n_3674),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_3961),
.B(n_3790),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_3961),
.B(n_3978),
.Y(n_4237)
);

OR2x2_ASAP7_75t_SL g4238 ( 
.A(n_4102),
.B(n_872),
.Y(n_4238)
);

OAI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_3920),
.A2(n_2651),
.B(n_2744),
.Y(n_4239)
);

OAI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_3945),
.A2(n_2880),
.B(n_2867),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_3867),
.Y(n_4241)
);

NOR2xp33_ASAP7_75t_L g4242 ( 
.A(n_3910),
.B(n_3636),
.Y(n_4242)
);

BUFx2_ASAP7_75t_SL g4243 ( 
.A(n_3909),
.Y(n_4243)
);

AOI21xp5_ASAP7_75t_L g4244 ( 
.A1(n_4171),
.A2(n_3782),
.B(n_3697),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3870),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_3889),
.B(n_4017),
.Y(n_4246)
);

AOI21xp5_ASAP7_75t_L g4247 ( 
.A1(n_4160),
.A2(n_3782),
.B(n_3697),
.Y(n_4247)
);

NAND2x1_ASAP7_75t_L g4248 ( 
.A(n_3928),
.B(n_3021),
.Y(n_4248)
);

OAI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_3863),
.A2(n_3686),
.B1(n_3683),
.B2(n_3029),
.Y(n_4249)
);

NOR2x1p5_ASAP7_75t_SL g4250 ( 
.A(n_4175),
.B(n_3518),
.Y(n_4250)
);

INVxp67_ASAP7_75t_L g4251 ( 
.A(n_4015),
.Y(n_4251)
);

AO21x1_ASAP7_75t_L g4252 ( 
.A1(n_3839),
.A2(n_3808),
.B(n_3807),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4005),
.B(n_3768),
.Y(n_4253)
);

O2A1O1Ixp33_ASAP7_75t_L g4254 ( 
.A1(n_4053),
.A2(n_788),
.B(n_829),
.C(n_755),
.Y(n_4254)
);

HB1xp67_ASAP7_75t_L g4255 ( 
.A(n_3983),
.Y(n_4255)
);

A2O1A1Ixp33_ASAP7_75t_L g4256 ( 
.A1(n_3988),
.A2(n_3814),
.B(n_3828),
.C(n_3823),
.Y(n_4256)
);

AND2x4_ASAP7_75t_L g4257 ( 
.A(n_3903),
.B(n_3946),
.Y(n_4257)
);

AOI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_4069),
.A2(n_3344),
.B(n_3313),
.Y(n_4258)
);

AOI21xp5_ASAP7_75t_L g4259 ( 
.A1(n_3840),
.A2(n_3929),
.B(n_3984),
.Y(n_4259)
);

INVx3_ASAP7_75t_L g4260 ( 
.A(n_4040),
.Y(n_4260)
);

INVx4_ASAP7_75t_L g4261 ( 
.A(n_3843),
.Y(n_4261)
);

NOR2xp33_ASAP7_75t_L g4262 ( 
.A(n_3880),
.B(n_2877),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_SL g4263 ( 
.A(n_3844),
.B(n_3777),
.Y(n_4263)
);

OR2x2_ASAP7_75t_L g4264 ( 
.A(n_4006),
.B(n_3787),
.Y(n_4264)
);

AOI22xp5_ASAP7_75t_L g4265 ( 
.A1(n_3873),
.A2(n_3786),
.B1(n_3804),
.B2(n_3803),
.Y(n_4265)
);

O2A1O1Ixp33_ASAP7_75t_L g4266 ( 
.A1(n_3866),
.A2(n_887),
.B(n_899),
.C(n_829),
.Y(n_4266)
);

AOI21xp5_ASAP7_75t_L g4267 ( 
.A1(n_3984),
.A2(n_3344),
.B(n_3313),
.Y(n_4267)
);

INVx3_ASAP7_75t_L g4268 ( 
.A(n_4067),
.Y(n_4268)
);

AND2x2_ASAP7_75t_L g4269 ( 
.A(n_3885),
.B(n_3792),
.Y(n_4269)
);

OAI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_4198),
.A2(n_2880),
.B(n_3211),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_3849),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_3888),
.Y(n_4272)
);

AOI21xp33_ASAP7_75t_L g4273 ( 
.A1(n_4044),
.A2(n_3226),
.B(n_3221),
.Y(n_4273)
);

AOI21xp5_ASAP7_75t_L g4274 ( 
.A1(n_4168),
.A2(n_3344),
.B(n_3313),
.Y(n_4274)
);

NAND2x1p5_ASAP7_75t_L g4275 ( 
.A(n_4020),
.B(n_3836),
.Y(n_4275)
);

OAI21xp33_ASAP7_75t_L g4276 ( 
.A1(n_4019),
.A2(n_2881),
.B(n_2878),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_SL g4277 ( 
.A(n_4034),
.B(n_3813),
.Y(n_4277)
);

NOR2xp33_ASAP7_75t_R g4278 ( 
.A(n_3913),
.B(n_3753),
.Y(n_4278)
);

INVx3_ASAP7_75t_L g4279 ( 
.A(n_3872),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_L g4280 ( 
.A(n_4018),
.B(n_3819),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4025),
.B(n_3834),
.Y(n_4281)
);

BUFx2_ASAP7_75t_SL g4282 ( 
.A(n_3876),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_3916),
.B(n_2884),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4050),
.B(n_3758),
.Y(n_4284)
);

AND2x2_ASAP7_75t_L g4285 ( 
.A(n_3959),
.B(n_2805),
.Y(n_4285)
);

AOI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_4168),
.A2(n_3825),
.B(n_3170),
.Y(n_4286)
);

NOR2xp33_ASAP7_75t_L g4287 ( 
.A(n_3991),
.B(n_1268),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_4051),
.B(n_3770),
.Y(n_4288)
);

NOR2xp33_ASAP7_75t_L g4289 ( 
.A(n_4148),
.B(n_1268),
.Y(n_4289)
);

INVx2_ASAP7_75t_L g4290 ( 
.A(n_3850),
.Y(n_4290)
);

AOI21xp5_ASAP7_75t_L g4291 ( 
.A1(n_4000),
.A2(n_4197),
.B(n_4048),
.Y(n_4291)
);

NOR2xp33_ASAP7_75t_L g4292 ( 
.A(n_3989),
.B(n_1268),
.Y(n_4292)
);

OAI21xp5_ASAP7_75t_L g4293 ( 
.A1(n_4153),
.A2(n_3233),
.B(n_3230),
.Y(n_4293)
);

AOI21xp5_ASAP7_75t_L g4294 ( 
.A1(n_4000),
.A2(n_3170),
.B(n_3166),
.Y(n_4294)
);

INVx2_ASAP7_75t_L g4295 ( 
.A(n_3854),
.Y(n_4295)
);

AOI21xp5_ASAP7_75t_L g4296 ( 
.A1(n_4197),
.A2(n_3170),
.B(n_3166),
.Y(n_4296)
);

OAI21xp5_ASAP7_75t_L g4297 ( 
.A1(n_4118),
.A2(n_3267),
.B(n_3234),
.Y(n_4297)
);

NOR2xp33_ASAP7_75t_L g4298 ( 
.A(n_3955),
.B(n_3822),
.Y(n_4298)
);

AOI21xp5_ASAP7_75t_L g4299 ( 
.A1(n_4045),
.A2(n_3178),
.B(n_3166),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_4056),
.B(n_3778),
.Y(n_4300)
);

OAI21xp5_ASAP7_75t_L g4301 ( 
.A1(n_4195),
.A2(n_4151),
.B(n_4128),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_4058),
.B(n_3793),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_3905),
.Y(n_4303)
);

AOI21xp5_ASAP7_75t_L g4304 ( 
.A1(n_3862),
.A2(n_3198),
.B(n_3178),
.Y(n_4304)
);

OR2x2_ASAP7_75t_L g4305 ( 
.A(n_3877),
.B(n_3447),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3927),
.Y(n_4306)
);

AOI21xp5_ASAP7_75t_L g4307 ( 
.A1(n_3862),
.A2(n_3198),
.B(n_3178),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_3952),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_3977),
.B(n_2806),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_4065),
.B(n_3798),
.Y(n_4310)
);

INVxp67_ASAP7_75t_L g4311 ( 
.A(n_4088),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3962),
.Y(n_4312)
);

NAND3xp33_ASAP7_75t_L g4313 ( 
.A(n_3993),
.B(n_939),
.C(n_938),
.Y(n_4313)
);

AOI21xp5_ASAP7_75t_L g4314 ( 
.A1(n_4156),
.A2(n_3201),
.B(n_3198),
.Y(n_4314)
);

AOI21x1_ASAP7_75t_L g4315 ( 
.A1(n_4093),
.A2(n_3746),
.B(n_3520),
.Y(n_4315)
);

AOI22xp33_ASAP7_75t_L g4316 ( 
.A1(n_4076),
.A2(n_3944),
.B1(n_3937),
.B2(n_4141),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_3970),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_3971),
.Y(n_4318)
);

INVx1_ASAP7_75t_SL g4319 ( 
.A(n_4140),
.Y(n_4319)
);

AOI21xp5_ASAP7_75t_L g4320 ( 
.A1(n_4052),
.A2(n_4206),
.B(n_4204),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3975),
.Y(n_4321)
);

INVxp67_ASAP7_75t_L g4322 ( 
.A(n_3893),
.Y(n_4322)
);

AOI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_4052),
.A2(n_3204),
.B(n_3201),
.Y(n_4323)
);

AOI21xp5_ASAP7_75t_L g4324 ( 
.A1(n_4075),
.A2(n_3204),
.B(n_3201),
.Y(n_4324)
);

NOR2xp33_ASAP7_75t_L g4325 ( 
.A(n_4072),
.B(n_3822),
.Y(n_4325)
);

AOI21xp5_ASAP7_75t_L g4326 ( 
.A1(n_4075),
.A2(n_3212),
.B(n_3204),
.Y(n_4326)
);

AOI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_3974),
.A2(n_3212),
.B(n_3071),
.Y(n_4327)
);

AOI21xp5_ASAP7_75t_L g4328 ( 
.A1(n_3974),
.A2(n_3212),
.B(n_3071),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_SL g4329 ( 
.A(n_3923),
.B(n_3518),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_3997),
.Y(n_4330)
);

BUFx3_ASAP7_75t_L g4331 ( 
.A(n_4001),
.Y(n_4331)
);

AOI21xp5_ASAP7_75t_L g4332 ( 
.A1(n_4146),
.A2(n_3071),
.B(n_3016),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_SL g4333 ( 
.A(n_3886),
.B(n_3518),
.Y(n_4333)
);

AO21x1_ASAP7_75t_L g4334 ( 
.A1(n_3926),
.A2(n_3815),
.B(n_3820),
.Y(n_4334)
);

OAI21xp5_ASAP7_75t_L g4335 ( 
.A1(n_4195),
.A2(n_3295),
.B(n_3268),
.Y(n_4335)
);

NOR2xp33_ASAP7_75t_L g4336 ( 
.A(n_3963),
.B(n_2806),
.Y(n_4336)
);

A2O1A1Ixp33_ASAP7_75t_L g4337 ( 
.A1(n_3924),
.A2(n_2813),
.B(n_2816),
.C(n_2815),
.Y(n_4337)
);

AOI21xp5_ASAP7_75t_L g4338 ( 
.A1(n_4077),
.A2(n_3085),
.B(n_3071),
.Y(n_4338)
);

A2O1A1Ixp33_ASAP7_75t_L g4339 ( 
.A1(n_3907),
.A2(n_2813),
.B(n_2816),
.C(n_2815),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_SL g4340 ( 
.A(n_3899),
.B(n_3518),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_3999),
.Y(n_4341)
);

AOI22xp5_ASAP7_75t_L g4342 ( 
.A1(n_4089),
.A2(n_3826),
.B1(n_3821),
.B2(n_2827),
.Y(n_4342)
);

OAI21xp5_ASAP7_75t_L g4343 ( 
.A1(n_4165),
.A2(n_3304),
.B(n_3285),
.Y(n_4343)
);

OAI22xp5_ASAP7_75t_L g4344 ( 
.A1(n_3896),
.A2(n_3322),
.B1(n_3321),
.B2(n_3085),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_3901),
.B(n_3809),
.Y(n_4345)
);

INVx2_ASAP7_75t_L g4346 ( 
.A(n_3864),
.Y(n_4346)
);

NOR2xp33_ASAP7_75t_L g4347 ( 
.A(n_4086),
.B(n_2826),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_SL g4348 ( 
.A(n_3904),
.B(n_3518),
.Y(n_4348)
);

AND2x2_ASAP7_75t_L g4349 ( 
.A(n_3985),
.B(n_2826),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_3994),
.B(n_4152),
.Y(n_4350)
);

BUFx12f_ASAP7_75t_L g4351 ( 
.A(n_4004),
.Y(n_4351)
);

BUFx6f_ASAP7_75t_L g4352 ( 
.A(n_4001),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4170),
.B(n_3816),
.Y(n_4353)
);

AOI21xp5_ASAP7_75t_L g4354 ( 
.A1(n_3845),
.A2(n_3085),
.B(n_3071),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_L g4355 ( 
.A(n_4032),
.B(n_3827),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_3868),
.Y(n_4356)
);

AND2x2_ASAP7_75t_L g4357 ( 
.A(n_3946),
.B(n_2827),
.Y(n_4357)
);

INVx4_ASAP7_75t_L g4358 ( 
.A(n_3843),
.Y(n_4358)
);

AO21x1_ASAP7_75t_L g4359 ( 
.A1(n_3884),
.A2(n_3387),
.B(n_3836),
.Y(n_4359)
);

NOR2xp67_ASAP7_75t_L g4360 ( 
.A(n_3892),
.B(n_3448),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_4177),
.B(n_2886),
.Y(n_4361)
);

CKINVDCx5p33_ASAP7_75t_R g4362 ( 
.A(n_4062),
.Y(n_4362)
);

NOR2xp33_ASAP7_75t_L g4363 ( 
.A(n_4123),
.B(n_2886),
.Y(n_4363)
);

INVx2_ASAP7_75t_SL g4364 ( 
.A(n_4179),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4014),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4027),
.Y(n_4366)
);

A2O1A1Ixp33_ASAP7_75t_L g4367 ( 
.A1(n_4049),
.A2(n_2887),
.B(n_2889),
.C(n_2888),
.Y(n_4367)
);

NOR2xp33_ASAP7_75t_L g4368 ( 
.A(n_4026),
.B(n_2887),
.Y(n_4368)
);

AOI21xp5_ASAP7_75t_L g4369 ( 
.A1(n_3845),
.A2(n_3110),
.B(n_3085),
.Y(n_4369)
);

AOI21xp5_ASAP7_75t_L g4370 ( 
.A1(n_4059),
.A2(n_3110),
.B(n_3085),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4037),
.Y(n_4371)
);

OAI21xp5_ASAP7_75t_L g4372 ( 
.A1(n_4002),
.A2(n_3347),
.B(n_3811),
.Y(n_4372)
);

AOI21xp5_ASAP7_75t_L g4373 ( 
.A1(n_3990),
.A2(n_3110),
.B(n_3144),
.Y(n_4373)
);

OAI22xp5_ASAP7_75t_L g4374 ( 
.A1(n_3900),
.A2(n_3321),
.B1(n_3322),
.B2(n_3110),
.Y(n_4374)
);

AOI21xp5_ASAP7_75t_L g4375 ( 
.A1(n_3990),
.A2(n_3110),
.B(n_3158),
.Y(n_4375)
);

NOR2xp33_ASAP7_75t_L g4376 ( 
.A(n_3911),
.B(n_2888),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_3931),
.B(n_3897),
.Y(n_4377)
);

AOI21xp5_ASAP7_75t_L g4378 ( 
.A1(n_4071),
.A2(n_3811),
.B(n_2985),
.Y(n_4378)
);

NOR2xp33_ASAP7_75t_L g4379 ( 
.A(n_3878),
.B(n_2889),
.Y(n_4379)
);

NOR2xp33_ASAP7_75t_L g4380 ( 
.A(n_4033),
.B(n_2892),
.Y(n_4380)
);

HB1xp67_ASAP7_75t_L g4381 ( 
.A(n_3981),
.Y(n_4381)
);

INVx2_ASAP7_75t_SL g4382 ( 
.A(n_4179),
.Y(n_4382)
);

AOI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_4071),
.A2(n_2985),
.B(n_2981),
.Y(n_4383)
);

OAI22xp5_ASAP7_75t_L g4384 ( 
.A1(n_4079),
.A2(n_3368),
.B1(n_3424),
.B2(n_3349),
.Y(n_4384)
);

NOR2xp33_ASAP7_75t_L g4385 ( 
.A(n_3895),
.B(n_2892),
.Y(n_4385)
);

OAI22xp5_ASAP7_75t_L g4386 ( 
.A1(n_3956),
.A2(n_1008),
.B1(n_1049),
.B2(n_887),
.Y(n_4386)
);

A2O1A1Ixp33_ASAP7_75t_L g4387 ( 
.A1(n_4193),
.A2(n_2897),
.B(n_2900),
.C(n_2898),
.Y(n_4387)
);

BUFx3_ASAP7_75t_L g4388 ( 
.A(n_3858),
.Y(n_4388)
);

BUFx2_ASAP7_75t_L g4389 ( 
.A(n_4029),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_SL g4390 ( 
.A(n_3917),
.B(n_3672),
.Y(n_4390)
);

AOI21xp5_ASAP7_75t_L g4391 ( 
.A1(n_3856),
.A2(n_3953),
.B(n_3958),
.Y(n_4391)
);

AOI21xp5_ASAP7_75t_L g4392 ( 
.A1(n_3856),
.A2(n_2985),
.B(n_2981),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_3874),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_3953),
.A2(n_3005),
.B(n_2981),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4068),
.Y(n_4395)
);

INVx2_ASAP7_75t_L g4396 ( 
.A(n_3883),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_SL g4397 ( 
.A(n_4074),
.B(n_3518),
.Y(n_4397)
);

OAI21xp5_ASAP7_75t_L g4398 ( 
.A1(n_4002),
.A2(n_2916),
.B(n_2738),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_4010),
.B(n_2897),
.Y(n_4399)
);

NOR2xp33_ASAP7_75t_L g4400 ( 
.A(n_3842),
.B(n_2898),
.Y(n_4400)
);

NOR2xp33_ASAP7_75t_L g4401 ( 
.A(n_3940),
.B(n_2900),
.Y(n_4401)
);

O2A1O1Ixp33_ASAP7_75t_SL g4402 ( 
.A1(n_3848),
.A2(n_3237),
.B(n_3244),
.C(n_3188),
.Y(n_4402)
);

AOI21xp5_ASAP7_75t_L g4403 ( 
.A1(n_3958),
.A2(n_3034),
.B(n_3005),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_3848),
.B(n_2901),
.Y(n_4404)
);

AOI21xp5_ASAP7_75t_L g4405 ( 
.A1(n_3861),
.A2(n_3034),
.B(n_3005),
.Y(n_4405)
);

AOI21xp5_ASAP7_75t_L g4406 ( 
.A1(n_3861),
.A2(n_3042),
.B(n_3034),
.Y(n_4406)
);

INVx2_ASAP7_75t_L g4407 ( 
.A(n_3891),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_4009),
.B(n_2901),
.Y(n_4408)
);

INVxp67_ASAP7_75t_L g4409 ( 
.A(n_4011),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_4041),
.B(n_2903),
.Y(n_4410)
);

O2A1O1Ixp33_ASAP7_75t_L g4411 ( 
.A1(n_3954),
.A2(n_1070),
.B(n_1105),
.C(n_1008),
.Y(n_4411)
);

AO21x1_ASAP7_75t_L g4412 ( 
.A1(n_3938),
.A2(n_3387),
.B(n_3249),
.Y(n_4412)
);

AND2x4_ASAP7_75t_L g4413 ( 
.A(n_3903),
.B(n_3406),
.Y(n_4413)
);

AOI21xp5_ASAP7_75t_L g4414 ( 
.A1(n_3980),
.A2(n_3153),
.B(n_3131),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_4012),
.B(n_2903),
.Y(n_4415)
);

AOI21xp5_ASAP7_75t_L g4416 ( 
.A1(n_3980),
.A2(n_3153),
.B(n_3422),
.Y(n_4416)
);

INVx11_ASAP7_75t_L g4417 ( 
.A(n_3843),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_SL g4418 ( 
.A(n_4046),
.B(n_3573),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_3914),
.Y(n_4419)
);

NOR2xp33_ASAP7_75t_R g4420 ( 
.A(n_4147),
.B(n_3508),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_3915),
.Y(n_4421)
);

AOI21xp5_ASAP7_75t_L g4422 ( 
.A1(n_4158),
.A2(n_3153),
.B(n_2785),
.Y(n_4422)
);

BUFx2_ASAP7_75t_L g4423 ( 
.A(n_4029),
.Y(n_4423)
);

AOI21xp5_ASAP7_75t_L g4424 ( 
.A1(n_3964),
.A2(n_2785),
.B(n_2765),
.Y(n_4424)
);

OAI22xp5_ASAP7_75t_L g4425 ( 
.A1(n_3956),
.A2(n_1105),
.B1(n_1135),
.B2(n_1126),
.Y(n_4425)
);

AOI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_3964),
.A2(n_2785),
.B(n_2765),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_4024),
.B(n_2904),
.Y(n_4427)
);

INVxp67_ASAP7_75t_L g4428 ( 
.A(n_3936),
.Y(n_4428)
);

AOI21xp5_ASAP7_75t_L g4429 ( 
.A1(n_4098),
.A2(n_2785),
.B(n_2765),
.Y(n_4429)
);

OAI21xp5_ASAP7_75t_L g4430 ( 
.A1(n_4188),
.A2(n_2916),
.B(n_2738),
.Y(n_4430)
);

AOI21xp5_ASAP7_75t_L g4431 ( 
.A1(n_4098),
.A2(n_2790),
.B(n_2785),
.Y(n_4431)
);

OAI21xp5_ASAP7_75t_L g4432 ( 
.A1(n_4188),
.A2(n_2738),
.B(n_2711),
.Y(n_4432)
);

OAI21xp33_ASAP7_75t_L g4433 ( 
.A1(n_3902),
.A2(n_1070),
.B(n_1126),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4024),
.B(n_2904),
.Y(n_4434)
);

AOI22xp5_ASAP7_75t_L g4435 ( 
.A1(n_4066),
.A2(n_2907),
.B1(n_3370),
.B2(n_3362),
.Y(n_4435)
);

AO21x1_ASAP7_75t_L g4436 ( 
.A1(n_3941),
.A2(n_3387),
.B(n_3251),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4078),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_3918),
.Y(n_4438)
);

NOR2xp33_ASAP7_75t_L g4439 ( 
.A(n_4092),
.B(n_2907),
.Y(n_4439)
);

NOR2xp33_ASAP7_75t_L g4440 ( 
.A(n_3987),
.B(n_1135),
.Y(n_4440)
);

AOI21xp5_ASAP7_75t_L g4441 ( 
.A1(n_3865),
.A2(n_2797),
.B(n_2790),
.Y(n_4441)
);

INVx3_ASAP7_75t_L g4442 ( 
.A(n_3872),
.Y(n_4442)
);

OAI21xp5_ASAP7_75t_L g4443 ( 
.A1(n_4163),
.A2(n_4159),
.B(n_3948),
.Y(n_4443)
);

AOI21xp5_ASAP7_75t_L g4444 ( 
.A1(n_3865),
.A2(n_2797),
.B(n_2790),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_L g4445 ( 
.A(n_4022),
.B(n_3428),
.Y(n_4445)
);

INVx4_ASAP7_75t_L g4446 ( 
.A(n_3872),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4016),
.B(n_3428),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_3922),
.Y(n_4448)
);

INVx2_ASAP7_75t_L g4449 ( 
.A(n_3930),
.Y(n_4449)
);

AOI21xp5_ASAP7_75t_L g4450 ( 
.A1(n_3887),
.A2(n_2797),
.B(n_2790),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_4008),
.B(n_3430),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4013),
.B(n_3430),
.Y(n_4452)
);

HB1xp67_ASAP7_75t_L g4453 ( 
.A(n_4036),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_3887),
.B(n_3431),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_3932),
.Y(n_4455)
);

INVx1_ASAP7_75t_SL g4456 ( 
.A(n_4036),
.Y(n_4456)
);

INVx1_ASAP7_75t_SL g4457 ( 
.A(n_4122),
.Y(n_4457)
);

INVx3_ASAP7_75t_L g4458 ( 
.A(n_3906),
.Y(n_4458)
);

INVx2_ASAP7_75t_SL g4459 ( 
.A(n_3908),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_4124),
.B(n_3431),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4095),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_4127),
.B(n_3337),
.Y(n_4462)
);

INVx1_ASAP7_75t_SL g4463 ( 
.A(n_4122),
.Y(n_4463)
);

NOR2xp33_ASAP7_75t_R g4464 ( 
.A(n_4205),
.B(n_3610),
.Y(n_4464)
);

OAI22xp5_ASAP7_75t_L g4465 ( 
.A1(n_3956),
.A2(n_1163),
.B1(n_1182),
.B2(n_1177),
.Y(n_4465)
);

AOI21xp5_ASAP7_75t_L g4466 ( 
.A1(n_4060),
.A2(n_2797),
.B(n_2790),
.Y(n_4466)
);

AOI21xp5_ASAP7_75t_L g4467 ( 
.A1(n_4081),
.A2(n_4202),
.B(n_4182),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_3934),
.Y(n_4468)
);

OAI22xp5_ASAP7_75t_L g4469 ( 
.A1(n_4100),
.A2(n_1163),
.B1(n_1182),
.B2(n_1177),
.Y(n_4469)
);

AND2x2_ASAP7_75t_L g4470 ( 
.A(n_3869),
.B(n_2843),
.Y(n_4470)
);

AOI21xp5_ASAP7_75t_L g4471 ( 
.A1(n_4202),
.A2(n_2799),
.B(n_2797),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4155),
.B(n_3337),
.Y(n_4472)
);

O2A1O1Ixp33_ASAP7_75t_L g4473 ( 
.A1(n_4096),
.A2(n_1198),
.B(n_1083),
.C(n_876),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_4189),
.B(n_3339),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_4191),
.B(n_3339),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_3869),
.B(n_2843),
.Y(n_4476)
);

AND2x6_ASAP7_75t_L g4477 ( 
.A(n_4184),
.B(n_3443),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4101),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_3948),
.B(n_3345),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4107),
.Y(n_4480)
);

AOI21xp5_ASAP7_75t_L g4481 ( 
.A1(n_4161),
.A2(n_2820),
.B(n_2799),
.Y(n_4481)
);

INVxp67_ASAP7_75t_L g4482 ( 
.A(n_4176),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_3871),
.B(n_3345),
.Y(n_4483)
);

AOI21xp5_ASAP7_75t_L g4484 ( 
.A1(n_4185),
.A2(n_2820),
.B(n_2799),
.Y(n_4484)
);

INVx1_ASAP7_75t_SL g4485 ( 
.A(n_4099),
.Y(n_4485)
);

AOI22xp5_ASAP7_75t_L g4486 ( 
.A1(n_4105),
.A2(n_3362),
.B1(n_3372),
.B2(n_3370),
.Y(n_4486)
);

BUFx4f_ASAP7_75t_L g4487 ( 
.A(n_3906),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4117),
.Y(n_4488)
);

AND2x4_ASAP7_75t_L g4489 ( 
.A(n_3860),
.B(n_3610),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4023),
.B(n_2843),
.Y(n_4490)
);

CKINVDCx5p33_ASAP7_75t_R g4491 ( 
.A(n_4061),
.Y(n_4491)
);

AOI21xp5_ASAP7_75t_L g4492 ( 
.A1(n_3949),
.A2(n_2820),
.B(n_2799),
.Y(n_4492)
);

NOR3xp33_ASAP7_75t_L g4493 ( 
.A(n_4116),
.B(n_876),
.C(n_872),
.Y(n_4493)
);

INVx2_ASAP7_75t_L g4494 ( 
.A(n_3942),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_4126),
.B(n_4149),
.Y(n_4495)
);

AOI21xp5_ASAP7_75t_L g4496 ( 
.A1(n_3949),
.A2(n_2820),
.B(n_2799),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_SL g4497 ( 
.A(n_4087),
.B(n_3672),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_4150),
.B(n_3361),
.Y(n_4498)
);

INVx3_ASAP7_75t_L g4499 ( 
.A(n_3906),
.Y(n_4499)
);

AOI21xp5_ASAP7_75t_L g4500 ( 
.A1(n_3951),
.A2(n_2825),
.B(n_2820),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4169),
.Y(n_4501)
);

AOI22xp5_ASAP7_75t_L g4502 ( 
.A1(n_4021),
.A2(n_3370),
.B1(n_3372),
.B2(n_3362),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_3943),
.Y(n_4503)
);

OAI21xp5_ASAP7_75t_L g4504 ( 
.A1(n_4125),
.A2(n_2738),
.B(n_2711),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4035),
.B(n_4145),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4181),
.Y(n_4506)
);

INVx3_ASAP7_75t_L g4507 ( 
.A(n_3921),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_SL g4508 ( 
.A(n_3950),
.B(n_3573),
.Y(n_4508)
);

INVx3_ASAP7_75t_L g4509 ( 
.A(n_3921),
.Y(n_4509)
);

AND2x2_ASAP7_75t_L g4510 ( 
.A(n_4145),
.B(n_2843),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_3947),
.B(n_3361),
.Y(n_4511)
);

NOR2xp67_ASAP7_75t_L g4512 ( 
.A(n_4162),
.B(n_3333),
.Y(n_4512)
);

AOI22xp5_ASAP7_75t_L g4513 ( 
.A1(n_4021),
.A2(n_3859),
.B1(n_4172),
.B2(n_4028),
.Y(n_4513)
);

O2A1O1Ixp5_ASAP7_75t_L g4514 ( 
.A1(n_4187),
.A2(n_2958),
.B(n_3149),
.C(n_3021),
.Y(n_4514)
);

AND2x2_ASAP7_75t_L g4515 ( 
.A(n_4028),
.B(n_1111),
.Y(n_4515)
);

OAI22xp5_ASAP7_75t_L g4516 ( 
.A1(n_4110),
.A2(n_3259),
.B1(n_3275),
.B2(n_3248),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_3951),
.B(n_3573),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_3957),
.B(n_1194),
.Y(n_4518)
);

O2A1O1Ixp33_ASAP7_75t_L g4519 ( 
.A1(n_4166),
.A2(n_4129),
.B(n_4203),
.C(n_4192),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4183),
.Y(n_4520)
);

BUFx2_ASAP7_75t_L g4521 ( 
.A(n_4104),
.Y(n_4521)
);

INVx2_ASAP7_75t_L g4522 ( 
.A(n_3967),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_3969),
.B(n_3380),
.Y(n_4523)
);

AOI21xp5_ASAP7_75t_L g4524 ( 
.A1(n_3973),
.A2(n_2855),
.B(n_2825),
.Y(n_4524)
);

INVx2_ASAP7_75t_L g4525 ( 
.A(n_3986),
.Y(n_4525)
);

OAI321xp33_ASAP7_75t_L g4526 ( 
.A1(n_4030),
.A2(n_3998),
.A3(n_894),
.B1(n_884),
.B2(n_898),
.C(n_893),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_3965),
.B(n_3380),
.Y(n_4527)
);

NOR2xp33_ASAP7_75t_L g4528 ( 
.A(n_3960),
.B(n_942),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_SL g4529 ( 
.A(n_3966),
.B(n_3573),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_3965),
.B(n_3385),
.Y(n_4530)
);

AOI21xp5_ASAP7_75t_L g4531 ( 
.A1(n_3973),
.A2(n_2855),
.B(n_2825),
.Y(n_4531)
);

BUFx6f_ASAP7_75t_L g4532 ( 
.A(n_4038),
.Y(n_4532)
);

O2A1O1Ixp33_ASAP7_75t_L g4533 ( 
.A1(n_4166),
.A2(n_884),
.B(n_893),
.C(n_881),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_3968),
.B(n_3385),
.Y(n_4534)
);

NAND2xp5_ASAP7_75t_SL g4535 ( 
.A(n_4200),
.B(n_4080),
.Y(n_4535)
);

BUFx6f_ASAP7_75t_L g4536 ( 
.A(n_4038),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_3968),
.B(n_3386),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_3995),
.B(n_3386),
.Y(n_4538)
);

A2O1A1Ixp33_ASAP7_75t_L g4539 ( 
.A1(n_4003),
.A2(n_3291),
.B(n_3359),
.C(n_3277),
.Y(n_4539)
);

AOI21xp5_ASAP7_75t_L g4540 ( 
.A1(n_3976),
.A2(n_2855),
.B(n_2825),
.Y(n_4540)
);

BUFx6f_ASAP7_75t_L g4541 ( 
.A(n_4038),
.Y(n_4541)
);

A2O1A1Ixp33_ASAP7_75t_L g4542 ( 
.A1(n_3939),
.A2(n_3378),
.B(n_3379),
.C(n_3365),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_3996),
.B(n_3388),
.Y(n_4543)
);

BUFx2_ASAP7_75t_SL g4544 ( 
.A(n_3875),
.Y(n_4544)
);

INVx3_ASAP7_75t_L g4545 ( 
.A(n_4047),
.Y(n_4545)
);

AOI21xp5_ASAP7_75t_L g4546 ( 
.A1(n_3976),
.A2(n_2855),
.B(n_2825),
.Y(n_4546)
);

NOR2xp33_ASAP7_75t_L g4547 ( 
.A(n_4135),
.B(n_943),
.Y(n_4547)
);

AO21x1_ASAP7_75t_L g4548 ( 
.A1(n_4167),
.A2(n_3317),
.B(n_3315),
.Y(n_4548)
);

INVx3_ASAP7_75t_L g4549 ( 
.A(n_4047),
.Y(n_4549)
);

BUFx3_ASAP7_75t_L g4550 ( 
.A(n_4047),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4186),
.Y(n_4551)
);

AND2x4_ASAP7_75t_L g4552 ( 
.A(n_4201),
.B(n_4166),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_SL g4553 ( 
.A(n_4085),
.B(n_3630),
.Y(n_4553)
);

AOI22xp5_ASAP7_75t_L g4554 ( 
.A1(n_3890),
.A2(n_3370),
.B1(n_3372),
.B2(n_3362),
.Y(n_4554)
);

HB1xp67_ASAP7_75t_L g4555 ( 
.A(n_4031),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4190),
.Y(n_4556)
);

NAND2xp5_ASAP7_75t_SL g4557 ( 
.A(n_3919),
.B(n_3645),
.Y(n_4557)
);

AOI21xp5_ASAP7_75t_L g4558 ( 
.A1(n_3935),
.A2(n_2863),
.B(n_2855),
.Y(n_4558)
);

AND2x2_ASAP7_75t_SL g4559 ( 
.A(n_4139),
.B(n_3443),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4042),
.Y(n_4560)
);

O2A1O1Ixp33_ASAP7_75t_L g4561 ( 
.A1(n_4180),
.A2(n_894),
.B(n_898),
.C(n_881),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_4043),
.B(n_4055),
.Y(n_4562)
);

INVxp67_ASAP7_75t_L g4563 ( 
.A(n_4194),
.Y(n_4563)
);

AOI21xp5_ASAP7_75t_L g4564 ( 
.A1(n_4157),
.A2(n_2908),
.B(n_2863),
.Y(n_4564)
);

INVx4_ASAP7_75t_L g4565 ( 
.A(n_4057),
.Y(n_4565)
);

A2O1A1Ixp33_ASAP7_75t_L g4566 ( 
.A1(n_4207),
.A2(n_2653),
.B(n_2601),
.C(n_2952),
.Y(n_4566)
);

BUFx6f_ASAP7_75t_L g4567 ( 
.A(n_4057),
.Y(n_4567)
);

AOI21xp5_ASAP7_75t_L g4568 ( 
.A1(n_4157),
.A2(n_2908),
.B(n_2863),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_4094),
.B(n_3388),
.Y(n_4569)
);

INVx3_ASAP7_75t_L g4570 ( 
.A(n_4057),
.Y(n_4570)
);

AOI21xp5_ASAP7_75t_L g4571 ( 
.A1(n_3838),
.A2(n_2908),
.B(n_2863),
.Y(n_4571)
);

AOI21xp5_ASAP7_75t_L g4572 ( 
.A1(n_3838),
.A2(n_2908),
.B(n_2863),
.Y(n_4572)
);

OAI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_4082),
.A2(n_2711),
.B(n_3315),
.Y(n_4573)
);

AOI21xp5_ASAP7_75t_L g4574 ( 
.A1(n_3853),
.A2(n_3933),
.B(n_4138),
.Y(n_4574)
);

AOI21xp5_ASAP7_75t_L g4575 ( 
.A1(n_3853),
.A2(n_2940),
.B(n_2908),
.Y(n_4575)
);

AOI21xp5_ASAP7_75t_L g4576 ( 
.A1(n_3933),
.A2(n_2945),
.B(n_2940),
.Y(n_4576)
);

OAI22xp5_ASAP7_75t_L g4577 ( 
.A1(n_4082),
.A2(n_3021),
.B1(n_3175),
.B2(n_3149),
.Y(n_4577)
);

OAI21xp5_ASAP7_75t_L g4578 ( 
.A1(n_4083),
.A2(n_2711),
.B(n_3317),
.Y(n_4578)
);

NOR2xp33_ASAP7_75t_L g4579 ( 
.A(n_4137),
.B(n_4131),
.Y(n_4579)
);

AOI21xp5_ASAP7_75t_L g4580 ( 
.A1(n_4083),
.A2(n_2945),
.B(n_2940),
.Y(n_4580)
);

AOI21xp5_ASAP7_75t_L g4581 ( 
.A1(n_4084),
.A2(n_2945),
.B(n_2940),
.Y(n_4581)
);

AND2x4_ASAP7_75t_L g4582 ( 
.A(n_4109),
.B(n_3610),
.Y(n_4582)
);

OAI21xp33_ASAP7_75t_L g4583 ( 
.A1(n_4196),
.A2(n_951),
.B(n_949),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_L g4584 ( 
.A(n_4113),
.B(n_3390),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4199),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_SL g4586 ( 
.A(n_4208),
.B(n_3573),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4114),
.B(n_3390),
.Y(n_4587)
);

AOI21xp5_ASAP7_75t_L g4588 ( 
.A1(n_4084),
.A2(n_2945),
.B(n_2940),
.Y(n_4588)
);

AOI21x1_ASAP7_75t_L g4589 ( 
.A1(n_4090),
.A2(n_3746),
.B(n_3520),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_SL g4590 ( 
.A(n_4178),
.B(n_3672),
.Y(n_4590)
);

AOI21xp5_ASAP7_75t_L g4591 ( 
.A1(n_4090),
.A2(n_2964),
.B(n_2945),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4064),
.B(n_1194),
.Y(n_4592)
);

INVx11_ASAP7_75t_L g4593 ( 
.A(n_4064),
.Y(n_4593)
);

O2A1O1Ixp33_ASAP7_75t_L g4594 ( 
.A1(n_4097),
.A2(n_903),
.B(n_905),
.C(n_900),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_3882),
.B(n_3402),
.Y(n_4595)
);

AOI21xp5_ASAP7_75t_L g4596 ( 
.A1(n_4097),
.A2(n_4119),
.B(n_4115),
.Y(n_4596)
);

NAND2xp5_ASAP7_75t_L g4597 ( 
.A(n_4106),
.B(n_4119),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_4106),
.B(n_3402),
.Y(n_4598)
);

AOI21xp5_ASAP7_75t_L g4599 ( 
.A1(n_4108),
.A2(n_2966),
.B(n_2964),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4108),
.B(n_3412),
.Y(n_4600)
);

AOI21xp5_ASAP7_75t_L g4601 ( 
.A1(n_4111),
.A2(n_4136),
.B(n_4134),
.Y(n_4601)
);

AOI22xp33_ASAP7_75t_L g4602 ( 
.A1(n_4111),
.A2(n_3372),
.B1(n_3362),
.B2(n_1201),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4064),
.B(n_1194),
.Y(n_4603)
);

BUFx3_ASAP7_75t_L g4604 ( 
.A(n_4521),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4215),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4225),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_SL g4607 ( 
.A(n_4237),
.B(n_4235),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4230),
.B(n_4112),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_4209),
.B(n_4242),
.Y(n_4609)
);

BUFx3_ASAP7_75t_L g4610 ( 
.A(n_4220),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4505),
.B(n_4103),
.Y(n_4611)
);

AOI22xp33_ASAP7_75t_L g4612 ( 
.A1(n_4226),
.A2(n_1194),
.B1(n_903),
.B2(n_905),
.Y(n_4612)
);

BUFx2_ASAP7_75t_L g4613 ( 
.A(n_4453),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_4271),
.Y(n_4614)
);

BUFx3_ASAP7_75t_L g4615 ( 
.A(n_4220),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_4485),
.B(n_4112),
.Y(n_4616)
);

HB1xp67_ASAP7_75t_L g4617 ( 
.A(n_4485),
.Y(n_4617)
);

OR2x6_ASAP7_75t_L g4618 ( 
.A(n_4320),
.B(n_4007),
.Y(n_4618)
);

HB1xp67_ASAP7_75t_L g4619 ( 
.A(n_4315),
.Y(n_4619)
);

INVx2_ASAP7_75t_L g4620 ( 
.A(n_4290),
.Y(n_4620)
);

NOR2xp67_ASAP7_75t_L g4621 ( 
.A(n_4482),
.B(n_4103),
.Y(n_4621)
);

NAND2xp5_ASAP7_75t_L g4622 ( 
.A(n_4214),
.B(n_4115),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4269),
.B(n_4211),
.Y(n_4623)
);

BUFx2_ASAP7_75t_L g4624 ( 
.A(n_4389),
.Y(n_4624)
);

INVx4_ASAP7_75t_L g4625 ( 
.A(n_4593),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4291),
.B(n_4121),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4391),
.B(n_4121),
.Y(n_4627)
);

AOI22xp33_ASAP7_75t_L g4628 ( 
.A1(n_4289),
.A2(n_909),
.B1(n_910),
.B2(n_900),
.Y(n_4628)
);

NOR2x1p5_ASAP7_75t_L g4629 ( 
.A(n_4331),
.B(n_3972),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4229),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4233),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4236),
.B(n_4130),
.Y(n_4632)
);

BUFx2_ASAP7_75t_L g4633 ( 
.A(n_4423),
.Y(n_4633)
);

CKINVDCx8_ASAP7_75t_R g4634 ( 
.A(n_4243),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4241),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_4218),
.B(n_4597),
.Y(n_4636)
);

INVx1_ASAP7_75t_SL g4637 ( 
.A(n_4456),
.Y(n_4637)
);

AND2x4_ASAP7_75t_L g4638 ( 
.A(n_4279),
.B(n_4103),
.Y(n_4638)
);

AND2x6_ASAP7_75t_SL g4639 ( 
.A(n_4579),
.B(n_4325),
.Y(n_4639)
);

INVx3_ASAP7_75t_L g4640 ( 
.A(n_4261),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4295),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4245),
.Y(n_4642)
);

AOI21xp5_ASAP7_75t_L g4643 ( 
.A1(n_4210),
.A2(n_2653),
.B(n_2601),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4283),
.B(n_909),
.Y(n_4644)
);

INVx5_ASAP7_75t_L g4645 ( 
.A(n_4477),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4596),
.B(n_4133),
.Y(n_4646)
);

INVx3_ASAP7_75t_L g4647 ( 
.A(n_4261),
.Y(n_4647)
);

INVx1_ASAP7_75t_SL g4648 ( 
.A(n_4456),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4601),
.B(n_4133),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4272),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4301),
.B(n_4134),
.Y(n_4651)
);

AOI22xp5_ASAP7_75t_L g4652 ( 
.A1(n_4287),
.A2(n_953),
.B1(n_955),
.B2(n_952),
.Y(n_4652)
);

INVx2_ASAP7_75t_L g4653 ( 
.A(n_4346),
.Y(n_4653)
);

AND2x2_ASAP7_75t_L g4654 ( 
.A(n_4457),
.B(n_910),
.Y(n_4654)
);

BUFx4f_ASAP7_75t_L g4655 ( 
.A(n_4220),
.Y(n_4655)
);

HB1xp67_ASAP7_75t_L g4656 ( 
.A(n_4381),
.Y(n_4656)
);

AND2x4_ASAP7_75t_L g4657 ( 
.A(n_4279),
.B(n_3710),
.Y(n_4657)
);

AND2x6_ASAP7_75t_L g4658 ( 
.A(n_4502),
.B(n_3443),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4303),
.Y(n_4659)
);

AOI22xp33_ASAP7_75t_L g4660 ( 
.A1(n_4528),
.A2(n_913),
.B1(n_915),
.B2(n_912),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4306),
.Y(n_4661)
);

BUFx3_ASAP7_75t_L g4662 ( 
.A(n_4352),
.Y(n_4662)
);

INVx2_ASAP7_75t_L g4663 ( 
.A(n_4356),
.Y(n_4663)
);

INVx3_ASAP7_75t_L g4664 ( 
.A(n_4358),
.Y(n_4664)
);

NOR2xp33_ASAP7_75t_R g4665 ( 
.A(n_4491),
.B(n_4362),
.Y(n_4665)
);

INVx4_ASAP7_75t_L g4666 ( 
.A(n_4417),
.Y(n_4666)
);

BUFx2_ASAP7_75t_L g4667 ( 
.A(n_4255),
.Y(n_4667)
);

NOR2xp33_ASAP7_75t_SL g4668 ( 
.A(n_4219),
.B(n_3092),
.Y(n_4668)
);

INVx2_ASAP7_75t_SL g4669 ( 
.A(n_4227),
.Y(n_4669)
);

HB1xp67_ASAP7_75t_L g4670 ( 
.A(n_4285),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4301),
.B(n_4443),
.Y(n_4671)
);

NOR2xp33_ASAP7_75t_L g4672 ( 
.A(n_4246),
.B(n_4054),
.Y(n_4672)
);

BUFx8_ASAP7_75t_L g4673 ( 
.A(n_4351),
.Y(n_4673)
);

INVx2_ASAP7_75t_L g4674 ( 
.A(n_4393),
.Y(n_4674)
);

NAND2xp33_ASAP7_75t_L g4675 ( 
.A(n_4352),
.B(n_3092),
.Y(n_4675)
);

OR2x6_ASAP7_75t_L g4676 ( 
.A(n_4259),
.B(n_4142),
.Y(n_4676)
);

CKINVDCx20_ASAP7_75t_R g4677 ( 
.A(n_4278),
.Y(n_4677)
);

BUFx2_ASAP7_75t_L g4678 ( 
.A(n_4464),
.Y(n_4678)
);

BUFx3_ASAP7_75t_L g4679 ( 
.A(n_4352),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4396),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4308),
.Y(n_4681)
);

BUFx6f_ASAP7_75t_L g4682 ( 
.A(n_4532),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4443),
.B(n_4142),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4350),
.B(n_4143),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_L g4685 ( 
.A(n_4228),
.B(n_4143),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4404),
.B(n_4144),
.Y(n_4686)
);

CKINVDCx5p33_ASAP7_75t_R g4687 ( 
.A(n_4420),
.Y(n_4687)
);

CKINVDCx5p33_ASAP7_75t_R g4688 ( 
.A(n_4282),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_L g4689 ( 
.A(n_4355),
.B(n_4144),
.Y(n_4689)
);

OR2x2_ASAP7_75t_L g4690 ( 
.A(n_4231),
.B(n_4174),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_4407),
.Y(n_4691)
);

BUFx8_ASAP7_75t_SL g4692 ( 
.A(n_4388),
.Y(n_4692)
);

AND2x4_ASAP7_75t_L g4693 ( 
.A(n_4442),
.B(n_3710),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_SL g4694 ( 
.A(n_4400),
.B(n_3573),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4353),
.B(n_3327),
.Y(n_4695)
);

AOI22x1_ASAP7_75t_L g4696 ( 
.A1(n_4319),
.A2(n_958),
.B1(n_959),
.B2(n_957),
.Y(n_4696)
);

INVx5_ASAP7_75t_L g4697 ( 
.A(n_4477),
.Y(n_4697)
);

OAI221xp5_ASAP7_75t_L g4698 ( 
.A1(n_4266),
.A2(n_915),
.B1(n_917),
.B2(n_913),
.C(n_912),
.Y(n_4698)
);

AND2x2_ASAP7_75t_L g4699 ( 
.A(n_4457),
.B(n_917),
.Y(n_4699)
);

OAI21xp5_ASAP7_75t_L g4700 ( 
.A1(n_4343),
.A2(n_2953),
.B(n_2952),
.Y(n_4700)
);

BUFx6f_ASAP7_75t_L g4701 ( 
.A(n_4532),
.Y(n_4701)
);

NOR2xp67_ASAP7_75t_L g4702 ( 
.A(n_4428),
.B(n_3412),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_4517),
.B(n_3327),
.Y(n_4703)
);

INVx2_ASAP7_75t_L g4704 ( 
.A(n_4419),
.Y(n_4704)
);

OR2x2_ASAP7_75t_L g4705 ( 
.A(n_4264),
.B(n_3329),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4312),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4317),
.Y(n_4707)
);

INVx3_ASAP7_75t_L g4708 ( 
.A(n_4358),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4318),
.Y(n_4709)
);

INVx2_ASAP7_75t_SL g4710 ( 
.A(n_4227),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4321),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4517),
.B(n_3329),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4421),
.Y(n_4713)
);

OAI22xp5_ASAP7_75t_L g4714 ( 
.A1(n_4559),
.A2(n_923),
.B1(n_924),
.B2(n_922),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4454),
.B(n_3330),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4438),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4448),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4330),
.Y(n_4718)
);

INVxp67_ASAP7_75t_L g4719 ( 
.A(n_4379),
.Y(n_4719)
);

OAI22xp5_ASAP7_75t_L g4720 ( 
.A1(n_4251),
.A2(n_923),
.B1(n_924),
.B2(n_922),
.Y(n_4720)
);

OR2x6_ASAP7_75t_L g4721 ( 
.A(n_4429),
.B(n_4431),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4341),
.Y(n_4722)
);

OAI22xp5_ASAP7_75t_L g4723 ( 
.A1(n_4386),
.A2(n_954),
.B1(n_962),
.B2(n_934),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4365),
.Y(n_4724)
);

BUFx4f_ASAP7_75t_L g4725 ( 
.A(n_4413),
.Y(n_4725)
);

NAND2x1p5_ASAP7_75t_L g4726 ( 
.A(n_4219),
.B(n_3743),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4410),
.B(n_3330),
.Y(n_4727)
);

BUFx2_ASAP7_75t_L g4728 ( 
.A(n_4463),
.Y(n_4728)
);

NOR2xp33_ASAP7_75t_SL g4729 ( 
.A(n_4219),
.B(n_4213),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4366),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_SL g4731 ( 
.A(n_4262),
.B(n_3630),
.Y(n_4731)
);

AND2x2_ASAP7_75t_L g4732 ( 
.A(n_4463),
.B(n_934),
.Y(n_4732)
);

INVx2_ASAP7_75t_L g4733 ( 
.A(n_4449),
.Y(n_4733)
);

AND3x1_ASAP7_75t_SL g4734 ( 
.A(n_4371),
.B(n_962),
.C(n_954),
.Y(n_4734)
);

INVx2_ASAP7_75t_SL g4735 ( 
.A(n_4459),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_L g4736 ( 
.A(n_4377),
.B(n_3332),
.Y(n_4736)
);

AND3x1_ASAP7_75t_SL g4737 ( 
.A(n_4395),
.B(n_979),
.C(n_977),
.Y(n_4737)
);

INVx2_ASAP7_75t_SL g4738 ( 
.A(n_4550),
.Y(n_4738)
);

INVx4_ASAP7_75t_L g4739 ( 
.A(n_4532),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4427),
.B(n_3332),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_4434),
.B(n_3419),
.Y(n_4741)
);

HB1xp67_ASAP7_75t_L g4742 ( 
.A(n_4309),
.Y(n_4742)
);

BUFx8_ASAP7_75t_L g4743 ( 
.A(n_4515),
.Y(n_4743)
);

INVx2_ASAP7_75t_L g4744 ( 
.A(n_4455),
.Y(n_4744)
);

AND2x4_ASAP7_75t_L g4745 ( 
.A(n_4442),
.B(n_3710),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_SL g4746 ( 
.A(n_4280),
.B(n_3630),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4349),
.B(n_3419),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4319),
.B(n_977),
.Y(n_4748)
);

INVx1_ASAP7_75t_SL g4749 ( 
.A(n_4495),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4253),
.B(n_3426),
.Y(n_4750)
);

AND2x4_ASAP7_75t_L g4751 ( 
.A(n_4458),
.B(n_3743),
.Y(n_4751)
);

INVx3_ASAP7_75t_L g4752 ( 
.A(n_4582),
.Y(n_4752)
);

NAND2xp5_ASAP7_75t_SL g4753 ( 
.A(n_4281),
.B(n_3630),
.Y(n_4753)
);

INVx1_ASAP7_75t_SL g4754 ( 
.A(n_4510),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4479),
.B(n_3426),
.Y(n_4755)
);

INVx2_ASAP7_75t_L g4756 ( 
.A(n_4468),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4437),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4461),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4478),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4494),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4445),
.B(n_3434),
.Y(n_4761)
);

O2A1O1Ixp33_ASAP7_75t_L g4762 ( 
.A1(n_4263),
.A2(n_1072),
.B(n_1084),
.C(n_1007),
.Y(n_4762)
);

INVx2_ASAP7_75t_L g4763 ( 
.A(n_4503),
.Y(n_4763)
);

BUFx2_ASAP7_75t_L g4764 ( 
.A(n_4322),
.Y(n_4764)
);

CKINVDCx20_ASAP7_75t_R g4765 ( 
.A(n_4513),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4527),
.B(n_3434),
.Y(n_4766)
);

BUFx4_ASAP7_75t_SL g4767 ( 
.A(n_4305),
.Y(n_4767)
);

INVx3_ASAP7_75t_SL g4768 ( 
.A(n_4364),
.Y(n_4768)
);

AND2x4_ASAP7_75t_L g4769 ( 
.A(n_4458),
.B(n_3743),
.Y(n_4769)
);

CKINVDCx5p33_ASAP7_75t_R g4770 ( 
.A(n_4544),
.Y(n_4770)
);

NOR2xp33_ASAP7_75t_L g4771 ( 
.A(n_4298),
.B(n_4164),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_4530),
.B(n_3435),
.Y(n_4772)
);

NOR3xp33_ASAP7_75t_L g4773 ( 
.A(n_4433),
.B(n_984),
.C(n_979),
.Y(n_4773)
);

INVx4_ASAP7_75t_L g4774 ( 
.A(n_4536),
.Y(n_4774)
);

INVx5_ASAP7_75t_L g4775 ( 
.A(n_4477),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4534),
.B(n_3435),
.Y(n_4776)
);

INVx6_ASAP7_75t_L g4777 ( 
.A(n_4219),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4537),
.B(n_3436),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4522),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4525),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_L g4781 ( 
.A(n_4480),
.B(n_3436),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_4488),
.B(n_3439),
.Y(n_4782)
);

INVx3_ASAP7_75t_L g4783 ( 
.A(n_4582),
.Y(n_4783)
);

INVx4_ASAP7_75t_L g4784 ( 
.A(n_4536),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4501),
.B(n_3439),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4506),
.Y(n_4786)
);

OR2x6_ASAP7_75t_L g4787 ( 
.A(n_4217),
.B(n_3743),
.Y(n_4787)
);

NAND2xp5_ASAP7_75t_L g4788 ( 
.A(n_4378),
.B(n_3135),
.Y(n_4788)
);

BUFx12f_ASAP7_75t_L g4789 ( 
.A(n_4382),
.Y(n_4789)
);

INVx2_ASAP7_75t_L g4790 ( 
.A(n_4560),
.Y(n_4790)
);

AND2x6_ASAP7_75t_L g4791 ( 
.A(n_4554),
.B(n_3773),
.Y(n_4791)
);

HB1xp67_ASAP7_75t_L g4792 ( 
.A(n_4311),
.Y(n_4792)
);

AOI22xp33_ASAP7_75t_SL g4793 ( 
.A1(n_4386),
.A2(n_988),
.B1(n_993),
.B2(n_984),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4256),
.B(n_3135),
.Y(n_4794)
);

BUFx6f_ASAP7_75t_L g4795 ( 
.A(n_4536),
.Y(n_4795)
);

AND2x2_ASAP7_75t_L g4796 ( 
.A(n_4555),
.B(n_988),
.Y(n_4796)
);

BUFx2_ASAP7_75t_L g4797 ( 
.A(n_4552),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4520),
.Y(n_4798)
);

INVx2_ASAP7_75t_SL g4799 ( 
.A(n_4541),
.Y(n_4799)
);

NAND2xp5_ASAP7_75t_SL g4800 ( 
.A(n_4363),
.B(n_3630),
.Y(n_4800)
);

INVx2_ASAP7_75t_SL g4801 ( 
.A(n_4541),
.Y(n_4801)
);

AND2x4_ASAP7_75t_L g4802 ( 
.A(n_4499),
.B(n_3773),
.Y(n_4802)
);

INVx3_ASAP7_75t_L g4803 ( 
.A(n_4507),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4551),
.Y(n_4804)
);

INVx2_ASAP7_75t_L g4805 ( 
.A(n_4556),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4585),
.Y(n_4806)
);

BUFx2_ASAP7_75t_L g4807 ( 
.A(n_4552),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4563),
.Y(n_4808)
);

BUFx6f_ASAP7_75t_L g4809 ( 
.A(n_4541),
.Y(n_4809)
);

INVx4_ASAP7_75t_L g4810 ( 
.A(n_4567),
.Y(n_4810)
);

INVx2_ASAP7_75t_L g4811 ( 
.A(n_4562),
.Y(n_4811)
);

INVx2_ASAP7_75t_L g4812 ( 
.A(n_4462),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_SL g4813 ( 
.A(n_4232),
.B(n_3630),
.Y(n_4813)
);

CKINVDCx5p33_ASAP7_75t_R g4814 ( 
.A(n_4409),
.Y(n_4814)
);

BUFx6f_ASAP7_75t_L g4815 ( 
.A(n_4567),
.Y(n_4815)
);

INVx3_ASAP7_75t_L g4816 ( 
.A(n_4507),
.Y(n_4816)
);

BUFx3_ASAP7_75t_L g4817 ( 
.A(n_4489),
.Y(n_4817)
);

BUFx3_ASAP7_75t_L g4818 ( 
.A(n_4489),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4498),
.Y(n_4819)
);

BUFx2_ASAP7_75t_L g4820 ( 
.A(n_4545),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4548),
.Y(n_4821)
);

NOR2xp33_ASAP7_75t_L g4822 ( 
.A(n_4292),
.B(n_961),
.Y(n_4822)
);

BUFx6f_ASAP7_75t_L g4823 ( 
.A(n_4567),
.Y(n_4823)
);

AND2x6_ASAP7_75t_L g4824 ( 
.A(n_4486),
.B(n_3773),
.Y(n_4824)
);

INVx5_ASAP7_75t_L g4825 ( 
.A(n_4477),
.Y(n_4825)
);

INVx2_ASAP7_75t_L g4826 ( 
.A(n_4472),
.Y(n_4826)
);

AND2x2_ASAP7_75t_SL g4827 ( 
.A(n_4487),
.B(n_3773),
.Y(n_4827)
);

BUFx6f_ASAP7_75t_L g4828 ( 
.A(n_4268),
.Y(n_4828)
);

NAND2xp5_ASAP7_75t_SL g4829 ( 
.A(n_4376),
.B(n_3645),
.Y(n_4829)
);

INVx3_ASAP7_75t_L g4830 ( 
.A(n_4509),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4589),
.Y(n_4831)
);

NAND2xp5_ASAP7_75t_SL g4832 ( 
.A(n_4347),
.B(n_3645),
.Y(n_4832)
);

INVx2_ASAP7_75t_L g4833 ( 
.A(n_4357),
.Y(n_4833)
);

INVx4_ASAP7_75t_L g4834 ( 
.A(n_4565),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4460),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4361),
.Y(n_4836)
);

AND2x2_ASAP7_75t_SL g4837 ( 
.A(n_4487),
.B(n_3789),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_L g4838 ( 
.A(n_4345),
.B(n_3137),
.Y(n_4838)
);

BUFx2_ASAP7_75t_L g4839 ( 
.A(n_4545),
.Y(n_4839)
);

BUFx6f_ASAP7_75t_L g4840 ( 
.A(n_4268),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4451),
.Y(n_4841)
);

BUFx2_ASAP7_75t_L g4842 ( 
.A(n_4549),
.Y(n_4842)
);

AND2x6_ASAP7_75t_L g4843 ( 
.A(n_4435),
.B(n_4222),
.Y(n_4843)
);

BUFx2_ASAP7_75t_L g4844 ( 
.A(n_4549),
.Y(n_4844)
);

AND2x2_ASAP7_75t_L g4845 ( 
.A(n_4490),
.B(n_993),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4452),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_L g4847 ( 
.A(n_4415),
.B(n_3137),
.Y(n_4847)
);

INVx2_ASAP7_75t_L g4848 ( 
.A(n_4509),
.Y(n_4848)
);

OR2x2_ASAP7_75t_L g4849 ( 
.A(n_4222),
.B(n_2574),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4598),
.B(n_3143),
.Y(n_4850)
);

INVx3_ASAP7_75t_L g4851 ( 
.A(n_4570),
.Y(n_4851)
);

NAND2xp5_ASAP7_75t_L g4852 ( 
.A(n_4600),
.B(n_3143),
.Y(n_4852)
);

INVx3_ASAP7_75t_L g4853 ( 
.A(n_4570),
.Y(n_4853)
);

HB1xp67_ASAP7_75t_L g4854 ( 
.A(n_4470),
.Y(n_4854)
);

NAND2xp5_ASAP7_75t_SL g4855 ( 
.A(n_4336),
.B(n_3645),
.Y(n_4855)
);

NOR2xp33_ASAP7_75t_L g4856 ( 
.A(n_4547),
.B(n_963),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4511),
.Y(n_4857)
);

AND2x4_ASAP7_75t_L g4858 ( 
.A(n_4446),
.B(n_4260),
.Y(n_4858)
);

HB1xp67_ASAP7_75t_L g4859 ( 
.A(n_4476),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4483),
.Y(n_4860)
);

NOR2xp33_ASAP7_75t_L g4861 ( 
.A(n_4257),
.B(n_4535),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4523),
.Y(n_4862)
);

NOR2xp33_ASAP7_75t_L g4863 ( 
.A(n_4257),
.B(n_964),
.Y(n_4863)
);

INVx2_ASAP7_75t_L g4864 ( 
.A(n_4538),
.Y(n_4864)
);

BUFx6f_ASAP7_75t_L g4865 ( 
.A(n_4413),
.Y(n_4865)
);

BUFx8_ASAP7_75t_L g4866 ( 
.A(n_4592),
.Y(n_4866)
);

INVx4_ASAP7_75t_L g4867 ( 
.A(n_4565),
.Y(n_4867)
);

BUFx6f_ASAP7_75t_L g4868 ( 
.A(n_4446),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4543),
.Y(n_4869)
);

AND2x2_ASAP7_75t_L g4870 ( 
.A(n_4385),
.B(n_994),
.Y(n_4870)
);

AND2x4_ASAP7_75t_L g4871 ( 
.A(n_4260),
.B(n_3789),
.Y(n_4871)
);

AND2x2_ASAP7_75t_L g4872 ( 
.A(n_4440),
.B(n_994),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_4467),
.B(n_3147),
.Y(n_4873)
);

INVx3_ASAP7_75t_L g4874 ( 
.A(n_4234),
.Y(n_4874)
);

CKINVDCx5p33_ASAP7_75t_R g4875 ( 
.A(n_4380),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_L g4876 ( 
.A(n_4474),
.B(n_3147),
.Y(n_4876)
);

AND2x2_ASAP7_75t_L g4877 ( 
.A(n_4368),
.B(n_1002),
.Y(n_4877)
);

OAI21xp5_ASAP7_75t_L g4878 ( 
.A1(n_4343),
.A2(n_2955),
.B(n_2953),
.Y(n_4878)
);

AND2x2_ASAP7_75t_L g4879 ( 
.A(n_4518),
.B(n_1002),
.Y(n_4879)
);

INVx2_ASAP7_75t_L g4880 ( 
.A(n_4569),
.Y(n_4880)
);

HB1xp67_ASAP7_75t_L g4881 ( 
.A(n_4360),
.Y(n_4881)
);

OR2x6_ASAP7_75t_L g4882 ( 
.A(n_4212),
.B(n_3789),
.Y(n_4882)
);

BUFx8_ASAP7_75t_L g4883 ( 
.A(n_4603),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_L g4884 ( 
.A(n_4475),
.B(n_3151),
.Y(n_4884)
);

CKINVDCx5p33_ASAP7_75t_R g4885 ( 
.A(n_4316),
.Y(n_4885)
);

OR2x2_ASAP7_75t_L g4886 ( 
.A(n_4348),
.B(n_4277),
.Y(n_4886)
);

NOR2xp33_ASAP7_75t_L g4887 ( 
.A(n_4238),
.B(n_965),
.Y(n_4887)
);

BUFx6f_ASAP7_75t_L g4888 ( 
.A(n_4234),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_SL g4889 ( 
.A(n_4313),
.B(n_3645),
.Y(n_4889)
);

INVx3_ASAP7_75t_L g4890 ( 
.A(n_4275),
.Y(n_4890)
);

NOR2xp67_ASAP7_75t_L g4891 ( 
.A(n_4401),
.B(n_3297),
.Y(n_4891)
);

HB1xp67_ASAP7_75t_L g4892 ( 
.A(n_4284),
.Y(n_4892)
);

BUFx3_ASAP7_75t_L g4893 ( 
.A(n_4439),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4447),
.B(n_3151),
.Y(n_4894)
);

INVx2_ASAP7_75t_L g4895 ( 
.A(n_4584),
.Y(n_4895)
);

A2O1A1Ixp33_ASAP7_75t_L g4896 ( 
.A1(n_4473),
.A2(n_1010),
.B(n_1013),
.C(n_1007),
.Y(n_4896)
);

INVx2_ASAP7_75t_L g4897 ( 
.A(n_4587),
.Y(n_4897)
);

INVx2_ASAP7_75t_L g4898 ( 
.A(n_4288),
.Y(n_4898)
);

INVx2_ASAP7_75t_L g4899 ( 
.A(n_4300),
.Y(n_4899)
);

INVx5_ASAP7_75t_L g4900 ( 
.A(n_4402),
.Y(n_4900)
);

BUFx2_ASAP7_75t_L g4901 ( 
.A(n_4595),
.Y(n_4901)
);

INVx2_ASAP7_75t_L g4902 ( 
.A(n_4302),
.Y(n_4902)
);

BUFx8_ASAP7_75t_L g4903 ( 
.A(n_4493),
.Y(n_4903)
);

INVx4_ASAP7_75t_L g4904 ( 
.A(n_4275),
.Y(n_4904)
);

AND2x2_ASAP7_75t_L g4905 ( 
.A(n_4310),
.B(n_1010),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4519),
.Y(n_4906)
);

AOI22xp5_ASAP7_75t_L g4907 ( 
.A1(n_4397),
.A2(n_969),
.B1(n_974),
.B2(n_973),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4586),
.Y(n_4908)
);

INVx2_ASAP7_75t_L g4909 ( 
.A(n_4223),
.Y(n_4909)
);

CKINVDCx5p33_ASAP7_75t_R g4910 ( 
.A(n_4425),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4252),
.Y(n_4911)
);

AND2x2_ASAP7_75t_L g4912 ( 
.A(n_4425),
.B(n_1013),
.Y(n_4912)
);

NAND2xp5_ASAP7_75t_L g4913 ( 
.A(n_4372),
.B(n_3645),
.Y(n_4913)
);

INVx2_ASAP7_75t_L g4914 ( 
.A(n_4408),
.Y(n_4914)
);

INVx2_ASAP7_75t_L g4915 ( 
.A(n_4399),
.Y(n_4915)
);

AND2x4_ASAP7_75t_L g4916 ( 
.A(n_4553),
.B(n_3789),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_L g4917 ( 
.A(n_4372),
.B(n_3672),
.Y(n_4917)
);

INVx2_ASAP7_75t_SL g4918 ( 
.A(n_4248),
.Y(n_4918)
);

CKINVDCx16_ASAP7_75t_R g4919 ( 
.A(n_4465),
.Y(n_4919)
);

NAND2xp5_ASAP7_75t_L g4920 ( 
.A(n_4273),
.B(n_3672),
.Y(n_4920)
);

BUFx12f_ASAP7_75t_L g4921 ( 
.A(n_4533),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_SL g4922 ( 
.A(n_4276),
.B(n_3672),
.Y(n_4922)
);

INVx2_ASAP7_75t_SL g4923 ( 
.A(n_4497),
.Y(n_4923)
);

CKINVDCx5p33_ASAP7_75t_R g4924 ( 
.A(n_4465),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4273),
.B(n_3767),
.Y(n_4925)
);

NOR2xp33_ASAP7_75t_L g4926 ( 
.A(n_4583),
.B(n_975),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_L g4927 ( 
.A(n_4247),
.B(n_4250),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_4412),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4333),
.B(n_3767),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_SL g4930 ( 
.A(n_4265),
.B(n_3767),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4249),
.B(n_3767),
.Y(n_4931)
);

INVxp67_ASAP7_75t_L g4932 ( 
.A(n_4516),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4436),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_L g4934 ( 
.A(n_4249),
.B(n_3767),
.Y(n_4934)
);

INVx2_ASAP7_75t_L g4935 ( 
.A(n_4590),
.Y(n_4935)
);

INVx2_ASAP7_75t_L g4936 ( 
.A(n_4514),
.Y(n_4936)
);

INVx2_ASAP7_75t_L g4937 ( 
.A(n_4329),
.Y(n_4937)
);

HB1xp67_ASAP7_75t_L g4938 ( 
.A(n_4374),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4573),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4573),
.Y(n_4940)
);

NOR2xp33_ASAP7_75t_R g4941 ( 
.A(n_4213),
.B(n_3810),
.Y(n_4941)
);

AOI22xp33_ASAP7_75t_L g4942 ( 
.A1(n_4529),
.A2(n_1019),
.B1(n_1020),
.B2(n_1015),
.Y(n_4942)
);

AND2x4_ASAP7_75t_L g4943 ( 
.A(n_4512),
.B(n_3810),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4578),
.Y(n_4944)
);

NOR2xp33_ASAP7_75t_L g4945 ( 
.A(n_4254),
.B(n_976),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4578),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4516),
.Y(n_4947)
);

NOR2xp33_ASAP7_75t_L g4948 ( 
.A(n_4469),
.B(n_978),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4344),
.B(n_3767),
.Y(n_4949)
);

AND2x2_ASAP7_75t_L g4950 ( 
.A(n_4342),
.B(n_1015),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4340),
.Y(n_4951)
);

BUFx3_ASAP7_75t_L g4952 ( 
.A(n_4334),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_4344),
.B(n_3297),
.Y(n_4953)
);

AOI21xp5_ASAP7_75t_L g4954 ( 
.A1(n_4216),
.A2(n_3175),
.B(n_3149),
.Y(n_4954)
);

BUFx12f_ASAP7_75t_L g4955 ( 
.A(n_4561),
.Y(n_4955)
);

NOR2xp67_ASAP7_75t_L g4956 ( 
.A(n_4574),
.B(n_3297),
.Y(n_4956)
);

BUFx6f_ASAP7_75t_L g4957 ( 
.A(n_4508),
.Y(n_4957)
);

AND2x6_ASAP7_75t_SL g4958 ( 
.A(n_4469),
.B(n_1019),
.Y(n_4958)
);

A2O1A1Ixp33_ASAP7_75t_L g4959 ( 
.A1(n_4411),
.A2(n_1022),
.B(n_1027),
.C(n_1020),
.Y(n_4959)
);

BUFx2_ASAP7_75t_L g4960 ( 
.A(n_4542),
.Y(n_4960)
);

INVx2_ASAP7_75t_SL g4961 ( 
.A(n_4418),
.Y(n_4961)
);

BUFx6f_ASAP7_75t_L g4962 ( 
.A(n_4557),
.Y(n_4962)
);

NOR2xp33_ASAP7_75t_L g4963 ( 
.A(n_4594),
.B(n_981),
.Y(n_4963)
);

AOI21xp5_ASAP7_75t_L g4964 ( 
.A1(n_4244),
.A2(n_4375),
.B(n_4373),
.Y(n_4964)
);

AOI22xp33_ASAP7_75t_L g4965 ( 
.A1(n_4390),
.A2(n_1027),
.B1(n_1030),
.B2(n_1022),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_L g4966 ( 
.A(n_4374),
.B(n_3316),
.Y(n_4966)
);

NAND3xp33_ASAP7_75t_L g4967 ( 
.A(n_4221),
.B(n_983),
.C(n_982),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4359),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4335),
.B(n_3316),
.Y(n_4969)
);

NOR2xp33_ASAP7_75t_L g4970 ( 
.A(n_4526),
.B(n_985),
.Y(n_4970)
);

AND3x1_ASAP7_75t_SL g4971 ( 
.A(n_4526),
.B(n_1039),
.C(n_1030),
.Y(n_4971)
);

INVx2_ASAP7_75t_L g4972 ( 
.A(n_4577),
.Y(n_4972)
);

AND2x6_ASAP7_75t_L g4973 ( 
.A(n_4221),
.B(n_3810),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4577),
.Y(n_4974)
);

NAND2xp5_ASAP7_75t_L g4975 ( 
.A(n_4335),
.B(n_3316),
.Y(n_4975)
);

INVx2_ASAP7_75t_L g4976 ( 
.A(n_4297),
.Y(n_4976)
);

NOR2xp33_ASAP7_75t_L g4977 ( 
.A(n_4293),
.B(n_986),
.Y(n_4977)
);

INVx1_ASAP7_75t_SL g4978 ( 
.A(n_4332),
.Y(n_4978)
);

INVx1_ASAP7_75t_L g4979 ( 
.A(n_4432),
.Y(n_4979)
);

BUFx8_ASAP7_75t_SL g4980 ( 
.A(n_4370),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_SL g4981 ( 
.A(n_4387),
.B(n_3810),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_SL g4982 ( 
.A(n_4297),
.B(n_3837),
.Y(n_4982)
);

INVx3_ASAP7_75t_L g4983 ( 
.A(n_4327),
.Y(n_4983)
);

AND2x2_ASAP7_75t_L g4984 ( 
.A(n_4270),
.B(n_1041),
.Y(n_4984)
);

AND2x2_ASAP7_75t_L g4985 ( 
.A(n_4270),
.B(n_1041),
.Y(n_4985)
);

BUFx2_ASAP7_75t_L g4986 ( 
.A(n_4539),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4354),
.B(n_3320),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4432),
.Y(n_4988)
);

BUFx3_ASAP7_75t_L g4989 ( 
.A(n_4384),
.Y(n_4989)
);

BUFx2_ASAP7_75t_L g4990 ( 
.A(n_4367),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4524),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_L g4992 ( 
.A(n_4369),
.B(n_4286),
.Y(n_4992)
);

AND2x4_ASAP7_75t_L g4993 ( 
.A(n_4328),
.B(n_3837),
.Y(n_4993)
);

NOR2xp33_ASAP7_75t_L g4994 ( 
.A(n_4338),
.B(n_987),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4531),
.Y(n_4995)
);

NAND2xp5_ASAP7_75t_L g4996 ( 
.A(n_4424),
.B(n_3320),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_SL g4997 ( 
.A(n_4267),
.B(n_3837),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4426),
.B(n_3320),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4540),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4546),
.Y(n_5000)
);

HB1xp67_ASAP7_75t_L g5001 ( 
.A(n_4224),
.Y(n_5001)
);

NAND2xp5_ASAP7_75t_L g5002 ( 
.A(n_4441),
.B(n_3837),
.Y(n_5002)
);

NAND2xp5_ASAP7_75t_L g5003 ( 
.A(n_4444),
.B(n_3333),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4450),
.B(n_3333),
.Y(n_5004)
);

HB1xp67_ASAP7_75t_SL g5005 ( 
.A(n_4384),
.Y(n_5005)
);

BUFx6f_ASAP7_75t_L g5006 ( 
.A(n_4571),
.Y(n_5006)
);

HB1xp67_ASAP7_75t_L g5007 ( 
.A(n_4392),
.Y(n_5007)
);

INVx2_ASAP7_75t_L g5008 ( 
.A(n_4398),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4492),
.B(n_3407),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4496),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4500),
.Y(n_5011)
);

AOI22xp33_ASAP7_75t_L g5012 ( 
.A1(n_4558),
.A2(n_1045),
.B1(n_1047),
.B2(n_1044),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_SL g5013 ( 
.A(n_4258),
.B(n_3250),
.Y(n_5013)
);

BUFx6f_ASAP7_75t_L g5014 ( 
.A(n_4572),
.Y(n_5014)
);

INVx3_ASAP7_75t_L g5015 ( 
.A(n_4575),
.Y(n_5015)
);

HB1xp67_ASAP7_75t_L g5016 ( 
.A(n_4224),
.Y(n_5016)
);

NOR2xp33_ASAP7_75t_L g5017 ( 
.A(n_4875),
.B(n_991),
.Y(n_5017)
);

OAI21x1_ASAP7_75t_L g5018 ( 
.A1(n_4964),
.A2(n_4274),
.B(n_4481),
.Y(n_5018)
);

BUFx6f_ASAP7_75t_L g5019 ( 
.A(n_4682),
.Y(n_5019)
);

OAI21x1_ASAP7_75t_L g5020 ( 
.A1(n_4964),
.A2(n_4484),
.B(n_4471),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_4606),
.Y(n_5021)
);

HB1xp67_ASAP7_75t_L g5022 ( 
.A(n_4617),
.Y(n_5022)
);

HB1xp67_ASAP7_75t_L g5023 ( 
.A(n_4617),
.Y(n_5023)
);

OR2x6_ASAP7_75t_L g5024 ( 
.A(n_4721),
.B(n_4304),
.Y(n_5024)
);

NOR2xp33_ASAP7_75t_L g5025 ( 
.A(n_4814),
.B(n_992),
.Y(n_5025)
);

NOR2xp33_ASAP7_75t_L g5026 ( 
.A(n_4609),
.B(n_995),
.Y(n_5026)
);

INVx2_ASAP7_75t_L g5027 ( 
.A(n_4805),
.Y(n_5027)
);

OAI22xp5_ASAP7_75t_L g5028 ( 
.A1(n_5005),
.A2(n_4602),
.B1(n_4566),
.B2(n_4339),
.Y(n_5028)
);

CKINVDCx5p33_ASAP7_75t_R g5029 ( 
.A(n_4665),
.Y(n_5029)
);

OR2x2_ASAP7_75t_L g5030 ( 
.A(n_4901),
.B(n_4504),
.Y(n_5030)
);

NAND2xp5_ASAP7_75t_L g5031 ( 
.A(n_4892),
.B(n_4307),
.Y(n_5031)
);

AOI21xp5_ASAP7_75t_L g5032 ( 
.A1(n_4646),
.A2(n_4323),
.B(n_4422),
.Y(n_5032)
);

NAND2xp5_ASAP7_75t_L g5033 ( 
.A(n_4749),
.B(n_4504),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_SL g5034 ( 
.A(n_4893),
.B(n_4294),
.Y(n_5034)
);

NOR2xp33_ASAP7_75t_L g5035 ( 
.A(n_4672),
.B(n_997),
.Y(n_5035)
);

OR2x6_ASAP7_75t_L g5036 ( 
.A(n_4721),
.B(n_4580),
.Y(n_5036)
);

BUFx6f_ASAP7_75t_SL g5037 ( 
.A(n_4625),
.Y(n_5037)
);

OAI21x1_ASAP7_75t_L g5038 ( 
.A1(n_4954),
.A2(n_4588),
.B(n_4581),
.Y(n_5038)
);

AOI22xp33_ASAP7_75t_L g5039 ( 
.A1(n_4955),
.A2(n_1045),
.B1(n_1047),
.B2(n_1044),
.Y(n_5039)
);

OAI21xp5_ASAP7_75t_L g5040 ( 
.A1(n_4977),
.A2(n_4337),
.B(n_4299),
.Y(n_5040)
);

O2A1O1Ixp33_ASAP7_75t_L g5041 ( 
.A1(n_4723),
.A2(n_1053),
.B(n_1056),
.C(n_1054),
.Y(n_5041)
);

INVx3_ASAP7_75t_L g5042 ( 
.A(n_4888),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_4749),
.B(n_4414),
.Y(n_5043)
);

INVxp67_ASAP7_75t_L g5044 ( 
.A(n_4656),
.Y(n_5044)
);

CKINVDCx8_ASAP7_75t_R g5045 ( 
.A(n_4687),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4630),
.Y(n_5046)
);

CKINVDCx5p33_ASAP7_75t_R g5047 ( 
.A(n_4692),
.Y(n_5047)
);

OR2x6_ASAP7_75t_SL g5048 ( 
.A(n_4910),
.B(n_998),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_4631),
.Y(n_5049)
);

AND2x2_ASAP7_75t_L g5050 ( 
.A(n_4623),
.B(n_4239),
.Y(n_5050)
);

AND2x4_ASAP7_75t_L g5051 ( 
.A(n_4858),
.B(n_4405),
.Y(n_5051)
);

NOR2xp33_ASAP7_75t_L g5052 ( 
.A(n_4771),
.B(n_4607),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4671),
.B(n_4406),
.Y(n_5053)
);

BUFx2_ASAP7_75t_L g5054 ( 
.A(n_4797),
.Y(n_5054)
);

INVx3_ASAP7_75t_L g5055 ( 
.A(n_4888),
.Y(n_5055)
);

BUFx10_ASAP7_75t_L g5056 ( 
.A(n_4770),
.Y(n_5056)
);

INVxp67_ASAP7_75t_L g5057 ( 
.A(n_4792),
.Y(n_5057)
);

INVx2_ASAP7_75t_L g5058 ( 
.A(n_4635),
.Y(n_5058)
);

INVx3_ASAP7_75t_L g5059 ( 
.A(n_4888),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_SL g5060 ( 
.A(n_4919),
.B(n_4314),
.Y(n_5060)
);

BUFx6f_ASAP7_75t_L g5061 ( 
.A(n_4682),
.Y(n_5061)
);

NOR2xp33_ASAP7_75t_L g5062 ( 
.A(n_4885),
.B(n_999),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4671),
.B(n_4591),
.Y(n_5063)
);

BUFx4f_ASAP7_75t_L g5064 ( 
.A(n_4828),
.Y(n_5064)
);

AND3x1_ASAP7_75t_SL g5065 ( 
.A(n_4698),
.B(n_1054),
.C(n_1053),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_4642),
.Y(n_5066)
);

AND2x2_ASAP7_75t_L g5067 ( 
.A(n_4854),
.B(n_4239),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_L g5068 ( 
.A(n_4636),
.B(n_4416),
.Y(n_5068)
);

BUFx6f_ASAP7_75t_L g5069 ( 
.A(n_4682),
.Y(n_5069)
);

A2O1A1Ixp33_ASAP7_75t_SL g5070 ( 
.A1(n_4948),
.A2(n_4240),
.B(n_1056),
.C(n_1071),
.Y(n_5070)
);

BUFx2_ASAP7_75t_L g5071 ( 
.A(n_4807),
.Y(n_5071)
);

AOI22xp5_ASAP7_75t_L g5072 ( 
.A1(n_4924),
.A2(n_1071),
.B1(n_1072),
.B2(n_1064),
.Y(n_5072)
);

BUFx3_ASAP7_75t_L g5073 ( 
.A(n_4789),
.Y(n_5073)
);

BUFx6f_ASAP7_75t_L g5074 ( 
.A(n_4701),
.Y(n_5074)
);

A2O1A1Ixp33_ASAP7_75t_L g5075 ( 
.A1(n_4945),
.A2(n_1077),
.B(n_1079),
.C(n_1064),
.Y(n_5075)
);

BUFx4_ASAP7_75t_SL g5076 ( 
.A(n_4677),
.Y(n_5076)
);

O2A1O1Ixp5_ASAP7_75t_L g5077 ( 
.A1(n_4714),
.A2(n_4599),
.B(n_4240),
.C(n_4403),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_4650),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_4659),
.Y(n_5079)
);

AOI22xp33_ASAP7_75t_L g5080 ( 
.A1(n_4989),
.A2(n_1079),
.B1(n_1080),
.B2(n_1077),
.Y(n_5080)
);

NOR2xp67_ASAP7_75t_L g5081 ( 
.A(n_4645),
.B(n_4394),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_4661),
.Y(n_5082)
);

BUFx4f_ASAP7_75t_SL g5083 ( 
.A(n_4673),
.Y(n_5083)
);

INVx4_ASAP7_75t_L g5084 ( 
.A(n_4828),
.Y(n_5084)
);

A2O1A1Ixp33_ASAP7_75t_L g5085 ( 
.A1(n_4963),
.A2(n_4960),
.B(n_4967),
.C(n_4926),
.Y(n_5085)
);

INVx2_ASAP7_75t_L g5086 ( 
.A(n_4681),
.Y(n_5086)
);

BUFx8_ASAP7_75t_L g5087 ( 
.A(n_4678),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_4636),
.B(n_4296),
.Y(n_5088)
);

NAND2x2_ASAP7_75t_L g5089 ( 
.A(n_4629),
.B(n_947),
.Y(n_5089)
);

INVx4_ASAP7_75t_L g5090 ( 
.A(n_4828),
.Y(n_5090)
);

BUFx12f_ASAP7_75t_L g5091 ( 
.A(n_4673),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_SL g5092 ( 
.A(n_4645),
.B(n_4324),
.Y(n_5092)
);

INVx3_ASAP7_75t_L g5093 ( 
.A(n_4868),
.Y(n_5093)
);

OAI22xp5_ASAP7_75t_L g5094 ( 
.A1(n_5005),
.A2(n_1084),
.B1(n_1085),
.B2(n_1080),
.Y(n_5094)
);

AOI22xp33_ASAP7_75t_L g5095 ( 
.A1(n_4921),
.A2(n_1092),
.B1(n_1095),
.B2(n_1085),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_4706),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_4707),
.Y(n_5097)
);

INVx2_ASAP7_75t_L g5098 ( 
.A(n_4709),
.Y(n_5098)
);

INVx2_ASAP7_75t_L g5099 ( 
.A(n_4711),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_4718),
.Y(n_5100)
);

AND2x2_ASAP7_75t_L g5101 ( 
.A(n_4859),
.B(n_4670),
.Y(n_5101)
);

CKINVDCx5p33_ASAP7_75t_R g5102 ( 
.A(n_4767),
.Y(n_5102)
);

NOR2xp67_ASAP7_75t_SL g5103 ( 
.A(n_4634),
.B(n_4576),
.Y(n_5103)
);

AND2x2_ASAP7_75t_L g5104 ( 
.A(n_4742),
.B(n_1092),
.Y(n_5104)
);

AOI22xp33_ASAP7_75t_L g5105 ( 
.A1(n_4856),
.A2(n_1100),
.B1(n_1103),
.B2(n_1095),
.Y(n_5105)
);

INVx1_ASAP7_75t_SL g5106 ( 
.A(n_4637),
.Y(n_5106)
);

INVx3_ASAP7_75t_L g5107 ( 
.A(n_4868),
.Y(n_5107)
);

AND2x2_ASAP7_75t_L g5108 ( 
.A(n_4754),
.B(n_1100),
.Y(n_5108)
);

AND2x4_ASAP7_75t_L g5109 ( 
.A(n_4858),
.B(n_4383),
.Y(n_5109)
);

AND2x6_ASAP7_75t_L g5110 ( 
.A(n_4957),
.B(n_3250),
.Y(n_5110)
);

INVx2_ASAP7_75t_L g5111 ( 
.A(n_4722),
.Y(n_5111)
);

INVxp67_ASAP7_75t_L g5112 ( 
.A(n_4764),
.Y(n_5112)
);

NAND2xp5_ASAP7_75t_L g5113 ( 
.A(n_4898),
.B(n_4326),
.Y(n_5113)
);

A2O1A1Ixp33_ASAP7_75t_L g5114 ( 
.A1(n_4986),
.A2(n_1116),
.B(n_1117),
.C(n_1103),
.Y(n_5114)
);

NAND2xp5_ASAP7_75t_SL g5115 ( 
.A(n_4645),
.B(n_4398),
.Y(n_5115)
);

AOI22xp5_ASAP7_75t_L g5116 ( 
.A1(n_4714),
.A2(n_1117),
.B1(n_1118),
.B2(n_1116),
.Y(n_5116)
);

INVx2_ASAP7_75t_L g5117 ( 
.A(n_4724),
.Y(n_5117)
);

OAI22xp33_ASAP7_75t_L g5118 ( 
.A1(n_4618),
.A2(n_1121),
.B1(n_1122),
.B2(n_1118),
.Y(n_5118)
);

BUFx2_ASAP7_75t_L g5119 ( 
.A(n_4667),
.Y(n_5119)
);

AND2x4_ASAP7_75t_L g5120 ( 
.A(n_4697),
.B(n_4564),
.Y(n_5120)
);

NOR2xp33_ASAP7_75t_L g5121 ( 
.A(n_4822),
.B(n_1000),
.Y(n_5121)
);

OAI22xp5_ASAP7_75t_L g5122 ( 
.A1(n_4793),
.A2(n_1122),
.B1(n_1124),
.B2(n_1121),
.Y(n_5122)
);

INVx3_ASAP7_75t_L g5123 ( 
.A(n_4868),
.Y(n_5123)
);

NOR2x1_ASAP7_75t_R g5124 ( 
.A(n_4697),
.B(n_1003),
.Y(n_5124)
);

HB1xp67_ASAP7_75t_L g5125 ( 
.A(n_4637),
.Y(n_5125)
);

INVx2_ASAP7_75t_L g5126 ( 
.A(n_4730),
.Y(n_5126)
);

AND2x2_ASAP7_75t_L g5127 ( 
.A(n_4754),
.B(n_1124),
.Y(n_5127)
);

BUFx2_ASAP7_75t_L g5128 ( 
.A(n_4604),
.Y(n_5128)
);

O2A1O1Ixp33_ASAP7_75t_L g5129 ( 
.A1(n_4723),
.A2(n_4698),
.B(n_4959),
.C(n_4896),
.Y(n_5129)
);

INVx1_ASAP7_75t_L g5130 ( 
.A(n_4757),
.Y(n_5130)
);

BUFx12f_ASAP7_75t_L g5131 ( 
.A(n_4866),
.Y(n_5131)
);

INVx4_ASAP7_75t_L g5132 ( 
.A(n_4840),
.Y(n_5132)
);

BUFx3_ASAP7_75t_L g5133 ( 
.A(n_4688),
.Y(n_5133)
);

INVx4_ASAP7_75t_L g5134 ( 
.A(n_4840),
.Y(n_5134)
);

OA21x2_ASAP7_75t_L g5135 ( 
.A1(n_4928),
.A2(n_4430),
.B(n_4568),
.Y(n_5135)
);

CKINVDCx5p33_ASAP7_75t_R g5136 ( 
.A(n_4767),
.Y(n_5136)
);

NAND2xp5_ASAP7_75t_L g5137 ( 
.A(n_4683),
.B(n_4430),
.Y(n_5137)
);

BUFx4f_ASAP7_75t_L g5138 ( 
.A(n_4840),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_4758),
.Y(n_5139)
);

INVx5_ASAP7_75t_L g5140 ( 
.A(n_4618),
.Y(n_5140)
);

AOI21xp5_ASAP7_75t_L g5141 ( 
.A1(n_4649),
.A2(n_4466),
.B(n_3182),
.Y(n_5141)
);

AOI22xp33_ASAP7_75t_L g5142 ( 
.A1(n_4970),
.A2(n_1131),
.B1(n_1136),
.B2(n_1128),
.Y(n_5142)
);

INVx2_ASAP7_75t_L g5143 ( 
.A(n_4759),
.Y(n_5143)
);

BUFx2_ASAP7_75t_L g5144 ( 
.A(n_4728),
.Y(n_5144)
);

INVx3_ASAP7_75t_L g5145 ( 
.A(n_4874),
.Y(n_5145)
);

OAI22xp5_ASAP7_75t_L g5146 ( 
.A1(n_4793),
.A2(n_1131),
.B1(n_1136),
.B2(n_1128),
.Y(n_5146)
);

AOI222xp33_ASAP7_75t_L g5147 ( 
.A1(n_4872),
.A2(n_1152),
.B1(n_1143),
.B2(n_1156),
.C1(n_1147),
.C2(n_1138),
.Y(n_5147)
);

INVx2_ASAP7_75t_L g5148 ( 
.A(n_4786),
.Y(n_5148)
);

AND2x2_ASAP7_75t_L g5149 ( 
.A(n_4611),
.B(n_1138),
.Y(n_5149)
);

AOI21xp5_ASAP7_75t_L g5150 ( 
.A1(n_4649),
.A2(n_3182),
.B(n_3175),
.Y(n_5150)
);

NAND2xp5_ASAP7_75t_L g5151 ( 
.A(n_4683),
.B(n_1143),
.Y(n_5151)
);

AND2x4_ASAP7_75t_L g5152 ( 
.A(n_4697),
.B(n_3250),
.Y(n_5152)
);

INVx2_ASAP7_75t_L g5153 ( 
.A(n_4798),
.Y(n_5153)
);

AND2x4_ASAP7_75t_L g5154 ( 
.A(n_4697),
.B(n_3261),
.Y(n_5154)
);

NOR2xp33_ASAP7_75t_L g5155 ( 
.A(n_4861),
.B(n_1004),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_SL g5156 ( 
.A(n_4775),
.B(n_1450),
.Y(n_5156)
);

INVx2_ASAP7_75t_L g5157 ( 
.A(n_4804),
.Y(n_5157)
);

AND2x2_ASAP7_75t_L g5158 ( 
.A(n_4833),
.B(n_4648),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_4947),
.B(n_1147),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_4806),
.Y(n_5160)
);

BUFx2_ASAP7_75t_L g5161 ( 
.A(n_4624),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_4808),
.Y(n_5162)
);

NOR2xp33_ASAP7_75t_L g5163 ( 
.A(n_4719),
.B(n_1005),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_4951),
.Y(n_5164)
);

OR2x2_ASAP7_75t_L g5165 ( 
.A(n_4886),
.B(n_1511),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_4911),
.Y(n_5166)
);

OAI321xp33_ASAP7_75t_L g5167 ( 
.A1(n_4618),
.A2(n_1160),
.A3(n_1156),
.B1(n_1161),
.B2(n_1158),
.C(n_1152),
.Y(n_5167)
);

INVx4_ASAP7_75t_L g5168 ( 
.A(n_4640),
.Y(n_5168)
);

BUFx3_ASAP7_75t_L g5169 ( 
.A(n_4768),
.Y(n_5169)
);

AOI21xp5_ASAP7_75t_L g5170 ( 
.A1(n_4627),
.A2(n_3223),
.B(n_3182),
.Y(n_5170)
);

INVx2_ASAP7_75t_L g5171 ( 
.A(n_4605),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_4937),
.Y(n_5172)
);

INVx2_ASAP7_75t_L g5173 ( 
.A(n_4614),
.Y(n_5173)
);

NOR2xp33_ASAP7_75t_L g5174 ( 
.A(n_4719),
.B(n_1006),
.Y(n_5174)
);

A2O1A1Ixp33_ASAP7_75t_L g5175 ( 
.A1(n_4887),
.A2(n_1160),
.B(n_1161),
.C(n_1158),
.Y(n_5175)
);

INVx2_ASAP7_75t_L g5176 ( 
.A(n_4620),
.Y(n_5176)
);

BUFx6f_ASAP7_75t_L g5177 ( 
.A(n_4701),
.Y(n_5177)
);

INVx3_ASAP7_75t_L g5178 ( 
.A(n_4874),
.Y(n_5178)
);

O2A1O1Ixp33_ASAP7_75t_L g5179 ( 
.A1(n_4870),
.A2(n_1162),
.B(n_1167),
.C(n_1166),
.Y(n_5179)
);

HB1xp67_ASAP7_75t_L g5180 ( 
.A(n_4648),
.Y(n_5180)
);

AOI22xp33_ASAP7_75t_L g5181 ( 
.A1(n_4903),
.A2(n_1166),
.B1(n_1167),
.B2(n_1162),
.Y(n_5181)
);

NOR2xp33_ASAP7_75t_L g5182 ( 
.A(n_4639),
.B(n_4863),
.Y(n_5182)
);

OAI22xp5_ASAP7_75t_L g5183 ( 
.A1(n_4628),
.A2(n_1169),
.B1(n_1170),
.B2(n_1168),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_4908),
.Y(n_5184)
);

BUFx6f_ASAP7_75t_SL g5185 ( 
.A(n_4625),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_4899),
.B(n_1011),
.Y(n_5186)
);

NAND2xp5_ASAP7_75t_L g5187 ( 
.A(n_4902),
.B(n_4684),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_4831),
.Y(n_5188)
);

AOI22xp5_ASAP7_75t_L g5189 ( 
.A1(n_4903),
.A2(n_1169),
.B1(n_1170),
.B2(n_1168),
.Y(n_5189)
);

O2A1O1Ixp33_ASAP7_75t_L g5190 ( 
.A1(n_4773),
.A2(n_1181),
.B(n_1190),
.C(n_1188),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_L g5191 ( 
.A(n_4684),
.B(n_1012),
.Y(n_5191)
);

BUFx6f_ASAP7_75t_L g5192 ( 
.A(n_4701),
.Y(n_5192)
);

INVx2_ASAP7_75t_L g5193 ( 
.A(n_4641),
.Y(n_5193)
);

NAND2xp5_ASAP7_75t_SL g5194 ( 
.A(n_4775),
.B(n_1511),
.Y(n_5194)
);

BUFx2_ASAP7_75t_SL g5195 ( 
.A(n_4621),
.Y(n_5195)
);

NAND2xp5_ASAP7_75t_L g5196 ( 
.A(n_4835),
.B(n_1014),
.Y(n_5196)
);

AOI22xp33_ASAP7_75t_L g5197 ( 
.A1(n_4990),
.A2(n_1188),
.B1(n_1190),
.B2(n_1181),
.Y(n_5197)
);

BUFx3_ASAP7_75t_L g5198 ( 
.A(n_4610),
.Y(n_5198)
);

INVx2_ASAP7_75t_L g5199 ( 
.A(n_4653),
.Y(n_5199)
);

INVx2_ASAP7_75t_L g5200 ( 
.A(n_4663),
.Y(n_5200)
);

AOI21xp33_ASAP7_75t_L g5201 ( 
.A1(n_4984),
.A2(n_2574),
.B(n_1205),
.Y(n_5201)
);

AO21x2_ASAP7_75t_L g5202 ( 
.A1(n_5013),
.A2(n_2534),
.B(n_2533),
.Y(n_5202)
);

AND2x4_ASAP7_75t_L g5203 ( 
.A(n_4775),
.B(n_3261),
.Y(n_5203)
);

CKINVDCx5p33_ASAP7_75t_R g5204 ( 
.A(n_4866),
.Y(n_5204)
);

NAND2xp5_ASAP7_75t_L g5205 ( 
.A(n_4915),
.B(n_1016),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4821),
.Y(n_5206)
);

NOR3xp33_ASAP7_75t_L g5207 ( 
.A(n_4994),
.B(n_1205),
.C(n_1193),
.Y(n_5207)
);

AOI221xp5_ASAP7_75t_L g5208 ( 
.A1(n_4720),
.A2(n_1018),
.B1(n_1023),
.B2(n_1021),
.C(n_1017),
.Y(n_5208)
);

BUFx2_ASAP7_75t_L g5209 ( 
.A(n_4633),
.Y(n_5209)
);

NAND2xp5_ASAP7_75t_L g5210 ( 
.A(n_4690),
.B(n_1024),
.Y(n_5210)
);

NAND2xp5_ASAP7_75t_L g5211 ( 
.A(n_4914),
.B(n_1026),
.Y(n_5211)
);

AOI22xp5_ASAP7_75t_L g5212 ( 
.A1(n_4773),
.A2(n_1193),
.B1(n_1029),
.B2(n_1032),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_4909),
.Y(n_5213)
);

AOI21xp5_ASAP7_75t_L g5214 ( 
.A1(n_4627),
.A2(n_3258),
.B(n_3223),
.Y(n_5214)
);

BUFx6f_ASAP7_75t_L g5215 ( 
.A(n_4795),
.Y(n_5215)
);

INVx2_ASAP7_75t_L g5216 ( 
.A(n_4674),
.Y(n_5216)
);

OR2x6_ASAP7_75t_L g5217 ( 
.A(n_4721),
.B(n_3261),
.Y(n_5217)
);

AO31x2_ASAP7_75t_L g5218 ( 
.A1(n_4933),
.A2(n_2535),
.A3(n_2557),
.B(n_2534),
.Y(n_5218)
);

CKINVDCx20_ASAP7_75t_R g5219 ( 
.A(n_4883),
.Y(n_5219)
);

A2O1A1Ixp33_ASAP7_75t_L g5220 ( 
.A1(n_4762),
.A2(n_1031),
.B(n_1035),
.C(n_1033),
.Y(n_5220)
);

BUFx6f_ASAP7_75t_L g5221 ( 
.A(n_4795),
.Y(n_5221)
);

A2O1A1Ixp33_ASAP7_75t_L g5222 ( 
.A1(n_4762),
.A2(n_1036),
.B(n_1050),
.C(n_1043),
.Y(n_5222)
);

BUFx6f_ASAP7_75t_L g5223 ( 
.A(n_4795),
.Y(n_5223)
);

INVx6_ASAP7_75t_L g5224 ( 
.A(n_4883),
.Y(n_5224)
);

O2A1O1Ixp33_ASAP7_75t_L g5225 ( 
.A1(n_4720),
.A2(n_2958),
.B(n_2955),
.C(n_2956),
.Y(n_5225)
);

NOR2xp33_ASAP7_75t_L g5226 ( 
.A(n_4765),
.B(n_1051),
.Y(n_5226)
);

AND2x4_ASAP7_75t_SL g5227 ( 
.A(n_4865),
.B(n_3261),
.Y(n_5227)
);

INVx3_ASAP7_75t_L g5228 ( 
.A(n_4638),
.Y(n_5228)
);

BUFx2_ASAP7_75t_L g5229 ( 
.A(n_4613),
.Y(n_5229)
);

A2O1A1Ixp33_ASAP7_75t_L g5230 ( 
.A1(n_4985),
.A2(n_1055),
.B(n_1058),
.C(n_1057),
.Y(n_5230)
);

OR2x2_ASAP7_75t_L g5231 ( 
.A(n_4913),
.B(n_1511),
.Y(n_5231)
);

INVx5_ASAP7_75t_L g5232 ( 
.A(n_4980),
.Y(n_5232)
);

OAI21xp5_ASAP7_75t_L g5233 ( 
.A1(n_5012),
.A2(n_2959),
.B(n_2956),
.Y(n_5233)
);

NAND2xp5_ASAP7_75t_L g5234 ( 
.A(n_4811),
.B(n_1059),
.Y(n_5234)
);

NOR2xp33_ASAP7_75t_L g5235 ( 
.A(n_4865),
.B(n_1060),
.Y(n_5235)
);

NOR2xp33_ASAP7_75t_L g5236 ( 
.A(n_4865),
.B(n_4735),
.Y(n_5236)
);

BUFx3_ASAP7_75t_L g5237 ( 
.A(n_4615),
.Y(n_5237)
);

A2O1A1Ixp33_ASAP7_75t_L g5238 ( 
.A1(n_4932),
.A2(n_1061),
.B(n_1063),
.C(n_1062),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_4976),
.Y(n_5239)
);

O2A1O1Ixp5_ASAP7_75t_SL g5240 ( 
.A1(n_4968),
.A2(n_2557),
.B(n_2535),
.C(n_2959),
.Y(n_5240)
);

AOI21xp5_ASAP7_75t_L g5241 ( 
.A1(n_4643),
.A2(n_3258),
.B(n_3223),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_4680),
.Y(n_5242)
);

INVx2_ASAP7_75t_SL g5243 ( 
.A(n_4809),
.Y(n_5243)
);

OAI22xp5_ASAP7_75t_L g5244 ( 
.A1(n_4775),
.A2(n_1066),
.B1(n_1074),
.B2(n_1068),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_4691),
.Y(n_5245)
);

BUFx12f_ASAP7_75t_L g5246 ( 
.A(n_4743),
.Y(n_5246)
);

AOI22xp33_ASAP7_75t_L g5247 ( 
.A1(n_4906),
.A2(n_1076),
.B1(n_1081),
.B2(n_1078),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_4704),
.Y(n_5248)
);

NOR2xp33_ASAP7_75t_SL g5249 ( 
.A(n_4825),
.B(n_3286),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_4812),
.B(n_1086),
.Y(n_5250)
);

INVx2_ASAP7_75t_L g5251 ( 
.A(n_4713),
.Y(n_5251)
);

INVx6_ASAP7_75t_L g5252 ( 
.A(n_4666),
.Y(n_5252)
);

AND2x4_ASAP7_75t_L g5253 ( 
.A(n_4825),
.B(n_3261),
.Y(n_5253)
);

INVx3_ASAP7_75t_L g5254 ( 
.A(n_4638),
.Y(n_5254)
);

INVx1_ASAP7_75t_SL g5255 ( 
.A(n_4820),
.Y(n_5255)
);

BUFx2_ASAP7_75t_L g5256 ( 
.A(n_4839),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_4716),
.Y(n_5257)
);

INVx2_ASAP7_75t_SL g5258 ( 
.A(n_4809),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_L g5259 ( 
.A(n_4932),
.B(n_1511),
.Y(n_5259)
);

INVx1_ASAP7_75t_L g5260 ( 
.A(n_4717),
.Y(n_5260)
);

INVx2_ASAP7_75t_L g5261 ( 
.A(n_4733),
.Y(n_5261)
);

INVx4_ASAP7_75t_L g5262 ( 
.A(n_4640),
.Y(n_5262)
);

BUFx6f_ASAP7_75t_L g5263 ( 
.A(n_4809),
.Y(n_5263)
);

INVx2_ASAP7_75t_L g5264 ( 
.A(n_4744),
.Y(n_5264)
);

BUFx6f_ASAP7_75t_L g5265 ( 
.A(n_4815),
.Y(n_5265)
);

AOI22xp5_ASAP7_75t_L g5266 ( 
.A1(n_4912),
.A2(n_1088),
.B1(n_1091),
.B2(n_1089),
.Y(n_5266)
);

AOI22xp5_ASAP7_75t_L g5267 ( 
.A1(n_4950),
.A2(n_1093),
.B1(n_1096),
.B2(n_1094),
.Y(n_5267)
);

AOI22xp33_ASAP7_75t_L g5268 ( 
.A1(n_4957),
.A2(n_1097),
.B1(n_1101),
.B2(n_1099),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_4756),
.Y(n_5269)
);

NOR2xp67_ASAP7_75t_L g5270 ( 
.A(n_4825),
.B(n_4927),
.Y(n_5270)
);

AOI21xp5_ASAP7_75t_L g5271 ( 
.A1(n_4643),
.A2(n_3294),
.B(n_3258),
.Y(n_5271)
);

INVx4_ASAP7_75t_L g5272 ( 
.A(n_4647),
.Y(n_5272)
);

BUFx6f_ASAP7_75t_L g5273 ( 
.A(n_4815),
.Y(n_5273)
);

INVx2_ASAP7_75t_L g5274 ( 
.A(n_4760),
.Y(n_5274)
);

INVx2_ASAP7_75t_L g5275 ( 
.A(n_4763),
.Y(n_5275)
);

AND2x4_ASAP7_75t_L g5276 ( 
.A(n_4825),
.B(n_3279),
.Y(n_5276)
);

OAI22xp5_ASAP7_75t_L g5277 ( 
.A1(n_4965),
.A2(n_1102),
.B1(n_1106),
.B2(n_1104),
.Y(n_5277)
);

AOI21xp5_ASAP7_75t_L g5278 ( 
.A1(n_4626),
.A2(n_3389),
.B(n_3294),
.Y(n_5278)
);

INVx3_ASAP7_75t_L g5279 ( 
.A(n_4803),
.Y(n_5279)
);

AOI22xp5_ASAP7_75t_L g5280 ( 
.A1(n_4612),
.A2(n_1109),
.B1(n_1112),
.B2(n_1110),
.Y(n_5280)
);

INVxp67_ASAP7_75t_L g5281 ( 
.A(n_4881),
.Y(n_5281)
);

AOI21xp5_ASAP7_75t_L g5282 ( 
.A1(n_4626),
.A2(n_3389),
.B(n_3294),
.Y(n_5282)
);

NAND2xp5_ASAP7_75t_L g5283 ( 
.A(n_4651),
.B(n_1678),
.Y(n_5283)
);

INVx2_ASAP7_75t_L g5284 ( 
.A(n_4779),
.Y(n_5284)
);

NAND2xp5_ASAP7_75t_SL g5285 ( 
.A(n_4904),
.B(n_1678),
.Y(n_5285)
);

INVx3_ASAP7_75t_L g5286 ( 
.A(n_4803),
.Y(n_5286)
);

BUFx4f_ASAP7_75t_SL g5287 ( 
.A(n_4743),
.Y(n_5287)
);

BUFx3_ASAP7_75t_L g5288 ( 
.A(n_4662),
.Y(n_5288)
);

OR2x6_ASAP7_75t_L g5289 ( 
.A(n_4676),
.B(n_3279),
.Y(n_5289)
);

INVx4_ASAP7_75t_L g5290 ( 
.A(n_4647),
.Y(n_5290)
);

A2O1A1Ixp33_ASAP7_75t_L g5291 ( 
.A1(n_4729),
.A2(n_1113),
.B(n_1115),
.C(n_1114),
.Y(n_5291)
);

INVx2_ASAP7_75t_L g5292 ( 
.A(n_4780),
.Y(n_5292)
);

OR2x6_ASAP7_75t_SL g5293 ( 
.A(n_4927),
.B(n_4651),
.Y(n_5293)
);

INVx5_ASAP7_75t_L g5294 ( 
.A(n_5006),
.Y(n_5294)
);

A2O1A1Ixp33_ASAP7_75t_L g5295 ( 
.A1(n_4729),
.A2(n_1119),
.B(n_1125),
.C(n_1120),
.Y(n_5295)
);

AND2x2_ASAP7_75t_L g5296 ( 
.A(n_4957),
.B(n_12),
.Y(n_5296)
);

INVx3_ASAP7_75t_L g5297 ( 
.A(n_4816),
.Y(n_5297)
);

INVx2_ASAP7_75t_L g5298 ( 
.A(n_4790),
.Y(n_5298)
);

NAND2xp5_ASAP7_75t_L g5299 ( 
.A(n_4836),
.B(n_1678),
.Y(n_5299)
);

INVxp67_ASAP7_75t_SL g5300 ( 
.A(n_4616),
.Y(n_5300)
);

NAND2xp5_ASAP7_75t_L g5301 ( 
.A(n_4826),
.B(n_1127),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_4860),
.Y(n_5302)
);

AND2x2_ASAP7_75t_L g5303 ( 
.A(n_4845),
.B(n_14),
.Y(n_5303)
);

AND2x4_ASAP7_75t_L g5304 ( 
.A(n_4890),
.B(n_4923),
.Y(n_5304)
);

INVx2_ASAP7_75t_L g5305 ( 
.A(n_4848),
.Y(n_5305)
);

INVx1_ASAP7_75t_L g5306 ( 
.A(n_4841),
.Y(n_5306)
);

BUFx2_ASAP7_75t_L g5307 ( 
.A(n_4842),
.Y(n_5307)
);

INVx2_ASAP7_75t_L g5308 ( 
.A(n_4705),
.Y(n_5308)
);

AND2x2_ASAP7_75t_L g5309 ( 
.A(n_4644),
.B(n_15),
.Y(n_5309)
);

NAND2xp5_ASAP7_75t_L g5310 ( 
.A(n_4846),
.B(n_1130),
.Y(n_5310)
);

NAND2x1_ASAP7_75t_L g5311 ( 
.A(n_4904),
.B(n_3389),
.Y(n_5311)
);

INVx1_ASAP7_75t_L g5312 ( 
.A(n_4935),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_4961),
.Y(n_5313)
);

NOR2xp33_ASAP7_75t_L g5314 ( 
.A(n_4958),
.B(n_1132),
.Y(n_5314)
);

OAI22xp5_ASAP7_75t_L g5315 ( 
.A1(n_4660),
.A2(n_1133),
.B1(n_1140),
.B2(n_1134),
.Y(n_5315)
);

BUFx12f_ASAP7_75t_L g5316 ( 
.A(n_4666),
.Y(n_5316)
);

AOI22xp5_ASAP7_75t_L g5317 ( 
.A1(n_4734),
.A2(n_1142),
.B1(n_1145),
.B2(n_1144),
.Y(n_5317)
);

AOI21xp5_ASAP7_75t_L g5318 ( 
.A1(n_4668),
.A2(n_3433),
.B(n_3366),
.Y(n_5318)
);

AND2x2_ASAP7_75t_L g5319 ( 
.A(n_4962),
.B(n_17),
.Y(n_5319)
);

BUFx2_ASAP7_75t_L g5320 ( 
.A(n_4844),
.Y(n_5320)
);

CKINVDCx20_ASAP7_75t_R g5321 ( 
.A(n_4817),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_4788),
.Y(n_5322)
);

NAND2xp5_ASAP7_75t_L g5323 ( 
.A(n_4819),
.B(n_1146),
.Y(n_5323)
);

OR2x6_ASAP7_75t_L g5324 ( 
.A(n_4676),
.B(n_3279),
.Y(n_5324)
);

AOI21xp5_ASAP7_75t_L g5325 ( 
.A1(n_4668),
.A2(n_3433),
.B(n_3366),
.Y(n_5325)
);

O2A1O1Ixp33_ASAP7_75t_L g5326 ( 
.A1(n_4694),
.A2(n_2954),
.B(n_2659),
.C(n_2669),
.Y(n_5326)
);

BUFx6f_ASAP7_75t_L g5327 ( 
.A(n_4815),
.Y(n_5327)
);

OAI21xp5_ASAP7_75t_L g5328 ( 
.A1(n_4700),
.A2(n_4878),
.B(n_4813),
.Y(n_5328)
);

BUFx6f_ASAP7_75t_L g5329 ( 
.A(n_4823),
.Y(n_5329)
);

AOI21xp5_ASAP7_75t_L g5330 ( 
.A1(n_4900),
.A2(n_3433),
.B(n_3366),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_4788),
.Y(n_5331)
);

INVx1_ASAP7_75t_SL g5332 ( 
.A(n_4952),
.Y(n_5332)
);

BUFx2_ASAP7_75t_L g5333 ( 
.A(n_4752),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_5007),
.Y(n_5334)
);

NAND2xp5_ASAP7_75t_L g5335 ( 
.A(n_4608),
.B(n_1148),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_4972),
.Y(n_5336)
);

INVx1_ASAP7_75t_SL g5337 ( 
.A(n_4978),
.Y(n_5337)
);

INVx2_ASAP7_75t_SL g5338 ( 
.A(n_4823),
.Y(n_5338)
);

NAND2xp5_ASAP7_75t_L g5339 ( 
.A(n_4608),
.B(n_1149),
.Y(n_5339)
);

CKINVDCx20_ASAP7_75t_R g5340 ( 
.A(n_4818),
.Y(n_5340)
);

INVx2_ASAP7_75t_SL g5341 ( 
.A(n_4823),
.Y(n_5341)
);

AND2x4_ASAP7_75t_L g5342 ( 
.A(n_4890),
.B(n_3279),
.Y(n_5342)
);

AND2x2_ASAP7_75t_L g5343 ( 
.A(n_4962),
.B(n_4654),
.Y(n_5343)
);

HB1xp67_ASAP7_75t_L g5344 ( 
.A(n_4962),
.Y(n_5344)
);

BUFx6f_ASAP7_75t_L g5345 ( 
.A(n_4655),
.Y(n_5345)
);

AND2x2_ASAP7_75t_L g5346 ( 
.A(n_4699),
.B(n_18),
.Y(n_5346)
);

INVx2_ASAP7_75t_L g5347 ( 
.A(n_4816),
.Y(n_5347)
);

NAND2xp5_ASAP7_75t_L g5348 ( 
.A(n_4622),
.B(n_1153),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_4974),
.Y(n_5349)
);

AOI21x1_ASAP7_75t_L g5350 ( 
.A1(n_4997),
.A2(n_2574),
.B(n_2947),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_4703),
.Y(n_5351)
);

OAI22xp5_ASAP7_75t_L g5352 ( 
.A1(n_4938),
.A2(n_1154),
.B1(n_1157),
.B2(n_1155),
.Y(n_5352)
);

NAND2xp5_ASAP7_75t_L g5353 ( 
.A(n_4622),
.B(n_1159),
.Y(n_5353)
);

OAI21xp33_ASAP7_75t_L g5354 ( 
.A1(n_4652),
.A2(n_1165),
.B(n_1164),
.Y(n_5354)
);

AOI22xp33_ASAP7_75t_L g5355 ( 
.A1(n_4843),
.A2(n_1171),
.B1(n_1178),
.B2(n_1172),
.Y(n_5355)
);

A2O1A1Ixp33_ASAP7_75t_L g5356 ( 
.A1(n_4907),
.A2(n_1179),
.B(n_1184),
.C(n_1180),
.Y(n_5356)
);

INVx4_ASAP7_75t_L g5357 ( 
.A(n_4664),
.Y(n_5357)
);

BUFx4f_ASAP7_75t_L g5358 ( 
.A(n_4669),
.Y(n_5358)
);

INVx2_ASAP7_75t_L g5359 ( 
.A(n_4830),
.Y(n_5359)
);

INVx2_ASAP7_75t_L g5360 ( 
.A(n_4830),
.Y(n_5360)
);

OAI21xp5_ASAP7_75t_L g5361 ( 
.A1(n_4700),
.A2(n_4878),
.B(n_4922),
.Y(n_5361)
);

AND2x4_ASAP7_75t_SL g5362 ( 
.A(n_4783),
.B(n_3279),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_4703),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_4712),
.Y(n_5364)
);

OR2x6_ASAP7_75t_L g5365 ( 
.A(n_4676),
.B(n_4777),
.Y(n_5365)
);

INVx1_ASAP7_75t_L g5366 ( 
.A(n_4712),
.Y(n_5366)
);

NAND2xp5_ASAP7_75t_SL g5367 ( 
.A(n_4827),
.B(n_1678),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_4781),
.Y(n_5368)
);

OAI22xp33_ASAP7_75t_L g5369 ( 
.A1(n_4931),
.A2(n_1202),
.B1(n_1189),
.B2(n_1192),
.Y(n_5369)
);

AND2x2_ASAP7_75t_L g5370 ( 
.A(n_4732),
.B(n_19),
.Y(n_5370)
);

O2A1O1Ixp5_ASAP7_75t_L g5371 ( 
.A1(n_4982),
.A2(n_2919),
.B(n_2921),
.C(n_2914),
.Y(n_5371)
);

O2A1O1Ixp33_ASAP7_75t_L g5372 ( 
.A1(n_4889),
.A2(n_2668),
.B(n_2676),
.C(n_2673),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_SL g5373 ( 
.A(n_4837),
.B(n_1678),
.Y(n_5373)
);

AND2x2_ASAP7_75t_L g5374 ( 
.A(n_4905),
.B(n_20),
.Y(n_5374)
);

AOI22xp33_ASAP7_75t_L g5375 ( 
.A1(n_4843),
.A2(n_1191),
.B1(n_1199),
.B2(n_1195),
.Y(n_5375)
);

INVx3_ASAP7_75t_L g5376 ( 
.A(n_4739),
.Y(n_5376)
);

BUFx6f_ASAP7_75t_L g5377 ( 
.A(n_4655),
.Y(n_5377)
);

BUFx6f_ASAP7_75t_L g5378 ( 
.A(n_4679),
.Y(n_5378)
);

AND2x2_ASAP7_75t_L g5379 ( 
.A(n_4783),
.B(n_21),
.Y(n_5379)
);

NAND2xp5_ASAP7_75t_L g5380 ( 
.A(n_4616),
.B(n_1678),
.Y(n_5380)
);

BUFx12f_ASAP7_75t_L g5381 ( 
.A(n_4710),
.Y(n_5381)
);

INVx1_ASAP7_75t_L g5382 ( 
.A(n_4782),
.Y(n_5382)
);

BUFx3_ASAP7_75t_L g5383 ( 
.A(n_4738),
.Y(n_5383)
);

OAI321xp33_ASAP7_75t_L g5384 ( 
.A1(n_4942),
.A2(n_25),
.A3(n_27),
.B1(n_28),
.B2(n_22),
.C(n_26),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_4782),
.Y(n_5385)
);

INVx2_ASAP7_75t_L g5386 ( 
.A(n_4851),
.Y(n_5386)
);

AOI22xp5_ASAP7_75t_L g5387 ( 
.A1(n_4737),
.A2(n_1200),
.B1(n_1208),
.B2(n_1678),
.Y(n_5387)
);

NAND2x1p5_ASAP7_75t_L g5388 ( 
.A(n_4664),
.B(n_3366),
.Y(n_5388)
);

BUFx3_ASAP7_75t_L g5389 ( 
.A(n_4799),
.Y(n_5389)
);

CKINVDCx5p33_ASAP7_75t_R g5390 ( 
.A(n_4725),
.Y(n_5390)
);

INVx1_ASAP7_75t_L g5391 ( 
.A(n_4785),
.Y(n_5391)
);

BUFx12f_ASAP7_75t_L g5392 ( 
.A(n_4748),
.Y(n_5392)
);

BUFx3_ASAP7_75t_L g5393 ( 
.A(n_4801),
.Y(n_5393)
);

BUFx12f_ASAP7_75t_L g5394 ( 
.A(n_4739),
.Y(n_5394)
);

INVxp67_ASAP7_75t_L g5395 ( 
.A(n_4796),
.Y(n_5395)
);

BUFx6f_ASAP7_75t_L g5396 ( 
.A(n_4774),
.Y(n_5396)
);

NAND2xp5_ASAP7_75t_SL g5397 ( 
.A(n_4725),
.B(n_1678),
.Y(n_5397)
);

BUFx3_ASAP7_75t_L g5398 ( 
.A(n_4851),
.Y(n_5398)
);

O2A1O1Ixp5_ASAP7_75t_SL g5399 ( 
.A1(n_4983),
.A2(n_3437),
.B(n_3441),
.C(n_3407),
.Y(n_5399)
);

INVx2_ASAP7_75t_L g5400 ( 
.A(n_4853),
.Y(n_5400)
);

INVx2_ASAP7_75t_L g5401 ( 
.A(n_4853),
.Y(n_5401)
);

INVx4_ASAP7_75t_L g5402 ( 
.A(n_4708),
.Y(n_5402)
);

OAI221xp5_ASAP7_75t_L g5403 ( 
.A1(n_4696),
.A2(n_947),
.B1(n_2587),
.B2(n_2576),
.C(n_2734),
.Y(n_5403)
);

CKINVDCx5p33_ASAP7_75t_R g5404 ( 
.A(n_4774),
.Y(n_5404)
);

NOR2xp33_ASAP7_75t_L g5405 ( 
.A(n_4877),
.B(n_26),
.Y(n_5405)
);

BUFx2_ASAP7_75t_L g5406 ( 
.A(n_4941),
.Y(n_5406)
);

INVx1_ASAP7_75t_L g5407 ( 
.A(n_4785),
.Y(n_5407)
);

BUFx2_ASAP7_75t_L g5408 ( 
.A(n_4784),
.Y(n_5408)
);

CKINVDCx6p67_ASAP7_75t_R g5409 ( 
.A(n_4784),
.Y(n_5409)
);

BUFx6f_ASAP7_75t_L g5410 ( 
.A(n_4810),
.Y(n_5410)
);

O2A1O1Ixp5_ASAP7_75t_L g5411 ( 
.A1(n_5085),
.A2(n_4731),
.B(n_4829),
.C(n_4753),
.Y(n_5411)
);

OAI21xp5_ASAP7_75t_L g5412 ( 
.A1(n_5207),
.A2(n_4879),
.B(n_4746),
.Y(n_5412)
);

AOI22xp33_ASAP7_75t_L g5413 ( 
.A1(n_5035),
.A2(n_4843),
.B1(n_4855),
.B2(n_5001),
.Y(n_5413)
);

INVx2_ASAP7_75t_L g5414 ( 
.A(n_5049),
.Y(n_5414)
);

BUFx3_ASAP7_75t_L g5415 ( 
.A(n_5381),
.Y(n_5415)
);

AND2x4_ASAP7_75t_L g5416 ( 
.A(n_5308),
.B(n_4983),
.Y(n_5416)
);

BUFx3_ASAP7_75t_L g5417 ( 
.A(n_5087),
.Y(n_5417)
);

CKINVDCx5p33_ASAP7_75t_R g5418 ( 
.A(n_5076),
.Y(n_5418)
);

OAI22xp5_ASAP7_75t_L g5419 ( 
.A1(n_5355),
.A2(n_4900),
.B1(n_4930),
.B2(n_4931),
.Y(n_5419)
);

BUFx2_ASAP7_75t_L g5420 ( 
.A(n_5256),
.Y(n_5420)
);

BUFx2_ASAP7_75t_L g5421 ( 
.A(n_5307),
.Y(n_5421)
);

NAND2xp5_ASAP7_75t_L g5422 ( 
.A(n_5300),
.B(n_4913),
.Y(n_5422)
);

NAND2xp5_ASAP7_75t_L g5423 ( 
.A(n_5125),
.B(n_4917),
.Y(n_5423)
);

NAND2xp5_ASAP7_75t_L g5424 ( 
.A(n_5180),
.B(n_4917),
.Y(n_5424)
);

NAND2x1p5_ASAP7_75t_L g5425 ( 
.A(n_5294),
.B(n_4900),
.Y(n_5425)
);

BUFx2_ASAP7_75t_L g5426 ( 
.A(n_5320),
.Y(n_5426)
);

INVx1_ASAP7_75t_L g5427 ( 
.A(n_5021),
.Y(n_5427)
);

NAND2xp5_ASAP7_75t_L g5428 ( 
.A(n_5106),
.B(n_4920),
.Y(n_5428)
);

INVx3_ASAP7_75t_L g5429 ( 
.A(n_5304),
.Y(n_5429)
);

NAND2xp5_ASAP7_75t_L g5430 ( 
.A(n_5106),
.B(n_4920),
.Y(n_5430)
);

INVx2_ASAP7_75t_L g5431 ( 
.A(n_5058),
.Y(n_5431)
);

AOI221xp5_ASAP7_75t_L g5432 ( 
.A1(n_5094),
.A2(n_5001),
.B1(n_5016),
.B2(n_4832),
.C(n_4800),
.Y(n_5432)
);

BUFx3_ASAP7_75t_L g5433 ( 
.A(n_5087),
.Y(n_5433)
);

INVx2_ASAP7_75t_L g5434 ( 
.A(n_5066),
.Y(n_5434)
);

HB1xp67_ASAP7_75t_L g5435 ( 
.A(n_5022),
.Y(n_5435)
);

INVx1_ASAP7_75t_SL g5436 ( 
.A(n_5128),
.Y(n_5436)
);

AOI22xp5_ASAP7_75t_L g5437 ( 
.A1(n_5182),
.A2(n_4843),
.B1(n_4934),
.B2(n_4971),
.Y(n_5437)
);

CKINVDCx6p67_ASAP7_75t_R g5438 ( 
.A(n_5232),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5046),
.Y(n_5439)
);

BUFx3_ASAP7_75t_L g5440 ( 
.A(n_5091),
.Y(n_5440)
);

INVx3_ASAP7_75t_L g5441 ( 
.A(n_5304),
.Y(n_5441)
);

BUFx6f_ASAP7_75t_L g5442 ( 
.A(n_5169),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_5078),
.Y(n_5443)
);

INVx1_ASAP7_75t_L g5444 ( 
.A(n_5079),
.Y(n_5444)
);

INVx2_ASAP7_75t_L g5445 ( 
.A(n_5086),
.Y(n_5445)
);

AOI22xp33_ASAP7_75t_L g5446 ( 
.A1(n_5060),
.A2(n_4843),
.B1(n_5016),
.B2(n_4824),
.Y(n_5446)
);

BUFx6f_ASAP7_75t_L g5447 ( 
.A(n_5396),
.Y(n_5447)
);

INVxp67_ASAP7_75t_SL g5448 ( 
.A(n_5334),
.Y(n_5448)
);

BUFx6f_ASAP7_75t_L g5449 ( 
.A(n_5396),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_5082),
.Y(n_5450)
);

INVx1_ASAP7_75t_L g5451 ( 
.A(n_5096),
.Y(n_5451)
);

BUFx6f_ASAP7_75t_L g5452 ( 
.A(n_5396),
.Y(n_5452)
);

AND2x2_ASAP7_75t_L g5453 ( 
.A(n_5101),
.B(n_4979),
.Y(n_5453)
);

OR2x6_ASAP7_75t_L g5454 ( 
.A(n_5365),
.B(n_4777),
.Y(n_5454)
);

AND2x6_ASAP7_75t_L g5455 ( 
.A(n_5332),
.B(n_4993),
.Y(n_5455)
);

AO21x1_ASAP7_75t_L g5456 ( 
.A1(n_5052),
.A2(n_5166),
.B(n_5313),
.Y(n_5456)
);

A2O1A1Ixp33_ASAP7_75t_L g5457 ( 
.A1(n_5212),
.A2(n_4900),
.B(n_4934),
.C(n_4992),
.Y(n_5457)
);

BUFx6f_ASAP7_75t_L g5458 ( 
.A(n_5410),
.Y(n_5458)
);

AND2x4_ASAP7_75t_L g5459 ( 
.A(n_5023),
.B(n_4978),
.Y(n_5459)
);

BUFx6f_ASAP7_75t_L g5460 ( 
.A(n_5410),
.Y(n_5460)
);

HB1xp67_ASAP7_75t_L g5461 ( 
.A(n_5337),
.Y(n_5461)
);

INVx3_ASAP7_75t_L g5462 ( 
.A(n_5042),
.Y(n_5462)
);

AND2x4_ASAP7_75t_L g5463 ( 
.A(n_5119),
.B(n_4993),
.Y(n_5463)
);

BUFx2_ASAP7_75t_L g5464 ( 
.A(n_5344),
.Y(n_5464)
);

AOI21xp5_ASAP7_75t_L g5465 ( 
.A1(n_5040),
.A2(n_4992),
.B(n_4675),
.Y(n_5465)
);

AOI21xp5_ASAP7_75t_L g5466 ( 
.A1(n_5040),
.A2(n_4981),
.B(n_4954),
.Y(n_5466)
);

AOI22xp33_ASAP7_75t_L g5467 ( 
.A1(n_5121),
.A2(n_4824),
.B1(n_4658),
.B2(n_4791),
.Y(n_5467)
);

INVx3_ASAP7_75t_L g5468 ( 
.A(n_5042),
.Y(n_5468)
);

AOI21xp5_ASAP7_75t_L g5469 ( 
.A1(n_5249),
.A2(n_4873),
.B(n_4794),
.Y(n_5469)
);

INVx3_ASAP7_75t_L g5470 ( 
.A(n_5055),
.Y(n_5470)
);

OAI21x1_ASAP7_75t_L g5471 ( 
.A1(n_5018),
.A2(n_5011),
.B(n_5010),
.Y(n_5471)
);

AND2x4_ASAP7_75t_L g5472 ( 
.A(n_5229),
.B(n_5015),
.Y(n_5472)
);

HB1xp67_ASAP7_75t_L g5473 ( 
.A(n_5337),
.Y(n_5473)
);

AOI21xp5_ASAP7_75t_L g5474 ( 
.A1(n_5249),
.A2(n_5070),
.B(n_5328),
.Y(n_5474)
);

AOI22xp33_ASAP7_75t_L g5475 ( 
.A1(n_5375),
.A2(n_4824),
.B1(n_4658),
.B2(n_4791),
.Y(n_5475)
);

AOI21xp5_ASAP7_75t_L g5476 ( 
.A1(n_5328),
.A2(n_4873),
.B(n_4794),
.Y(n_5476)
);

O2A1O1Ixp5_ASAP7_75t_SL g5477 ( 
.A1(n_5206),
.A2(n_5015),
.B(n_4991),
.C(n_4999),
.Y(n_5477)
);

OAI221xp5_ASAP7_75t_L g5478 ( 
.A1(n_5105),
.A2(n_4702),
.B1(n_4685),
.B2(n_4632),
.C(n_4689),
.Y(n_5478)
);

AOI21xp5_ASAP7_75t_L g5479 ( 
.A1(n_5028),
.A2(n_4787),
.B(n_4956),
.Y(n_5479)
);

A2O1A1Ixp33_ASAP7_75t_L g5480 ( 
.A1(n_5212),
.A2(n_4891),
.B(n_4685),
.C(n_4632),
.Y(n_5480)
);

AOI22xp5_ASAP7_75t_L g5481 ( 
.A1(n_5118),
.A2(n_4824),
.B1(n_4658),
.B2(n_4791),
.Y(n_5481)
);

O2A1O1Ixp33_ASAP7_75t_L g5482 ( 
.A1(n_5094),
.A2(n_5238),
.B(n_5230),
.C(n_5075),
.Y(n_5482)
);

NAND2xp5_ASAP7_75t_L g5483 ( 
.A(n_5044),
.B(n_4925),
.Y(n_5483)
);

OR2x6_ASAP7_75t_L g5484 ( 
.A(n_5365),
.B(n_4777),
.Y(n_5484)
);

BUFx6f_ASAP7_75t_L g5485 ( 
.A(n_5410),
.Y(n_5485)
);

INVx3_ASAP7_75t_L g5486 ( 
.A(n_5055),
.Y(n_5486)
);

AOI21xp5_ASAP7_75t_L g5487 ( 
.A1(n_5028),
.A2(n_4787),
.B(n_4686),
.Y(n_5487)
);

INVx3_ASAP7_75t_L g5488 ( 
.A(n_5059),
.Y(n_5488)
);

INVx4_ASAP7_75t_L g5489 ( 
.A(n_5232),
.Y(n_5489)
);

BUFx3_ASAP7_75t_L g5490 ( 
.A(n_5131),
.Y(n_5490)
);

AND2x2_ASAP7_75t_L g5491 ( 
.A(n_5144),
.B(n_4988),
.Y(n_5491)
);

AOI21xp5_ASAP7_75t_L g5492 ( 
.A1(n_5032),
.A2(n_4787),
.B(n_4686),
.Y(n_5492)
);

AOI22xp33_ASAP7_75t_L g5493 ( 
.A1(n_5314),
.A2(n_4824),
.B1(n_4658),
.B2(n_4791),
.Y(n_5493)
);

BUFx2_ASAP7_75t_L g5494 ( 
.A(n_5054),
.Y(n_5494)
);

AND2x4_ASAP7_75t_L g5495 ( 
.A(n_5365),
.B(n_5002),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5097),
.Y(n_5496)
);

BUFx6f_ASAP7_75t_L g5497 ( 
.A(n_5394),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5100),
.Y(n_5498)
);

BUFx3_ASAP7_75t_L g5499 ( 
.A(n_5224),
.Y(n_5499)
);

INVxp67_ASAP7_75t_SL g5500 ( 
.A(n_5043),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_5057),
.B(n_4925),
.Y(n_5501)
);

OR2x6_ASAP7_75t_L g5502 ( 
.A(n_5270),
.B(n_4726),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_5130),
.Y(n_5503)
);

AOI21xp5_ASAP7_75t_L g5504 ( 
.A1(n_5092),
.A2(n_4736),
.B(n_4882),
.Y(n_5504)
);

AND2x4_ASAP7_75t_L g5505 ( 
.A(n_5164),
.B(n_5002),
.Y(n_5505)
);

OAI22xp5_ASAP7_75t_L g5506 ( 
.A1(n_5232),
.A2(n_4929),
.B1(n_4949),
.B2(n_4689),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_5160),
.Y(n_5507)
);

AND2x2_ASAP7_75t_L g5508 ( 
.A(n_5071),
.B(n_5008),
.Y(n_5508)
);

BUFx2_ASAP7_75t_R g5509 ( 
.A(n_5102),
.Y(n_5509)
);

BUFx6f_ASAP7_75t_L g5510 ( 
.A(n_5378),
.Y(n_5510)
);

OR2x6_ASAP7_75t_L g5511 ( 
.A(n_5270),
.B(n_5195),
.Y(n_5511)
);

AND2x2_ASAP7_75t_L g5512 ( 
.A(n_5161),
.B(n_4939),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_5188),
.Y(n_5513)
);

INVx2_ASAP7_75t_L g5514 ( 
.A(n_5098),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_5099),
.Y(n_5515)
);

BUFx2_ASAP7_75t_L g5516 ( 
.A(n_5209),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_5111),
.Y(n_5517)
);

INVx2_ASAP7_75t_L g5518 ( 
.A(n_5117),
.Y(n_5518)
);

AOI21xp5_ASAP7_75t_L g5519 ( 
.A1(n_5361),
.A2(n_4882),
.B(n_4969),
.Y(n_5519)
);

NAND2xp5_ASAP7_75t_L g5520 ( 
.A(n_5187),
.B(n_4940),
.Y(n_5520)
);

HB1xp67_ASAP7_75t_L g5521 ( 
.A(n_5255),
.Y(n_5521)
);

AOI22xp33_ASAP7_75t_L g5522 ( 
.A1(n_5034),
.A2(n_4658),
.B1(n_4791),
.B2(n_4973),
.Y(n_5522)
);

NAND3xp33_ASAP7_75t_L g5523 ( 
.A(n_5147),
.B(n_5000),
.C(n_4995),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_5126),
.Y(n_5524)
);

INVx2_ASAP7_75t_SL g5525 ( 
.A(n_5383),
.Y(n_5525)
);

NAND2xp5_ASAP7_75t_L g5526 ( 
.A(n_5158),
.B(n_4944),
.Y(n_5526)
);

INVx2_ASAP7_75t_L g5527 ( 
.A(n_5139),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5143),
.Y(n_5528)
);

AND2x4_ASAP7_75t_L g5529 ( 
.A(n_5184),
.B(n_5006),
.Y(n_5529)
);

INVx1_ASAP7_75t_L g5530 ( 
.A(n_5148),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_5153),
.Y(n_5531)
);

BUFx3_ASAP7_75t_L g5532 ( 
.A(n_5224),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_5157),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_5162),
.Y(n_5534)
);

HB1xp67_ASAP7_75t_L g5535 ( 
.A(n_5255),
.Y(n_5535)
);

INVx4_ASAP7_75t_L g5536 ( 
.A(n_5136),
.Y(n_5536)
);

BUFx6f_ASAP7_75t_L g5537 ( 
.A(n_5378),
.Y(n_5537)
);

BUFx5_ASAP7_75t_L g5538 ( 
.A(n_5110),
.Y(n_5538)
);

AND2x4_ASAP7_75t_L g5539 ( 
.A(n_5333),
.B(n_5014),
.Y(n_5539)
);

AND2x6_ASAP7_75t_L g5540 ( 
.A(n_5332),
.B(n_4871),
.Y(n_5540)
);

AND2x2_ASAP7_75t_L g5541 ( 
.A(n_5050),
.B(n_4946),
.Y(n_5541)
);

NAND2xp5_ASAP7_75t_L g5542 ( 
.A(n_5306),
.B(n_4862),
.Y(n_5542)
);

INVx1_ASAP7_75t_L g5543 ( 
.A(n_5302),
.Y(n_5543)
);

BUFx3_ASAP7_75t_L g5544 ( 
.A(n_5246),
.Y(n_5544)
);

AOI21xp5_ASAP7_75t_L g5545 ( 
.A1(n_5361),
.A2(n_4975),
.B(n_4969),
.Y(n_5545)
);

AND2x2_ASAP7_75t_L g5546 ( 
.A(n_5343),
.B(n_4751),
.Y(n_5546)
);

NAND2xp5_ASAP7_75t_L g5547 ( 
.A(n_5172),
.B(n_4869),
.Y(n_5547)
);

INVx1_ASAP7_75t_L g5548 ( 
.A(n_5027),
.Y(n_5548)
);

INVx3_ASAP7_75t_L g5549 ( 
.A(n_5059),
.Y(n_5549)
);

NOR2xp67_ASAP7_75t_L g5550 ( 
.A(n_5281),
.B(n_4918),
.Y(n_5550)
);

BUFx2_ASAP7_75t_L g5551 ( 
.A(n_5228),
.Y(n_5551)
);

AND2x4_ASAP7_75t_L g5552 ( 
.A(n_5140),
.B(n_5014),
.Y(n_5552)
);

AOI21xp5_ASAP7_75t_L g5553 ( 
.A1(n_5318),
.A2(n_4975),
.B(n_4953),
.Y(n_5553)
);

INVx5_ASAP7_75t_L g5554 ( 
.A(n_5252),
.Y(n_5554)
);

BUFx2_ASAP7_75t_L g5555 ( 
.A(n_5228),
.Y(n_5555)
);

BUFx3_ASAP7_75t_L g5556 ( 
.A(n_5133),
.Y(n_5556)
);

AOI21xp5_ASAP7_75t_L g5557 ( 
.A1(n_5325),
.A2(n_4953),
.B(n_4966),
.Y(n_5557)
);

BUFx3_ASAP7_75t_L g5558 ( 
.A(n_5045),
.Y(n_5558)
);

BUFx6f_ASAP7_75t_L g5559 ( 
.A(n_5378),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_5213),
.Y(n_5560)
);

INVx1_ASAP7_75t_SL g5561 ( 
.A(n_5321),
.Y(n_5561)
);

INVx2_ASAP7_75t_L g5562 ( 
.A(n_5312),
.Y(n_5562)
);

INVx2_ASAP7_75t_SL g5563 ( 
.A(n_5358),
.Y(n_5563)
);

INVx2_ASAP7_75t_SL g5564 ( 
.A(n_5358),
.Y(n_5564)
);

INVx2_ASAP7_75t_SL g5565 ( 
.A(n_5198),
.Y(n_5565)
);

NAND2xp5_ASAP7_75t_L g5566 ( 
.A(n_5031),
.B(n_4857),
.Y(n_5566)
);

INVx2_ASAP7_75t_SL g5567 ( 
.A(n_5237),
.Y(n_5567)
);

AND2x2_ASAP7_75t_L g5568 ( 
.A(n_5112),
.B(n_4751),
.Y(n_5568)
);

NAND2xp5_ASAP7_75t_L g5569 ( 
.A(n_5293),
.B(n_4864),
.Y(n_5569)
);

INVx2_ASAP7_75t_L g5570 ( 
.A(n_5242),
.Y(n_5570)
);

BUFx6f_ASAP7_75t_L g5571 ( 
.A(n_5316),
.Y(n_5571)
);

NAND2xp5_ASAP7_75t_L g5572 ( 
.A(n_5351),
.B(n_5363),
.Y(n_5572)
);

INVx1_ASAP7_75t_L g5573 ( 
.A(n_5245),
.Y(n_5573)
);

NAND2xp5_ASAP7_75t_L g5574 ( 
.A(n_5364),
.B(n_4880),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_5248),
.Y(n_5575)
);

O2A1O1Ixp5_ASAP7_75t_L g5576 ( 
.A1(n_5103),
.A2(n_4834),
.B(n_4867),
.C(n_4810),
.Y(n_5576)
);

AND2x4_ASAP7_75t_L g5577 ( 
.A(n_5140),
.B(n_5051),
.Y(n_5577)
);

INVx1_ASAP7_75t_SL g5578 ( 
.A(n_5340),
.Y(n_5578)
);

CKINVDCx5p33_ASAP7_75t_R g5579 ( 
.A(n_5047),
.Y(n_5579)
);

AND2x4_ASAP7_75t_L g5580 ( 
.A(n_5140),
.B(n_4973),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_5257),
.Y(n_5581)
);

INVx1_ASAP7_75t_L g5582 ( 
.A(n_5322),
.Y(n_5582)
);

INVx2_ASAP7_75t_SL g5583 ( 
.A(n_5288),
.Y(n_5583)
);

INVx1_ASAP7_75t_SL g5584 ( 
.A(n_5056),
.Y(n_5584)
);

INVxp67_ASAP7_75t_L g5585 ( 
.A(n_5104),
.Y(n_5585)
);

BUFx2_ASAP7_75t_L g5586 ( 
.A(n_5254),
.Y(n_5586)
);

NAND2xp5_ASAP7_75t_L g5587 ( 
.A(n_5366),
.B(n_5088),
.Y(n_5587)
);

INVx3_ASAP7_75t_L g5588 ( 
.A(n_5168),
.Y(n_5588)
);

INVx3_ASAP7_75t_R g5589 ( 
.A(n_5408),
.Y(n_5589)
);

INVx2_ASAP7_75t_SL g5590 ( 
.A(n_5056),
.Y(n_5590)
);

BUFx4f_ASAP7_75t_SL g5591 ( 
.A(n_5219),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5331),
.Y(n_5592)
);

O2A1O1Ixp33_ASAP7_75t_L g5593 ( 
.A1(n_5129),
.A2(n_4695),
.B(n_4747),
.C(n_4750),
.Y(n_5593)
);

AOI222xp33_ASAP7_75t_L g5594 ( 
.A1(n_5354),
.A2(n_4973),
.B1(n_4747),
.B2(n_4727),
.C1(n_4897),
.C2(n_4895),
.Y(n_5594)
);

NOR2xp33_ASAP7_75t_L g5595 ( 
.A(n_5392),
.B(n_4834),
.Y(n_5595)
);

NOR3xp33_ASAP7_75t_L g5596 ( 
.A(n_5167),
.B(n_4867),
.C(n_4750),
.Y(n_5596)
);

OAI21x1_ASAP7_75t_L g5597 ( 
.A1(n_5038),
.A2(n_5020),
.B(n_5077),
.Y(n_5597)
);

BUFx6f_ASAP7_75t_L g5598 ( 
.A(n_5019),
.Y(n_5598)
);

AOI22xp33_ASAP7_75t_L g5599 ( 
.A1(n_5226),
.A2(n_4973),
.B1(n_4916),
.B2(n_4871),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_5260),
.Y(n_5600)
);

O2A1O1Ixp33_ASAP7_75t_SL g5601 ( 
.A1(n_5189),
.A2(n_4727),
.B(n_4715),
.C(n_4740),
.Y(n_5601)
);

BUFx2_ASAP7_75t_L g5602 ( 
.A(n_5254),
.Y(n_5602)
);

INVxp67_ASAP7_75t_L g5603 ( 
.A(n_5149),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_5239),
.Y(n_5604)
);

INVx2_ASAP7_75t_L g5605 ( 
.A(n_5269),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5336),
.Y(n_5606)
);

AND2x4_ASAP7_75t_L g5607 ( 
.A(n_5051),
.B(n_4973),
.Y(n_5607)
);

AOI22xp33_ASAP7_75t_L g5608 ( 
.A1(n_5142),
.A2(n_5062),
.B1(n_5405),
.B2(n_5095),
.Y(n_5608)
);

NAND2xp5_ASAP7_75t_L g5609 ( 
.A(n_5068),
.B(n_5368),
.Y(n_5609)
);

HB1xp67_ASAP7_75t_L g5610 ( 
.A(n_5067),
.Y(n_5610)
);

AOI22xp33_ASAP7_75t_L g5611 ( 
.A1(n_5039),
.A2(n_4916),
.B1(n_4802),
.B2(n_4769),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_5349),
.Y(n_5612)
);

OR2x6_ASAP7_75t_L g5613 ( 
.A(n_5406),
.B(n_4726),
.Y(n_5613)
);

OAI21xp33_ASAP7_75t_L g5614 ( 
.A1(n_5072),
.A2(n_5004),
.B(n_5003),
.Y(n_5614)
);

OR2x2_ASAP7_75t_L g5615 ( 
.A(n_5030),
.B(n_4619),
.Y(n_5615)
);

AND2x2_ASAP7_75t_L g5616 ( 
.A(n_5395),
.B(n_4769),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5171),
.Y(n_5617)
);

AND2x2_ASAP7_75t_L g5618 ( 
.A(n_5236),
.B(n_4802),
.Y(n_5618)
);

INVx3_ASAP7_75t_L g5619 ( 
.A(n_5168),
.Y(n_5619)
);

AND2x4_ASAP7_75t_L g5620 ( 
.A(n_5109),
.B(n_4619),
.Y(n_5620)
);

NAND2xp5_ASAP7_75t_L g5621 ( 
.A(n_5382),
.B(n_4849),
.Y(n_5621)
);

NAND2xp5_ASAP7_75t_L g5622 ( 
.A(n_5385),
.B(n_4936),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_5218),
.Y(n_5623)
);

BUFx6f_ASAP7_75t_L g5624 ( 
.A(n_5019),
.Y(n_5624)
);

INVx2_ASAP7_75t_SL g5625 ( 
.A(n_5389),
.Y(n_5625)
);

INVx3_ASAP7_75t_L g5626 ( 
.A(n_5262),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5218),
.Y(n_5627)
);

AND2x2_ASAP7_75t_L g5628 ( 
.A(n_5347),
.B(n_4657),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_5305),
.Y(n_5629)
);

OAI22xp5_ASAP7_75t_L g5630 ( 
.A1(n_5116),
.A2(n_5197),
.B1(n_5267),
.B2(n_5189),
.Y(n_5630)
);

CKINVDCx20_ASAP7_75t_R g5631 ( 
.A(n_5083),
.Y(n_5631)
);

INVx1_ASAP7_75t_L g5632 ( 
.A(n_5218),
.Y(n_5632)
);

AND2x4_ASAP7_75t_L g5633 ( 
.A(n_5109),
.B(n_4657),
.Y(n_5633)
);

CKINVDCx6p67_ASAP7_75t_R g5634 ( 
.A(n_5037),
.Y(n_5634)
);

INVx2_ASAP7_75t_L g5635 ( 
.A(n_5173),
.Y(n_5635)
);

CKINVDCx5p33_ASAP7_75t_R g5636 ( 
.A(n_5029),
.Y(n_5636)
);

INVx1_ASAP7_75t_SL g5637 ( 
.A(n_5404),
.Y(n_5637)
);

AND2x4_ASAP7_75t_L g5638 ( 
.A(n_5217),
.B(n_4693),
.Y(n_5638)
);

AND2x2_ASAP7_75t_L g5639 ( 
.A(n_5359),
.B(n_4693),
.Y(n_5639)
);

O2A1O1Ixp5_ASAP7_75t_L g5640 ( 
.A1(n_5115),
.A2(n_4745),
.B(n_5009),
.C(n_5004),
.Y(n_5640)
);

OR2x2_ASAP7_75t_L g5641 ( 
.A(n_5231),
.B(n_5003),
.Y(n_5641)
);

NAND2xp5_ASAP7_75t_L g5642 ( 
.A(n_5391),
.B(n_5009),
.Y(n_5642)
);

BUFx4f_ASAP7_75t_SL g5643 ( 
.A(n_5073),
.Y(n_5643)
);

INVx1_ASAP7_75t_L g5644 ( 
.A(n_5176),
.Y(n_5644)
);

INVx2_ASAP7_75t_L g5645 ( 
.A(n_5193),
.Y(n_5645)
);

INVx1_ASAP7_75t_L g5646 ( 
.A(n_5199),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_5200),
.Y(n_5647)
);

AND2x4_ASAP7_75t_L g5648 ( 
.A(n_5217),
.B(n_4745),
.Y(n_5648)
);

INVx3_ASAP7_75t_L g5649 ( 
.A(n_5262),
.Y(n_5649)
);

NOR2xp33_ASAP7_75t_L g5650 ( 
.A(n_5155),
.B(n_4943),
.Y(n_5650)
);

INVx1_ASAP7_75t_L g5651 ( 
.A(n_5216),
.Y(n_5651)
);

INVx1_ASAP7_75t_L g5652 ( 
.A(n_5251),
.Y(n_5652)
);

AND2x4_ASAP7_75t_L g5653 ( 
.A(n_5217),
.B(n_4987),
.Y(n_5653)
);

NAND3xp33_ASAP7_75t_L g5654 ( 
.A(n_5147),
.B(n_4987),
.C(n_4838),
.Y(n_5654)
);

NAND2xp5_ASAP7_75t_L g5655 ( 
.A(n_5407),
.B(n_4715),
.Y(n_5655)
);

AND2x4_ASAP7_75t_L g5656 ( 
.A(n_5145),
.B(n_4996),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_5261),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_5360),
.B(n_4943),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_5264),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_5274),
.Y(n_5660)
);

INVx2_ASAP7_75t_L g5661 ( 
.A(n_5275),
.Y(n_5661)
);

AND2x2_ASAP7_75t_L g5662 ( 
.A(n_5279),
.B(n_4966),
.Y(n_5662)
);

INVx2_ASAP7_75t_L g5663 ( 
.A(n_5284),
.Y(n_5663)
);

INVx2_ASAP7_75t_L g5664 ( 
.A(n_5292),
.Y(n_5664)
);

INVx1_ASAP7_75t_SL g5665 ( 
.A(n_5393),
.Y(n_5665)
);

INVx2_ASAP7_75t_L g5666 ( 
.A(n_5298),
.Y(n_5666)
);

CKINVDCx16_ASAP7_75t_R g5667 ( 
.A(n_5048),
.Y(n_5667)
);

NAND2xp5_ASAP7_75t_L g5668 ( 
.A(n_5033),
.B(n_4838),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_5113),
.Y(n_5669)
);

INVx2_ASAP7_75t_SL g5670 ( 
.A(n_5064),
.Y(n_5670)
);

BUFx6f_ASAP7_75t_L g5671 ( 
.A(n_5019),
.Y(n_5671)
);

INVx2_ASAP7_75t_SL g5672 ( 
.A(n_5064),
.Y(n_5672)
);

CKINVDCx5p33_ASAP7_75t_R g5673 ( 
.A(n_5204),
.Y(n_5673)
);

AOI21xp33_ASAP7_75t_SL g5674 ( 
.A1(n_5026),
.A2(n_28),
.B(n_29),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5063),
.Y(n_5675)
);

NAND2xp5_ASAP7_75t_L g5676 ( 
.A(n_5053),
.B(n_4740),
.Y(n_5676)
);

INVx2_ASAP7_75t_L g5677 ( 
.A(n_5386),
.Y(n_5677)
);

NAND2x1_ASAP7_75t_L g5678 ( 
.A(n_5145),
.B(n_4996),
.Y(n_5678)
);

OAI21x1_ASAP7_75t_SL g5679 ( 
.A1(n_5151),
.A2(n_4761),
.B(n_4894),
.Y(n_5679)
);

NOR2xp33_ASAP7_75t_L g5680 ( 
.A(n_5348),
.B(n_29),
.Y(n_5680)
);

INVx1_ASAP7_75t_SL g5681 ( 
.A(n_5398),
.Y(n_5681)
);

INVx2_ASAP7_75t_L g5682 ( 
.A(n_5400),
.Y(n_5682)
);

BUFx4_ASAP7_75t_SL g5683 ( 
.A(n_5390),
.Y(n_5683)
);

AOI21xp5_ASAP7_75t_L g5684 ( 
.A1(n_5156),
.A2(n_5194),
.B(n_5141),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_5053),
.Y(n_5685)
);

INVx2_ASAP7_75t_L g5686 ( 
.A(n_5401),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5063),
.Y(n_5687)
);

AND2x4_ASAP7_75t_L g5688 ( 
.A(n_5178),
.B(n_4998),
.Y(n_5688)
);

INVx2_ASAP7_75t_L g5689 ( 
.A(n_5279),
.Y(n_5689)
);

CKINVDCx20_ASAP7_75t_R g5690 ( 
.A(n_5287),
.Y(n_5690)
);

AOI21x1_ASAP7_75t_L g5691 ( 
.A1(n_5159),
.A2(n_4884),
.B(n_4876),
.Y(n_5691)
);

AOI21xp33_ASAP7_75t_L g5692 ( 
.A1(n_5369),
.A2(n_4884),
.B(n_4876),
.Y(n_5692)
);

AND2x2_ASAP7_75t_L g5693 ( 
.A(n_5286),
.B(n_5297),
.Y(n_5693)
);

CKINVDCx5p33_ASAP7_75t_R g5694 ( 
.A(n_5037),
.Y(n_5694)
);

AO22x1_ASAP7_75t_L g5695 ( 
.A1(n_5108),
.A2(n_4894),
.B1(n_4847),
.B2(n_4741),
.Y(n_5695)
);

CKINVDCx6p67_ASAP7_75t_R g5696 ( 
.A(n_5185),
.Y(n_5696)
);

BUFx2_ASAP7_75t_L g5697 ( 
.A(n_5178),
.Y(n_5697)
);

O2A1O1Ixp33_ASAP7_75t_L g5698 ( 
.A1(n_5114),
.A2(n_5356),
.B(n_5291),
.C(n_5295),
.Y(n_5698)
);

NAND2xp5_ASAP7_75t_L g5699 ( 
.A(n_5137),
.B(n_4755),
.Y(n_5699)
);

AND2x2_ASAP7_75t_L g5700 ( 
.A(n_5286),
.B(n_5297),
.Y(n_5700)
);

AND2x2_ASAP7_75t_L g5701 ( 
.A(n_5127),
.B(n_4755),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_5165),
.Y(n_5702)
);

BUFx2_ASAP7_75t_L g5703 ( 
.A(n_5093),
.Y(n_5703)
);

BUFx6f_ASAP7_75t_L g5704 ( 
.A(n_5061),
.Y(n_5704)
);

INVx1_ASAP7_75t_L g5705 ( 
.A(n_5159),
.Y(n_5705)
);

INVx1_ASAP7_75t_SL g5706 ( 
.A(n_5409),
.Y(n_5706)
);

NAND2x1p5_ASAP7_75t_L g5707 ( 
.A(n_5272),
.B(n_4766),
.Y(n_5707)
);

INVx2_ASAP7_75t_L g5708 ( 
.A(n_5135),
.Y(n_5708)
);

INVx2_ASAP7_75t_SL g5709 ( 
.A(n_5138),
.Y(n_5709)
);

A2O1A1Ixp33_ASAP7_75t_L g5710 ( 
.A1(n_5384),
.A2(n_4847),
.B(n_4741),
.C(n_4772),
.Y(n_5710)
);

NAND2xp5_ASAP7_75t_L g5711 ( 
.A(n_5137),
.B(n_4766),
.Y(n_5711)
);

INVx5_ASAP7_75t_L g5712 ( 
.A(n_5252),
.Y(n_5712)
);

OR2x6_ASAP7_75t_L g5713 ( 
.A(n_5289),
.B(n_4772),
.Y(n_5713)
);

AOI22xp33_ASAP7_75t_L g5714 ( 
.A1(n_5354),
.A2(n_4778),
.B1(n_4776),
.B2(n_4850),
.Y(n_5714)
);

NAND2xp5_ASAP7_75t_L g5715 ( 
.A(n_5380),
.B(n_5283),
.Y(n_5715)
);

OAI22xp5_ASAP7_75t_L g5716 ( 
.A1(n_5116),
.A2(n_4778),
.B1(n_4776),
.B2(n_4850),
.Y(n_5716)
);

BUFx6f_ASAP7_75t_L g5717 ( 
.A(n_5061),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_5299),
.Y(n_5718)
);

BUFx2_ASAP7_75t_L g5719 ( 
.A(n_5093),
.Y(n_5719)
);

NAND2xp5_ASAP7_75t_L g5720 ( 
.A(n_5380),
.B(n_4852),
.Y(n_5720)
);

AND2x4_ASAP7_75t_L g5721 ( 
.A(n_5289),
.B(n_4852),
.Y(n_5721)
);

AOI22xp33_ASAP7_75t_L g5722 ( 
.A1(n_5181),
.A2(n_2587),
.B1(n_2576),
.B2(n_2734),
.Y(n_5722)
);

AND2x4_ASAP7_75t_L g5723 ( 
.A(n_5289),
.B(n_30),
.Y(n_5723)
);

NAND2xp5_ASAP7_75t_L g5724 ( 
.A(n_5283),
.B(n_31),
.Y(n_5724)
);

AND2x4_ASAP7_75t_L g5725 ( 
.A(n_5324),
.B(n_32),
.Y(n_5725)
);

INVx2_ASAP7_75t_L g5726 ( 
.A(n_5135),
.Y(n_5726)
);

INVx1_ASAP7_75t_L g5727 ( 
.A(n_5036),
.Y(n_5727)
);

NAND2x1p5_ASAP7_75t_L g5728 ( 
.A(n_5272),
.B(n_3367),
.Y(n_5728)
);

AND2x2_ASAP7_75t_L g5729 ( 
.A(n_5296),
.B(n_32),
.Y(n_5729)
);

BUFx6f_ASAP7_75t_L g5730 ( 
.A(n_5061),
.Y(n_5730)
);

BUFx12f_ASAP7_75t_L g5731 ( 
.A(n_5345),
.Y(n_5731)
);

INVx2_ASAP7_75t_SL g5732 ( 
.A(n_5138),
.Y(n_5732)
);

NAND2xp5_ASAP7_75t_L g5733 ( 
.A(n_5191),
.B(n_33),
.Y(n_5733)
);

AND2x4_ASAP7_75t_L g5734 ( 
.A(n_5324),
.B(n_33),
.Y(n_5734)
);

BUFx6f_ASAP7_75t_L g5735 ( 
.A(n_5069),
.Y(n_5735)
);

NAND2xp5_ASAP7_75t_L g5736 ( 
.A(n_5353),
.B(n_35),
.Y(n_5736)
);

INVxp67_ASAP7_75t_L g5737 ( 
.A(n_5163),
.Y(n_5737)
);

AOI22xp5_ASAP7_75t_L g5738 ( 
.A1(n_5065),
.A2(n_2587),
.B1(n_2734),
.B2(n_2947),
.Y(n_5738)
);

OAI21xp33_ASAP7_75t_SL g5739 ( 
.A1(n_5285),
.A2(n_5402),
.B(n_5357),
.Y(n_5739)
);

BUFx2_ASAP7_75t_L g5740 ( 
.A(n_5107),
.Y(n_5740)
);

BUFx4_ASAP7_75t_SL g5741 ( 
.A(n_5185),
.Y(n_5741)
);

NAND2xp5_ASAP7_75t_L g5742 ( 
.A(n_5335),
.B(n_36),
.Y(n_5742)
);

O2A1O1Ixp5_ASAP7_75t_SL g5743 ( 
.A1(n_5376),
.A2(n_3437),
.B(n_3441),
.C(n_3407),
.Y(n_5743)
);

INVx2_ASAP7_75t_L g5744 ( 
.A(n_5202),
.Y(n_5744)
);

AOI22xp33_ASAP7_75t_L g5745 ( 
.A1(n_5017),
.A2(n_5374),
.B1(n_5174),
.B2(n_5309),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5036),
.Y(n_5746)
);

AOI21xp5_ASAP7_75t_L g5747 ( 
.A1(n_5150),
.A2(n_3374),
.B(n_3367),
.Y(n_5747)
);

OAI21x1_ASAP7_75t_L g5748 ( 
.A1(n_5477),
.A2(n_5240),
.B(n_5350),
.Y(n_5748)
);

AND2x4_ASAP7_75t_L g5749 ( 
.A(n_5620),
.B(n_5036),
.Y(n_5749)
);

OAI21x1_ASAP7_75t_SL g5750 ( 
.A1(n_5456),
.A2(n_5259),
.B(n_5290),
.Y(n_5750)
);

INVx1_ASAP7_75t_L g5751 ( 
.A(n_5513),
.Y(n_5751)
);

AOI22xp33_ASAP7_75t_L g5752 ( 
.A1(n_5630),
.A2(n_5024),
.B1(n_5397),
.B2(n_5247),
.Y(n_5752)
);

AOI22xp5_ASAP7_75t_L g5753 ( 
.A1(n_5608),
.A2(n_5122),
.B1(n_5146),
.B2(n_5267),
.Y(n_5753)
);

OAI21xp5_ASAP7_75t_L g5754 ( 
.A1(n_5457),
.A2(n_5167),
.B(n_5384),
.Y(n_5754)
);

NAND2x1p5_ASAP7_75t_L g5755 ( 
.A(n_5554),
.B(n_5120),
.Y(n_5755)
);

INVx2_ASAP7_75t_SL g5756 ( 
.A(n_5442),
.Y(n_5756)
);

INVx2_ASAP7_75t_L g5757 ( 
.A(n_5464),
.Y(n_5757)
);

NAND2x1p5_ASAP7_75t_L g5758 ( 
.A(n_5554),
.B(n_5120),
.Y(n_5758)
);

INVx1_ASAP7_75t_L g5759 ( 
.A(n_5513),
.Y(n_5759)
);

O2A1O1Ixp33_ASAP7_75t_SL g5760 ( 
.A1(n_5674),
.A2(n_5175),
.B(n_5210),
.C(n_5339),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_5515),
.Y(n_5761)
);

BUFx2_ASAP7_75t_L g5762 ( 
.A(n_5511),
.Y(n_5762)
);

OAI21x1_ASAP7_75t_L g5763 ( 
.A1(n_5597),
.A2(n_5399),
.B(n_5259),
.Y(n_5763)
);

AO21x2_ASAP7_75t_L g5764 ( 
.A1(n_5708),
.A2(n_5081),
.B(n_5299),
.Y(n_5764)
);

INVx3_ASAP7_75t_L g5765 ( 
.A(n_5429),
.Y(n_5765)
);

OAI21x1_ASAP7_75t_L g5766 ( 
.A1(n_5471),
.A2(n_5081),
.B(n_5371),
.Y(n_5766)
);

OAI21x1_ASAP7_75t_L g5767 ( 
.A1(n_5479),
.A2(n_5282),
.B(n_5278),
.Y(n_5767)
);

OAI21x1_ASAP7_75t_L g5768 ( 
.A1(n_5466),
.A2(n_5214),
.B(n_5170),
.Y(n_5768)
);

NAND3xp33_ASAP7_75t_L g5769 ( 
.A(n_5680),
.B(n_5266),
.C(n_5179),
.Y(n_5769)
);

OAI22xp33_ASAP7_75t_L g5770 ( 
.A1(n_5481),
.A2(n_5324),
.B1(n_5024),
.B2(n_5266),
.Y(n_5770)
);

OAI21x1_ASAP7_75t_L g5771 ( 
.A1(n_5726),
.A2(n_5123),
.B(n_5330),
.Y(n_5771)
);

NOR2xp33_ASAP7_75t_L g5772 ( 
.A(n_5489),
.B(n_5310),
.Y(n_5772)
);

CKINVDCx5p33_ASAP7_75t_R g5773 ( 
.A(n_5418),
.Y(n_5773)
);

NOR2xp67_ASAP7_75t_SL g5774 ( 
.A(n_5489),
.B(n_5345),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_5515),
.Y(n_5775)
);

AOI221xp5_ASAP7_75t_L g5776 ( 
.A1(n_5601),
.A2(n_5352),
.B1(n_5315),
.B2(n_5183),
.C(n_5146),
.Y(n_5776)
);

AO31x2_ASAP7_75t_L g5777 ( 
.A1(n_5623),
.A2(n_5357),
.A3(n_5402),
.B(n_5290),
.Y(n_5777)
);

BUFx12f_ASAP7_75t_L g5778 ( 
.A(n_5673),
.Y(n_5778)
);

NAND2x1p5_ASAP7_75t_L g5779 ( 
.A(n_5554),
.B(n_5084),
.Y(n_5779)
);

INVx1_ASAP7_75t_SL g5780 ( 
.A(n_5569),
.Y(n_5780)
);

OAI21x1_ASAP7_75t_SL g5781 ( 
.A1(n_5679),
.A2(n_5090),
.B(n_5084),
.Y(n_5781)
);

INVx2_ASAP7_75t_L g5782 ( 
.A(n_5517),
.Y(n_5782)
);

CKINVDCx11_ASAP7_75t_R g5783 ( 
.A(n_5631),
.Y(n_5783)
);

OAI22xp5_ASAP7_75t_L g5784 ( 
.A1(n_5437),
.A2(n_5475),
.B1(n_5467),
.B2(n_5493),
.Y(n_5784)
);

OAI21x1_ASAP7_75t_L g5785 ( 
.A1(n_5492),
.A2(n_5123),
.B(n_5241),
.Y(n_5785)
);

OA21x2_ASAP7_75t_L g5786 ( 
.A1(n_5727),
.A2(n_5196),
.B(n_5323),
.Y(n_5786)
);

AO21x1_ASAP7_75t_L g5787 ( 
.A1(n_5500),
.A2(n_5244),
.B(n_5352),
.Y(n_5787)
);

INVx2_ASAP7_75t_L g5788 ( 
.A(n_5517),
.Y(n_5788)
);

AOI222xp33_ASAP7_75t_L g5789 ( 
.A1(n_5733),
.A2(n_5122),
.B1(n_5183),
.B2(n_5080),
.C1(n_5315),
.C2(n_5208),
.Y(n_5789)
);

INVx2_ASAP7_75t_L g5790 ( 
.A(n_5524),
.Y(n_5790)
);

O2A1O1Ixp33_ASAP7_75t_SL g5791 ( 
.A1(n_5584),
.A2(n_5186),
.B(n_5211),
.C(n_5205),
.Y(n_5791)
);

AO21x2_ASAP7_75t_L g5792 ( 
.A1(n_5623),
.A2(n_5201),
.B(n_5250),
.Y(n_5792)
);

INVx2_ASAP7_75t_L g5793 ( 
.A(n_5524),
.Y(n_5793)
);

BUFx6f_ASAP7_75t_L g5794 ( 
.A(n_5442),
.Y(n_5794)
);

OA21x2_ASAP7_75t_L g5795 ( 
.A1(n_5727),
.A2(n_5301),
.B(n_5234),
.Y(n_5795)
);

OAI221xp5_ASAP7_75t_L g5796 ( 
.A1(n_5482),
.A2(n_5268),
.B1(n_5280),
.B2(n_5317),
.C(n_5190),
.Y(n_5796)
);

BUFx6f_ASAP7_75t_L g5797 ( 
.A(n_5442),
.Y(n_5797)
);

OAI21x1_ASAP7_75t_L g5798 ( 
.A1(n_5747),
.A2(n_5271),
.B(n_5376),
.Y(n_5798)
);

OA21x2_ASAP7_75t_L g5799 ( 
.A1(n_5746),
.A2(n_5319),
.B(n_5201),
.Y(n_5799)
);

AND2x4_ASAP7_75t_L g5800 ( 
.A(n_5620),
.B(n_5024),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5528),
.Y(n_5801)
);

AO31x2_ASAP7_75t_L g5802 ( 
.A1(n_5627),
.A2(n_5090),
.A3(n_5134),
.B(n_5132),
.Y(n_5802)
);

OA21x2_ASAP7_75t_L g5803 ( 
.A1(n_5746),
.A2(n_5379),
.B(n_5373),
.Y(n_5803)
);

INVx3_ASAP7_75t_L g5804 ( 
.A(n_5429),
.Y(n_5804)
);

OA21x2_ASAP7_75t_L g5805 ( 
.A1(n_5627),
.A2(n_5367),
.B(n_5258),
.Y(n_5805)
);

OAI21x1_ASAP7_75t_L g5806 ( 
.A1(n_5465),
.A2(n_5311),
.B(n_5388),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5528),
.Y(n_5807)
);

BUFx6f_ASAP7_75t_L g5808 ( 
.A(n_5447),
.Y(n_5808)
);

OAI21x1_ASAP7_75t_SL g5809 ( 
.A1(n_5487),
.A2(n_5134),
.B(n_5132),
.Y(n_5809)
);

AOI22xp33_ASAP7_75t_L g5810 ( 
.A1(n_5614),
.A2(n_5523),
.B1(n_5594),
.B2(n_5413),
.Y(n_5810)
);

AND2x2_ASAP7_75t_L g5811 ( 
.A(n_5610),
.B(n_5243),
.Y(n_5811)
);

OAI21x1_ASAP7_75t_L g5812 ( 
.A1(n_5744),
.A2(n_5244),
.B(n_5326),
.Y(n_5812)
);

HB1xp67_ASAP7_75t_L g5813 ( 
.A(n_5461),
.Y(n_5813)
);

OAI21x1_ASAP7_75t_L g5814 ( 
.A1(n_5678),
.A2(n_5372),
.B(n_5225),
.Y(n_5814)
);

OAI21x1_ASAP7_75t_SL g5815 ( 
.A1(n_5593),
.A2(n_5338),
.B(n_5341),
.Y(n_5815)
);

AND2x4_ASAP7_75t_L g5816 ( 
.A(n_5577),
.B(n_5069),
.Y(n_5816)
);

INVx3_ASAP7_75t_L g5817 ( 
.A(n_5441),
.Y(n_5817)
);

OAI21x1_ASAP7_75t_L g5818 ( 
.A1(n_5469),
.A2(n_5041),
.B(n_5233),
.Y(n_5818)
);

BUFx6f_ASAP7_75t_L g5819 ( 
.A(n_5447),
.Y(n_5819)
);

INVx1_ASAP7_75t_L g5820 ( 
.A(n_5530),
.Y(n_5820)
);

OAI22xp5_ASAP7_75t_L g5821 ( 
.A1(n_5446),
.A2(n_5522),
.B1(n_5480),
.B2(n_5603),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5530),
.Y(n_5822)
);

O2A1O1Ixp33_ASAP7_75t_SL g5823 ( 
.A1(n_5706),
.A2(n_5220),
.B(n_5222),
.C(n_5025),
.Y(n_5823)
);

AO21x2_ASAP7_75t_L g5824 ( 
.A1(n_5632),
.A2(n_5474),
.B(n_5622),
.Y(n_5824)
);

INVx2_ASAP7_75t_L g5825 ( 
.A(n_5531),
.Y(n_5825)
);

OAI21x1_ASAP7_75t_L g5826 ( 
.A1(n_5640),
.A2(n_5233),
.B(n_5303),
.Y(n_5826)
);

AND2x4_ASAP7_75t_L g5827 ( 
.A(n_5577),
.B(n_5069),
.Y(n_5827)
);

NAND2xp5_ASAP7_75t_L g5828 ( 
.A(n_5675),
.B(n_5074),
.Y(n_5828)
);

O2A1O1Ixp33_ASAP7_75t_L g5829 ( 
.A1(n_5698),
.A2(n_5277),
.B(n_5370),
.C(n_5346),
.Y(n_5829)
);

OR2x2_ASAP7_75t_L g5830 ( 
.A(n_5615),
.B(n_5074),
.Y(n_5830)
);

OA21x2_ASAP7_75t_L g5831 ( 
.A1(n_5632),
.A2(n_5675),
.B(n_5687),
.Y(n_5831)
);

AOI221xp5_ASAP7_75t_L g5832 ( 
.A1(n_5736),
.A2(n_5277),
.B1(n_5280),
.B2(n_5317),
.C(n_5235),
.Y(n_5832)
);

NAND2x1p5_ASAP7_75t_L g5833 ( 
.A(n_5712),
.B(n_5152),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_5531),
.Y(n_5834)
);

BUFx12f_ASAP7_75t_L g5835 ( 
.A(n_5579),
.Y(n_5835)
);

AO21x2_ASAP7_75t_L g5836 ( 
.A1(n_5506),
.A2(n_5403),
.B(n_5387),
.Y(n_5836)
);

AND2x2_ASAP7_75t_L g5837 ( 
.A(n_5420),
.B(n_5421),
.Y(n_5837)
);

INVx2_ASAP7_75t_L g5838 ( 
.A(n_5426),
.Y(n_5838)
);

OAI21x1_ASAP7_75t_L g5839 ( 
.A1(n_5557),
.A2(n_5387),
.B(n_5124),
.Y(n_5839)
);

BUFx2_ASAP7_75t_L g5840 ( 
.A(n_5511),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5427),
.Y(n_5841)
);

INVx3_ASAP7_75t_L g5842 ( 
.A(n_5441),
.Y(n_5842)
);

AOI21x1_ASAP7_75t_L g5843 ( 
.A1(n_5695),
.A2(n_5342),
.B(n_5154),
.Y(n_5843)
);

O2A1O1Ixp33_ASAP7_75t_SL g5844 ( 
.A1(n_5563),
.A2(n_5124),
.B(n_5089),
.C(n_5345),
.Y(n_5844)
);

NOR2xp33_ASAP7_75t_SL g5845 ( 
.A(n_5509),
.B(n_5377),
.Y(n_5845)
);

INVx6_ASAP7_75t_SL g5846 ( 
.A(n_5613),
.Y(n_5846)
);

NOR2x1_ASAP7_75t_SL g5847 ( 
.A(n_5454),
.B(n_5377),
.Y(n_5847)
);

INVx1_ASAP7_75t_SL g5848 ( 
.A(n_5697),
.Y(n_5848)
);

BUFx3_ASAP7_75t_L g5849 ( 
.A(n_5690),
.Y(n_5849)
);

INVx2_ASAP7_75t_L g5850 ( 
.A(n_5582),
.Y(n_5850)
);

AO21x2_ASAP7_75t_L g5851 ( 
.A1(n_5476),
.A2(n_5342),
.B(n_5154),
.Y(n_5851)
);

NOR2xp33_ASAP7_75t_L g5852 ( 
.A(n_5737),
.B(n_5377),
.Y(n_5852)
);

INVx1_ASAP7_75t_SL g5853 ( 
.A(n_5473),
.Y(n_5853)
);

AND2x2_ASAP7_75t_L g5854 ( 
.A(n_5494),
.B(n_5074),
.Y(n_5854)
);

INVx2_ASAP7_75t_SL g5855 ( 
.A(n_5516),
.Y(n_5855)
);

OAI21x1_ASAP7_75t_L g5856 ( 
.A1(n_5519),
.A2(n_2558),
.B(n_2531),
.Y(n_5856)
);

OAI21xp5_ASAP7_75t_L g5857 ( 
.A1(n_5419),
.A2(n_5654),
.B(n_5411),
.Y(n_5857)
);

INVx2_ASAP7_75t_L g5858 ( 
.A(n_5582),
.Y(n_5858)
);

AO21x2_ASAP7_75t_L g5859 ( 
.A1(n_5550),
.A2(n_5203),
.B(n_5152),
.Y(n_5859)
);

INVx2_ASAP7_75t_L g5860 ( 
.A(n_5592),
.Y(n_5860)
);

NOR2x1_ASAP7_75t_R g5861 ( 
.A(n_5417),
.B(n_5433),
.Y(n_5861)
);

HB1xp67_ASAP7_75t_L g5862 ( 
.A(n_5521),
.Y(n_5862)
);

OAI22xp33_ASAP7_75t_L g5863 ( 
.A1(n_5738),
.A2(n_5177),
.B1(n_5215),
.B2(n_5192),
.Y(n_5863)
);

OAI21x1_ASAP7_75t_L g5864 ( 
.A1(n_5425),
.A2(n_5504),
.B(n_5553),
.Y(n_5864)
);

NAND2xp5_ASAP7_75t_L g5865 ( 
.A(n_5685),
.B(n_5177),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5439),
.Y(n_5866)
);

INVx2_ASAP7_75t_L g5867 ( 
.A(n_5592),
.Y(n_5867)
);

INVx2_ASAP7_75t_L g5868 ( 
.A(n_5534),
.Y(n_5868)
);

AOI22xp33_ASAP7_75t_L g5869 ( 
.A1(n_5669),
.A2(n_5110),
.B1(n_5253),
.B2(n_5203),
.Y(n_5869)
);

INVx2_ASAP7_75t_L g5870 ( 
.A(n_5443),
.Y(n_5870)
);

OR2x6_ASAP7_75t_L g5871 ( 
.A(n_5454),
.B(n_5253),
.Y(n_5871)
);

BUFx8_ASAP7_75t_L g5872 ( 
.A(n_5571),
.Y(n_5872)
);

OAI21xp5_ASAP7_75t_L g5873 ( 
.A1(n_5545),
.A2(n_5412),
.B(n_5478),
.Y(n_5873)
);

NAND2xp5_ASAP7_75t_L g5874 ( 
.A(n_5541),
.B(n_5177),
.Y(n_5874)
);

HB1xp67_ASAP7_75t_L g5875 ( 
.A(n_5535),
.Y(n_5875)
);

AOI22xp33_ASAP7_75t_L g5876 ( 
.A1(n_5463),
.A2(n_5110),
.B1(n_5276),
.B2(n_5215),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_5444),
.Y(n_5877)
);

INVx1_ASAP7_75t_L g5878 ( 
.A(n_5450),
.Y(n_5878)
);

OR2x2_ASAP7_75t_L g5879 ( 
.A(n_5423),
.B(n_5424),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_5451),
.Y(n_5880)
);

AND2x4_ASAP7_75t_L g5881 ( 
.A(n_5607),
.B(n_5192),
.Y(n_5881)
);

AND2x2_ASAP7_75t_L g5882 ( 
.A(n_5453),
.B(n_5192),
.Y(n_5882)
);

NAND2xp5_ASAP7_75t_L g5883 ( 
.A(n_5587),
.B(n_5215),
.Y(n_5883)
);

OAI21x1_ASAP7_75t_L g5884 ( 
.A1(n_5691),
.A2(n_2558),
.B(n_2531),
.Y(n_5884)
);

INVx2_ASAP7_75t_SL g5885 ( 
.A(n_5499),
.Y(n_5885)
);

O2A1O1Ixp33_ASAP7_75t_L g5886 ( 
.A1(n_5742),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_5886)
);

INVx1_ASAP7_75t_L g5887 ( 
.A(n_5496),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_5498),
.Y(n_5888)
);

INVx1_ASAP7_75t_L g5889 ( 
.A(n_5503),
.Y(n_5889)
);

BUFx12f_ASAP7_75t_L g5890 ( 
.A(n_5636),
.Y(n_5890)
);

AOI21xp5_ASAP7_75t_L g5891 ( 
.A1(n_5684),
.A2(n_5362),
.B(n_5227),
.Y(n_5891)
);

AO21x2_ASAP7_75t_L g5892 ( 
.A1(n_5642),
.A2(n_5110),
.B(n_5221),
.Y(n_5892)
);

AOI221xp5_ASAP7_75t_L g5893 ( 
.A1(n_5724),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.C(n_40),
.Y(n_5893)
);

OR2x6_ASAP7_75t_L g5894 ( 
.A(n_5484),
.B(n_5221),
.Y(n_5894)
);

BUFx3_ASAP7_75t_L g5895 ( 
.A(n_5591),
.Y(n_5895)
);

AO21x2_ASAP7_75t_L g5896 ( 
.A1(n_5422),
.A2(n_5223),
.B(n_5221),
.Y(n_5896)
);

BUFx2_ASAP7_75t_L g5897 ( 
.A(n_5455),
.Y(n_5897)
);

OR2x2_ASAP7_75t_L g5898 ( 
.A(n_5428),
.B(n_5223),
.Y(n_5898)
);

OAI21x1_ASAP7_75t_L g5899 ( 
.A1(n_5743),
.A2(n_2558),
.B(n_2531),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5507),
.Y(n_5900)
);

OAI21xp5_ASAP7_75t_L g5901 ( 
.A1(n_5432),
.A2(n_39),
.B(n_40),
.Y(n_5901)
);

INVx4_ASAP7_75t_SL g5902 ( 
.A(n_5643),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5543),
.Y(n_5903)
);

INVx6_ASAP7_75t_L g5904 ( 
.A(n_5536),
.Y(n_5904)
);

OR2x2_ASAP7_75t_L g5905 ( 
.A(n_5430),
.B(n_5223),
.Y(n_5905)
);

AND2x2_ASAP7_75t_L g5906 ( 
.A(n_5512),
.B(n_5263),
.Y(n_5906)
);

OR2x2_ASAP7_75t_L g5907 ( 
.A(n_5483),
.B(n_5263),
.Y(n_5907)
);

INVx2_ASAP7_75t_L g5908 ( 
.A(n_5689),
.Y(n_5908)
);

INVx1_ASAP7_75t_L g5909 ( 
.A(n_5533),
.Y(n_5909)
);

OAI22xp5_ASAP7_75t_L g5910 ( 
.A1(n_5585),
.A2(n_5265),
.B1(n_5273),
.B2(n_5263),
.Y(n_5910)
);

OAI21x1_ASAP7_75t_L g5911 ( 
.A1(n_5588),
.A2(n_2614),
.B(n_2600),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5562),
.Y(n_5912)
);

OR2x6_ASAP7_75t_L g5913 ( 
.A(n_5484),
.B(n_5265),
.Y(n_5913)
);

OR2x2_ASAP7_75t_L g5914 ( 
.A(n_5501),
.B(n_5265),
.Y(n_5914)
);

AND2x4_ASAP7_75t_L g5915 ( 
.A(n_5607),
.B(n_5273),
.Y(n_5915)
);

NAND2x1p5_ASAP7_75t_L g5916 ( 
.A(n_5712),
.B(n_5273),
.Y(n_5916)
);

INVx3_ASAP7_75t_L g5917 ( 
.A(n_5472),
.Y(n_5917)
);

OAI21xp5_ASAP7_75t_L g5918 ( 
.A1(n_5576),
.A2(n_41),
.B(n_42),
.Y(n_5918)
);

AOI22xp5_ASAP7_75t_L g5919 ( 
.A1(n_5667),
.A2(n_5327),
.B1(n_5329),
.B2(n_2587),
.Y(n_5919)
);

OAI21x1_ASAP7_75t_L g5920 ( 
.A1(n_5588),
.A2(n_5626),
.B(n_5619),
.Y(n_5920)
);

INVx2_ASAP7_75t_L g5921 ( 
.A(n_5570),
.Y(n_5921)
);

OAI21x1_ASAP7_75t_L g5922 ( 
.A1(n_5619),
.A2(n_5649),
.B(n_5626),
.Y(n_5922)
);

AOI22xp33_ASAP7_75t_L g5923 ( 
.A1(n_5463),
.A2(n_5495),
.B1(n_5692),
.B2(n_5596),
.Y(n_5923)
);

AND2x2_ASAP7_75t_L g5924 ( 
.A(n_5551),
.B(n_5327),
.Y(n_5924)
);

AOI22xp33_ASAP7_75t_L g5925 ( 
.A1(n_5495),
.A2(n_5327),
.B1(n_5329),
.B2(n_2587),
.Y(n_5925)
);

A2O1A1Ixp33_ASAP7_75t_L g5926 ( 
.A1(n_5739),
.A2(n_5329),
.B(n_46),
.C(n_49),
.Y(n_5926)
);

INVx4_ASAP7_75t_SL g5927 ( 
.A(n_5571),
.Y(n_5927)
);

OAI21x1_ASAP7_75t_L g5928 ( 
.A1(n_5649),
.A2(n_3105),
.B(n_3089),
.Y(n_5928)
);

INVx1_ASAP7_75t_L g5929 ( 
.A(n_5573),
.Y(n_5929)
);

CKINVDCx5p33_ASAP7_75t_R g5930 ( 
.A(n_5683),
.Y(n_5930)
);

AOI21xp5_ASAP7_75t_L g5931 ( 
.A1(n_5502),
.A2(n_3374),
.B(n_3367),
.Y(n_5931)
);

HB1xp67_ASAP7_75t_L g5932 ( 
.A(n_5435),
.Y(n_5932)
);

AND2x4_ASAP7_75t_L g5933 ( 
.A(n_5472),
.B(n_43),
.Y(n_5933)
);

INVx2_ASAP7_75t_L g5934 ( 
.A(n_5600),
.Y(n_5934)
);

CKINVDCx5p33_ASAP7_75t_R g5935 ( 
.A(n_5741),
.Y(n_5935)
);

NAND2xp5_ASAP7_75t_L g5936 ( 
.A(n_5505),
.B(n_44),
.Y(n_5936)
);

OAI21x1_ASAP7_75t_L g5937 ( 
.A1(n_5707),
.A2(n_3105),
.B(n_3089),
.Y(n_5937)
);

CKINVDCx20_ASAP7_75t_R g5938 ( 
.A(n_5438),
.Y(n_5938)
);

INVx2_ASAP7_75t_L g5939 ( 
.A(n_5605),
.Y(n_5939)
);

INVx1_ASAP7_75t_L g5940 ( 
.A(n_5575),
.Y(n_5940)
);

AND2x6_ASAP7_75t_L g5941 ( 
.A(n_5723),
.B(n_3367),
.Y(n_5941)
);

OAI21x1_ASAP7_75t_L g5942 ( 
.A1(n_5641),
.A2(n_5609),
.B(n_5705),
.Y(n_5942)
);

OAI21x1_ASAP7_75t_L g5943 ( 
.A1(n_5462),
.A2(n_3128),
.B(n_2919),
.Y(n_5943)
);

INVx2_ASAP7_75t_L g5944 ( 
.A(n_5414),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5581),
.Y(n_5945)
);

A2O1A1Ixp33_ASAP7_75t_L g5946 ( 
.A1(n_5650),
.A2(n_54),
.B(n_55),
.C(n_51),
.Y(n_5946)
);

BUFx12f_ASAP7_75t_L g5947 ( 
.A(n_5571),
.Y(n_5947)
);

AO21x2_ASAP7_75t_L g5948 ( 
.A1(n_5560),
.A2(n_2950),
.B(n_2949),
.Y(n_5948)
);

OAI21x1_ASAP7_75t_L g5949 ( 
.A1(n_5468),
.A2(n_2933),
.B(n_2914),
.Y(n_5949)
);

INVx6_ASAP7_75t_L g5950 ( 
.A(n_5536),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5604),
.Y(n_5951)
);

AOI22xp33_ASAP7_75t_L g5952 ( 
.A1(n_5715),
.A2(n_2224),
.B1(n_2226),
.B2(n_2219),
.Y(n_5952)
);

AND2x2_ASAP7_75t_L g5953 ( 
.A(n_5555),
.B(n_50),
.Y(n_5953)
);

OAI21xp5_ASAP7_75t_L g5954 ( 
.A1(n_5710),
.A2(n_50),
.B(n_51),
.Y(n_5954)
);

CKINVDCx5p33_ASAP7_75t_R g5955 ( 
.A(n_5558),
.Y(n_5955)
);

INVx2_ASAP7_75t_L g5956 ( 
.A(n_5431),
.Y(n_5956)
);

NOR2xp67_ASAP7_75t_L g5957 ( 
.A(n_5712),
.B(n_56),
.Y(n_5957)
);

AND2x4_ASAP7_75t_L g5958 ( 
.A(n_5505),
.B(n_57),
.Y(n_5958)
);

AND2x2_ASAP7_75t_L g5959 ( 
.A(n_5586),
.B(n_58),
.Y(n_5959)
);

OA21x2_ASAP7_75t_L g5960 ( 
.A1(n_5520),
.A2(n_5572),
.B(n_5448),
.Y(n_5960)
);

AOI22xp33_ASAP7_75t_L g5961 ( 
.A1(n_5702),
.A2(n_5633),
.B1(n_5718),
.B2(n_5653),
.Y(n_5961)
);

AO21x2_ASAP7_75t_L g5962 ( 
.A1(n_5604),
.A2(n_2950),
.B(n_2949),
.Y(n_5962)
);

AND2x2_ASAP7_75t_L g5963 ( 
.A(n_5602),
.B(n_58),
.Y(n_5963)
);

NOR2x1_ASAP7_75t_SL g5964 ( 
.A(n_5502),
.B(n_1250),
.Y(n_5964)
);

AOI21x1_ASAP7_75t_L g5965 ( 
.A1(n_5590),
.A2(n_2948),
.B(n_2935),
.Y(n_5965)
);

INVx2_ASAP7_75t_L g5966 ( 
.A(n_5434),
.Y(n_5966)
);

INVx2_ASAP7_75t_L g5967 ( 
.A(n_5445),
.Y(n_5967)
);

INVx3_ASAP7_75t_L g5968 ( 
.A(n_5470),
.Y(n_5968)
);

BUFx6f_ASAP7_75t_L g5969 ( 
.A(n_5447),
.Y(n_5969)
);

AND2x4_ASAP7_75t_L g5970 ( 
.A(n_5416),
.B(n_59),
.Y(n_5970)
);

AO21x2_ASAP7_75t_L g5971 ( 
.A1(n_5606),
.A2(n_5612),
.B(n_5676),
.Y(n_5971)
);

OAI21x1_ASAP7_75t_SL g5972 ( 
.A1(n_5542),
.A2(n_59),
.B(n_60),
.Y(n_5972)
);

AOI21xp33_ASAP7_75t_SL g5973 ( 
.A1(n_5694),
.A2(n_61),
.B(n_62),
.Y(n_5973)
);

OAI21x1_ASAP7_75t_L g5974 ( 
.A1(n_5470),
.A2(n_2948),
.B(n_2935),
.Y(n_5974)
);

INVx2_ASAP7_75t_L g5975 ( 
.A(n_5514),
.Y(n_5975)
);

NAND2xp5_ASAP7_75t_L g5976 ( 
.A(n_5548),
.B(n_62),
.Y(n_5976)
);

AO31x2_ASAP7_75t_L g5977 ( 
.A1(n_5703),
.A2(n_65),
.A3(n_63),
.B(n_64),
.Y(n_5977)
);

CKINVDCx5p33_ASAP7_75t_R g5978 ( 
.A(n_5634),
.Y(n_5978)
);

INVx4_ASAP7_75t_L g5979 ( 
.A(n_5696),
.Y(n_5979)
);

CKINVDCx20_ASAP7_75t_R g5980 ( 
.A(n_5440),
.Y(n_5980)
);

AO21x2_ASAP7_75t_L g5981 ( 
.A1(n_5566),
.A2(n_2944),
.B(n_77),
.Y(n_5981)
);

NOR2xp33_ASAP7_75t_L g5982 ( 
.A(n_5497),
.B(n_66),
.Y(n_5982)
);

OAI21x1_ASAP7_75t_L g5983 ( 
.A1(n_5486),
.A2(n_2951),
.B(n_2944),
.Y(n_5983)
);

OAI21x1_ASAP7_75t_L g5984 ( 
.A1(n_5486),
.A2(n_2951),
.B(n_2769),
.Y(n_5984)
);

INVx1_ASAP7_75t_SL g5985 ( 
.A(n_5719),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5518),
.Y(n_5986)
);

OAI21x1_ASAP7_75t_L g5987 ( 
.A1(n_5488),
.A2(n_2951),
.B(n_2769),
.Y(n_5987)
);

OA21x2_ASAP7_75t_L g5988 ( 
.A1(n_5526),
.A2(n_2673),
.B(n_2668),
.Y(n_5988)
);

OA21x2_ASAP7_75t_L g5989 ( 
.A1(n_5547),
.A2(n_2680),
.B(n_2676),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5527),
.Y(n_5990)
);

NAND2xp5_ASAP7_75t_L g5991 ( 
.A(n_5617),
.B(n_66),
.Y(n_5991)
);

CKINVDCx5p33_ASAP7_75t_R g5992 ( 
.A(n_5731),
.Y(n_5992)
);

AO21x2_ASAP7_75t_L g5993 ( 
.A1(n_5668),
.A2(n_79),
.B(n_68),
.Y(n_5993)
);

INVx1_ASAP7_75t_L g5994 ( 
.A(n_5644),
.Y(n_5994)
);

NOR3xp33_ASAP7_75t_SL g5995 ( 
.A(n_5595),
.B(n_68),
.C(n_69),
.Y(n_5995)
);

INVx2_ASAP7_75t_L g5996 ( 
.A(n_5677),
.Y(n_5996)
);

NOR2xp33_ASAP7_75t_L g5997 ( 
.A(n_5497),
.B(n_5637),
.Y(n_5997)
);

OAI21x1_ASAP7_75t_L g5998 ( 
.A1(n_5488),
.A2(n_2769),
.B(n_2763),
.Y(n_5998)
);

O2A1O1Ixp33_ASAP7_75t_L g5999 ( 
.A1(n_5716),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_5999)
);

A2O1A1Ixp33_ASAP7_75t_L g6000 ( 
.A1(n_5723),
.A2(n_75),
.B(n_77),
.C(n_73),
.Y(n_6000)
);

AOI21xp5_ASAP7_75t_L g6001 ( 
.A1(n_5580),
.A2(n_3374),
.B(n_3367),
.Y(n_6001)
);

AO31x2_ASAP7_75t_L g6002 ( 
.A1(n_5740),
.A2(n_79),
.A3(n_72),
.B(n_73),
.Y(n_6002)
);

OA21x2_ASAP7_75t_L g6003 ( 
.A1(n_5699),
.A2(n_2681),
.B(n_2680),
.Y(n_6003)
);

NOR2xp33_ASAP7_75t_SL g6004 ( 
.A(n_5580),
.B(n_5552),
.Y(n_6004)
);

NAND2xp5_ASAP7_75t_L g6005 ( 
.A(n_5646),
.B(n_80),
.Y(n_6005)
);

INVx2_ASAP7_75t_L g6006 ( 
.A(n_5682),
.Y(n_6006)
);

AOI22xp33_ASAP7_75t_L g6007 ( 
.A1(n_5633),
.A2(n_2227),
.B1(n_2226),
.B2(n_2964),
.Y(n_6007)
);

INVx2_ASAP7_75t_L g6008 ( 
.A(n_5686),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5647),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5651),
.Y(n_6010)
);

O2A1O1Ixp33_ASAP7_75t_SL g6011 ( 
.A1(n_5564),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_6011)
);

AOI22xp33_ASAP7_75t_L g6012 ( 
.A1(n_5653),
.A2(n_2227),
.B1(n_2226),
.B2(n_2964),
.Y(n_6012)
);

NAND2xp5_ASAP7_75t_L g6013 ( 
.A(n_5652),
.B(n_83),
.Y(n_6013)
);

OA21x2_ASAP7_75t_L g6014 ( 
.A1(n_5711),
.A2(n_2683),
.B(n_2681),
.Y(n_6014)
);

NOR2x1_ASAP7_75t_L g6015 ( 
.A(n_5459),
.B(n_3374),
.Y(n_6015)
);

AOI21xp5_ASAP7_75t_L g6016 ( 
.A1(n_5552),
.A2(n_3381),
.B(n_3374),
.Y(n_6016)
);

OR2x6_ASAP7_75t_L g6017 ( 
.A(n_5613),
.B(n_3381),
.Y(n_6017)
);

HB1xp67_ASAP7_75t_L g6018 ( 
.A(n_5459),
.Y(n_6018)
);

BUFx2_ASAP7_75t_L g6019 ( 
.A(n_5455),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_5657),
.Y(n_6020)
);

NAND2x1p5_ASAP7_75t_L g6021 ( 
.A(n_6015),
.B(n_5539),
.Y(n_6021)
);

OAI21xp5_ASAP7_75t_L g6022 ( 
.A1(n_5857),
.A2(n_5873),
.B(n_5901),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_5751),
.Y(n_6023)
);

INVx1_ASAP7_75t_L g6024 ( 
.A(n_5759),
.Y(n_6024)
);

BUFx3_ASAP7_75t_L g6025 ( 
.A(n_5778),
.Y(n_6025)
);

OR2x2_ASAP7_75t_L g6026 ( 
.A(n_5780),
.B(n_5491),
.Y(n_6026)
);

INVx2_ASAP7_75t_L g6027 ( 
.A(n_5896),
.Y(n_6027)
);

INVx4_ASAP7_75t_L g6028 ( 
.A(n_5902),
.Y(n_6028)
);

NAND2xp5_ASAP7_75t_L g6029 ( 
.A(n_5960),
.B(n_5659),
.Y(n_6029)
);

INVx2_ASAP7_75t_L g6030 ( 
.A(n_5850),
.Y(n_6030)
);

INVx1_ASAP7_75t_L g6031 ( 
.A(n_5951),
.Y(n_6031)
);

AOI22xp33_ASAP7_75t_SL g6032 ( 
.A1(n_5901),
.A2(n_5725),
.B1(n_5734),
.B2(n_5729),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_5761),
.Y(n_6033)
);

HB1xp67_ASAP7_75t_L g6034 ( 
.A(n_5960),
.Y(n_6034)
);

AOI22xp33_ASAP7_75t_L g6035 ( 
.A1(n_5857),
.A2(n_5455),
.B1(n_5599),
.B2(n_5725),
.Y(n_6035)
);

AOI22xp33_ASAP7_75t_L g6036 ( 
.A1(n_5787),
.A2(n_5734),
.B1(n_5497),
.B2(n_5701),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_5775),
.Y(n_6037)
);

BUFx4_ASAP7_75t_SL g6038 ( 
.A(n_5935),
.Y(n_6038)
);

OR2x2_ASAP7_75t_L g6039 ( 
.A(n_5780),
.B(n_5508),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5807),
.Y(n_6040)
);

INVx5_ASAP7_75t_SL g6041 ( 
.A(n_5993),
.Y(n_6041)
);

CKINVDCx5p33_ASAP7_75t_R g6042 ( 
.A(n_5783),
.Y(n_6042)
);

INVx1_ASAP7_75t_L g6043 ( 
.A(n_5820),
.Y(n_6043)
);

OAI22xp33_ASAP7_75t_L g6044 ( 
.A1(n_5873),
.A2(n_5753),
.B1(n_5754),
.B2(n_6004),
.Y(n_6044)
);

BUFx10_ASAP7_75t_L g6045 ( 
.A(n_5982),
.Y(n_6045)
);

AOI22xp33_ASAP7_75t_L g6046 ( 
.A1(n_5769),
.A2(n_5416),
.B1(n_5540),
.B2(n_5745),
.Y(n_6046)
);

BUFx5_ASAP7_75t_L g6047 ( 
.A(n_5941),
.Y(n_6047)
);

INVx2_ASAP7_75t_L g6048 ( 
.A(n_5858),
.Y(n_6048)
);

INVx2_ASAP7_75t_L g6049 ( 
.A(n_5860),
.Y(n_6049)
);

NAND2xp5_ASAP7_75t_L g6050 ( 
.A(n_5971),
.B(n_5660),
.Y(n_6050)
);

AND2x2_ASAP7_75t_L g6051 ( 
.A(n_5762),
.B(n_5436),
.Y(n_6051)
);

CKINVDCx20_ASAP7_75t_R g6052 ( 
.A(n_5980),
.Y(n_6052)
);

NAND2xp5_ASAP7_75t_SL g6053 ( 
.A(n_5845),
.B(n_5449),
.Y(n_6053)
);

OAI22xp33_ASAP7_75t_L g6054 ( 
.A1(n_5753),
.A2(n_5713),
.B1(n_5681),
.B2(n_5720),
.Y(n_6054)
);

INVx4_ASAP7_75t_SL g6055 ( 
.A(n_5977),
.Y(n_6055)
);

NOR2xp33_ASAP7_75t_L g6056 ( 
.A(n_5979),
.B(n_5490),
.Y(n_6056)
);

INVx2_ASAP7_75t_L g6057 ( 
.A(n_5867),
.Y(n_6057)
);

AND2x4_ASAP7_75t_L g6058 ( 
.A(n_5840),
.B(n_5529),
.Y(n_6058)
);

NAND2xp5_ASAP7_75t_L g6059 ( 
.A(n_5971),
.B(n_5635),
.Y(n_6059)
);

INVx1_ASAP7_75t_L g6060 ( 
.A(n_5822),
.Y(n_6060)
);

INVx2_ASAP7_75t_L g6061 ( 
.A(n_5782),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_5834),
.Y(n_6062)
);

INVx2_ASAP7_75t_SL g6063 ( 
.A(n_5904),
.Y(n_6063)
);

AOI22xp33_ASAP7_75t_L g6064 ( 
.A1(n_5769),
.A2(n_5810),
.B1(n_5954),
.B2(n_5754),
.Y(n_6064)
);

OR2x2_ASAP7_75t_L g6065 ( 
.A(n_5879),
.B(n_5629),
.Y(n_6065)
);

AOI22xp33_ASAP7_75t_L g6066 ( 
.A1(n_5954),
.A2(n_5540),
.B1(n_5714),
.B2(n_5648),
.Y(n_6066)
);

INVx1_ASAP7_75t_L g6067 ( 
.A(n_5841),
.Y(n_6067)
);

INVx1_ASAP7_75t_L g6068 ( 
.A(n_5866),
.Y(n_6068)
);

OR2x6_ASAP7_75t_L g6069 ( 
.A(n_5864),
.B(n_5713),
.Y(n_6069)
);

OAI22xp5_ASAP7_75t_L g6070 ( 
.A1(n_5752),
.A2(n_5611),
.B1(n_5665),
.B2(n_5722),
.Y(n_6070)
);

INVx8_ASAP7_75t_L g6071 ( 
.A(n_5947),
.Y(n_6071)
);

INVxp67_ASAP7_75t_SL g6072 ( 
.A(n_5831),
.Y(n_6072)
);

INVx2_ASAP7_75t_L g6073 ( 
.A(n_5788),
.Y(n_6073)
);

AO21x2_ASAP7_75t_L g6074 ( 
.A1(n_5824),
.A2(n_5574),
.B(n_5645),
.Y(n_6074)
);

AOI22xp33_ASAP7_75t_L g6075 ( 
.A1(n_5789),
.A2(n_5540),
.B1(n_5648),
.B2(n_5638),
.Y(n_6075)
);

AOI22xp33_ASAP7_75t_SL g6076 ( 
.A1(n_5918),
.A2(n_5540),
.B1(n_5578),
.B2(n_5561),
.Y(n_6076)
);

INVx2_ASAP7_75t_L g6077 ( 
.A(n_5790),
.Y(n_6077)
);

CKINVDCx5p33_ASAP7_75t_R g6078 ( 
.A(n_5773),
.Y(n_6078)
);

HB1xp67_ASAP7_75t_L g6079 ( 
.A(n_5813),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_5877),
.Y(n_6080)
);

AND2x2_ASAP7_75t_L g6081 ( 
.A(n_5917),
.B(n_5837),
.Y(n_6081)
);

HB1xp67_ASAP7_75t_L g6082 ( 
.A(n_5831),
.Y(n_6082)
);

OAI21x1_ASAP7_75t_L g6083 ( 
.A1(n_5843),
.A2(n_5549),
.B(n_5655),
.Y(n_6083)
);

BUFx8_ASAP7_75t_L g6084 ( 
.A(n_5835),
.Y(n_6084)
);

CKINVDCx5p33_ASAP7_75t_R g6085 ( 
.A(n_5890),
.Y(n_6085)
);

AOI22xp33_ASAP7_75t_L g6086 ( 
.A1(n_5789),
.A2(n_5638),
.B1(n_5529),
.B2(n_5656),
.Y(n_6086)
);

AOI22xp33_ASAP7_75t_SL g6087 ( 
.A1(n_5918),
.A2(n_5532),
.B1(n_5556),
.B2(n_5544),
.Y(n_6087)
);

CKINVDCx20_ASAP7_75t_R g6088 ( 
.A(n_5938),
.Y(n_6088)
);

BUFx2_ASAP7_75t_L g6089 ( 
.A(n_5846),
.Y(n_6089)
);

INVx2_ASAP7_75t_L g6090 ( 
.A(n_5793),
.Y(n_6090)
);

INVx2_ASAP7_75t_L g6091 ( 
.A(n_5801),
.Y(n_6091)
);

NAND2xp5_ASAP7_75t_L g6092 ( 
.A(n_5942),
.B(n_5661),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_5878),
.Y(n_6093)
);

OAI22xp33_ASAP7_75t_L g6094 ( 
.A1(n_6004),
.A2(n_5525),
.B1(n_5625),
.B2(n_5567),
.Y(n_6094)
);

BUFx3_ASAP7_75t_L g6095 ( 
.A(n_5872),
.Y(n_6095)
);

AND2x4_ASAP7_75t_L g6096 ( 
.A(n_5859),
.B(n_5693),
.Y(n_6096)
);

INVx1_ASAP7_75t_L g6097 ( 
.A(n_5880),
.Y(n_6097)
);

BUFx10_ASAP7_75t_L g6098 ( 
.A(n_5978),
.Y(n_6098)
);

INVx1_ASAP7_75t_L g6099 ( 
.A(n_5887),
.Y(n_6099)
);

INVx2_ASAP7_75t_L g6100 ( 
.A(n_5825),
.Y(n_6100)
);

INVx1_ASAP7_75t_L g6101 ( 
.A(n_5888),
.Y(n_6101)
);

INVx2_ASAP7_75t_L g6102 ( 
.A(n_5968),
.Y(n_6102)
);

OAI21x1_ASAP7_75t_L g6103 ( 
.A1(n_5771),
.A2(n_5922),
.B(n_5920),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5889),
.Y(n_6104)
);

NAND2x1p5_ASAP7_75t_L g6105 ( 
.A(n_6015),
.B(n_5539),
.Y(n_6105)
);

AOI21x1_ASAP7_75t_L g6106 ( 
.A1(n_5774),
.A2(n_5583),
.B(n_5565),
.Y(n_6106)
);

INVx4_ASAP7_75t_L g6107 ( 
.A(n_5902),
.Y(n_6107)
);

INVx1_ASAP7_75t_L g6108 ( 
.A(n_5900),
.Y(n_6108)
);

AOI22xp33_ASAP7_75t_L g6109 ( 
.A1(n_5836),
.A2(n_5688),
.B1(n_5656),
.B2(n_5721),
.Y(n_6109)
);

INVx1_ASAP7_75t_L g6110 ( 
.A(n_5903),
.Y(n_6110)
);

AOI22xp33_ASAP7_75t_SL g6111 ( 
.A1(n_5796),
.A2(n_5415),
.B1(n_5538),
.B2(n_5616),
.Y(n_6111)
);

AO21x2_ASAP7_75t_L g6112 ( 
.A1(n_5824),
.A2(n_5664),
.B(n_5663),
.Y(n_6112)
);

INVx3_ASAP7_75t_L g6113 ( 
.A(n_5846),
.Y(n_6113)
);

BUFx2_ASAP7_75t_L g6114 ( 
.A(n_5779),
.Y(n_6114)
);

AND2x4_ASAP7_75t_L g6115 ( 
.A(n_5859),
.B(n_5700),
.Y(n_6115)
);

INVx2_ASAP7_75t_L g6116 ( 
.A(n_5968),
.Y(n_6116)
);

INVx2_ASAP7_75t_L g6117 ( 
.A(n_5765),
.Y(n_6117)
);

AOI22xp33_ASAP7_75t_SL g6118 ( 
.A1(n_5796),
.A2(n_5538),
.B1(n_5721),
.B2(n_5589),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5868),
.Y(n_6119)
);

INVx1_ASAP7_75t_SL g6120 ( 
.A(n_5985),
.Y(n_6120)
);

AND2x4_ASAP7_75t_L g6121 ( 
.A(n_5847),
.B(n_5688),
.Y(n_6121)
);

AND2x2_ASAP7_75t_L g6122 ( 
.A(n_5917),
.B(n_5568),
.Y(n_6122)
);

INVx4_ASAP7_75t_L g6123 ( 
.A(n_5927),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_5870),
.Y(n_6124)
);

INVx1_ASAP7_75t_L g6125 ( 
.A(n_5929),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5940),
.Y(n_6126)
);

INVx1_ASAP7_75t_L g6127 ( 
.A(n_5945),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_5909),
.Y(n_6128)
);

HB1xp67_ASAP7_75t_L g6129 ( 
.A(n_5862),
.Y(n_6129)
);

AOI22xp33_ASAP7_75t_L g6130 ( 
.A1(n_5836),
.A2(n_5546),
.B1(n_5662),
.B2(n_5618),
.Y(n_6130)
);

INVx4_ASAP7_75t_L g6131 ( 
.A(n_5927),
.Y(n_6131)
);

BUFx2_ASAP7_75t_SL g6132 ( 
.A(n_5957),
.Y(n_6132)
);

INVx2_ASAP7_75t_L g6133 ( 
.A(n_5765),
.Y(n_6133)
);

AOI22xp33_ASAP7_75t_L g6134 ( 
.A1(n_5776),
.A2(n_5658),
.B1(n_5639),
.B2(n_5628),
.Y(n_6134)
);

BUFx2_ASAP7_75t_L g6135 ( 
.A(n_5779),
.Y(n_6135)
);

AOI22xp33_ASAP7_75t_SL g6136 ( 
.A1(n_5786),
.A2(n_5538),
.B1(n_5537),
.B2(n_5510),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_5994),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_6009),
.Y(n_6138)
);

INVx2_ASAP7_75t_SL g6139 ( 
.A(n_5904),
.Y(n_6139)
);

AOI21x1_ASAP7_75t_L g6140 ( 
.A1(n_5976),
.A2(n_5666),
.B(n_5621),
.Y(n_6140)
);

OAI22xp5_ASAP7_75t_L g6141 ( 
.A1(n_5946),
.A2(n_5670),
.B1(n_5709),
.B2(n_5672),
.Y(n_6141)
);

AOI22xp33_ASAP7_75t_L g6142 ( 
.A1(n_5776),
.A2(n_5537),
.B1(n_5559),
.B2(n_5510),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_6010),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_6020),
.Y(n_6144)
);

INVx1_ASAP7_75t_SL g6145 ( 
.A(n_5985),
.Y(n_6145)
);

AOI22xp5_ASAP7_75t_L g6146 ( 
.A1(n_5893),
.A2(n_5732),
.B1(n_5538),
.B2(n_5537),
.Y(n_6146)
);

INVx2_ASAP7_75t_L g6147 ( 
.A(n_5804),
.Y(n_6147)
);

AND2x2_ASAP7_75t_L g6148 ( 
.A(n_6018),
.B(n_5510),
.Y(n_6148)
);

INVx2_ASAP7_75t_L g6149 ( 
.A(n_5817),
.Y(n_6149)
);

CKINVDCx11_ASAP7_75t_R g6150 ( 
.A(n_5849),
.Y(n_6150)
);

INVx2_ASAP7_75t_L g6151 ( 
.A(n_5817),
.Y(n_6151)
);

HB1xp67_ASAP7_75t_SL g6152 ( 
.A(n_5872),
.Y(n_6152)
);

INVx2_ASAP7_75t_L g6153 ( 
.A(n_5842),
.Y(n_6153)
);

INVx2_ASAP7_75t_L g6154 ( 
.A(n_5842),
.Y(n_6154)
);

INVxp33_ASAP7_75t_L g6155 ( 
.A(n_5861),
.Y(n_6155)
);

AND2x4_ASAP7_75t_L g6156 ( 
.A(n_5800),
.B(n_5449),
.Y(n_6156)
);

INVx1_ASAP7_75t_L g6157 ( 
.A(n_5912),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_5986),
.Y(n_6158)
);

INVx2_ASAP7_75t_L g6159 ( 
.A(n_5802),
.Y(n_6159)
);

INVx2_ASAP7_75t_L g6160 ( 
.A(n_5802),
.Y(n_6160)
);

INVx1_ASAP7_75t_L g6161 ( 
.A(n_5990),
.Y(n_6161)
);

BUFx12f_ASAP7_75t_L g6162 ( 
.A(n_5930),
.Y(n_6162)
);

AOI21x1_ASAP7_75t_L g6163 ( 
.A1(n_5976),
.A2(n_5452),
.B(n_5449),
.Y(n_6163)
);

INVx1_ASAP7_75t_L g6164 ( 
.A(n_5932),
.Y(n_6164)
);

INVx2_ASAP7_75t_L g6165 ( 
.A(n_5802),
.Y(n_6165)
);

BUFx6f_ASAP7_75t_L g6166 ( 
.A(n_5794),
.Y(n_6166)
);

BUFx3_ASAP7_75t_L g6167 ( 
.A(n_5895),
.Y(n_6167)
);

CKINVDCx5p33_ASAP7_75t_R g6168 ( 
.A(n_5955),
.Y(n_6168)
);

HB1xp67_ASAP7_75t_L g6169 ( 
.A(n_5875),
.Y(n_6169)
);

INVx6_ASAP7_75t_L g6170 ( 
.A(n_5794),
.Y(n_6170)
);

AOI22xp5_ASAP7_75t_L g6171 ( 
.A1(n_5893),
.A2(n_5538),
.B1(n_5559),
.B2(n_5458),
.Y(n_6171)
);

HB1xp67_ASAP7_75t_L g6172 ( 
.A(n_5853),
.Y(n_6172)
);

INVx1_ASAP7_75t_SL g6173 ( 
.A(n_5848),
.Y(n_6173)
);

CKINVDCx6p67_ASAP7_75t_R g6174 ( 
.A(n_5979),
.Y(n_6174)
);

AOI22xp5_ASAP7_75t_L g6175 ( 
.A1(n_5832),
.A2(n_5458),
.B1(n_5460),
.B2(n_5452),
.Y(n_6175)
);

INVx1_ASAP7_75t_SL g6176 ( 
.A(n_5848),
.Y(n_6176)
);

INVx2_ASAP7_75t_L g6177 ( 
.A(n_5781),
.Y(n_6177)
);

AO21x1_ASAP7_75t_L g6178 ( 
.A1(n_5973),
.A2(n_5728),
.B(n_84),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_5921),
.Y(n_6179)
);

AND2x2_ASAP7_75t_L g6180 ( 
.A(n_5854),
.B(n_5452),
.Y(n_6180)
);

CKINVDCx6p67_ASAP7_75t_R g6181 ( 
.A(n_5953),
.Y(n_6181)
);

AOI21x1_ASAP7_75t_L g6182 ( 
.A1(n_5991),
.A2(n_5460),
.B(n_5458),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_5934),
.Y(n_6183)
);

INVx2_ASAP7_75t_L g6184 ( 
.A(n_5939),
.Y(n_6184)
);

AOI21x1_ASAP7_75t_L g6185 ( 
.A1(n_5991),
.A2(n_5485),
.B(n_5460),
.Y(n_6185)
);

BUFx6f_ASAP7_75t_L g6186 ( 
.A(n_5794),
.Y(n_6186)
);

OAI21x1_ASAP7_75t_L g6187 ( 
.A1(n_5785),
.A2(n_5750),
.B(n_5758),
.Y(n_6187)
);

OAI21xp5_ASAP7_75t_SL g6188 ( 
.A1(n_5832),
.A2(n_5485),
.B(n_5598),
.Y(n_6188)
);

INVx2_ASAP7_75t_L g6189 ( 
.A(n_5908),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_5944),
.Y(n_6190)
);

INVx3_ASAP7_75t_L g6191 ( 
.A(n_5816),
.Y(n_6191)
);

HB1xp67_ASAP7_75t_L g6192 ( 
.A(n_5795),
.Y(n_6192)
);

INVx2_ASAP7_75t_L g6193 ( 
.A(n_5830),
.Y(n_6193)
);

INVx2_ASAP7_75t_L g6194 ( 
.A(n_5757),
.Y(n_6194)
);

AND2x2_ASAP7_75t_L g6195 ( 
.A(n_5906),
.B(n_5485),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_5956),
.Y(n_6196)
);

INVx1_ASAP7_75t_L g6197 ( 
.A(n_5966),
.Y(n_6197)
);

INVx6_ASAP7_75t_L g6198 ( 
.A(n_5797),
.Y(n_6198)
);

CKINVDCx20_ASAP7_75t_R g6199 ( 
.A(n_5992),
.Y(n_6199)
);

AOI22xp33_ASAP7_75t_SL g6200 ( 
.A1(n_5786),
.A2(n_5624),
.B1(n_5671),
.B2(n_5598),
.Y(n_6200)
);

OAI21x1_ASAP7_75t_L g6201 ( 
.A1(n_5758),
.A2(n_5624),
.B(n_5598),
.Y(n_6201)
);

BUFx6f_ASAP7_75t_SL g6202 ( 
.A(n_5797),
.Y(n_6202)
);

INVx1_ASAP7_75t_L g6203 ( 
.A(n_5967),
.Y(n_6203)
);

INVx1_ASAP7_75t_L g6204 ( 
.A(n_5975),
.Y(n_6204)
);

AOI22xp33_ASAP7_75t_L g6205 ( 
.A1(n_5784),
.A2(n_5821),
.B1(n_5770),
.B2(n_5923),
.Y(n_6205)
);

INVxp33_ASAP7_75t_L g6206 ( 
.A(n_5861),
.Y(n_6206)
);

INVx3_ASAP7_75t_L g6207 ( 
.A(n_5816),
.Y(n_6207)
);

BUFx2_ASAP7_75t_L g6208 ( 
.A(n_5755),
.Y(n_6208)
);

INVx1_ASAP7_75t_SL g6209 ( 
.A(n_5795),
.Y(n_6209)
);

INVx2_ASAP7_75t_L g6210 ( 
.A(n_5996),
.Y(n_6210)
);

HB1xp67_ASAP7_75t_L g6211 ( 
.A(n_5851),
.Y(n_6211)
);

BUFx3_ASAP7_75t_L g6212 ( 
.A(n_5797),
.Y(n_6212)
);

INVx2_ASAP7_75t_L g6213 ( 
.A(n_6006),
.Y(n_6213)
);

NAND2xp5_ASAP7_75t_SL g6214 ( 
.A(n_5845),
.B(n_5624),
.Y(n_6214)
);

OAI21x1_ASAP7_75t_L g6215 ( 
.A1(n_5931),
.A2(n_5704),
.B(n_5671),
.Y(n_6215)
);

INVx2_ASAP7_75t_SL g6216 ( 
.A(n_5950),
.Y(n_6216)
);

OAI21x1_ASAP7_75t_L g6217 ( 
.A1(n_5931),
.A2(n_5704),
.B(n_5671),
.Y(n_6217)
);

OAI22xp33_ASAP7_75t_L g6218 ( 
.A1(n_5784),
.A2(n_5717),
.B1(n_5730),
.B2(n_5704),
.Y(n_6218)
);

AOI22xp33_ASAP7_75t_L g6219 ( 
.A1(n_5821),
.A2(n_5717),
.B1(n_5735),
.B2(n_5730),
.Y(n_6219)
);

AND2x2_ASAP7_75t_L g6220 ( 
.A(n_5882),
.B(n_5717),
.Y(n_6220)
);

AND2x2_ASAP7_75t_L g6221 ( 
.A(n_5924),
.B(n_5811),
.Y(n_6221)
);

NOR2xp33_ASAP7_75t_L g6222 ( 
.A(n_5950),
.B(n_5730),
.Y(n_6222)
);

INVx2_ASAP7_75t_L g6223 ( 
.A(n_6008),
.Y(n_6223)
);

HB1xp67_ASAP7_75t_L g6224 ( 
.A(n_5851),
.Y(n_6224)
);

INVx2_ASAP7_75t_L g6225 ( 
.A(n_5777),
.Y(n_6225)
);

BUFx3_ASAP7_75t_L g6226 ( 
.A(n_5885),
.Y(n_6226)
);

INVx2_ASAP7_75t_L g6227 ( 
.A(n_5777),
.Y(n_6227)
);

INVx1_ASAP7_75t_L g6228 ( 
.A(n_5828),
.Y(n_6228)
);

AOI22xp33_ASAP7_75t_L g6229 ( 
.A1(n_5818),
.A2(n_5735),
.B1(n_2227),
.B2(n_2966),
.Y(n_6229)
);

BUFx2_ASAP7_75t_L g6230 ( 
.A(n_5894),
.Y(n_6230)
);

AND2x2_ASAP7_75t_L g6231 ( 
.A(n_5855),
.B(n_5735),
.Y(n_6231)
);

INVx2_ASAP7_75t_L g6232 ( 
.A(n_5777),
.Y(n_6232)
);

AND2x4_ASAP7_75t_L g6233 ( 
.A(n_5800),
.B(n_86),
.Y(n_6233)
);

OAI22xp33_ASAP7_75t_L g6234 ( 
.A1(n_5894),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_6234)
);

NAND2x1p5_ASAP7_75t_L g6235 ( 
.A(n_5805),
.B(n_3381),
.Y(n_6235)
);

HB1xp67_ASAP7_75t_L g6236 ( 
.A(n_5981),
.Y(n_6236)
);

INVx1_ASAP7_75t_L g6237 ( 
.A(n_5828),
.Y(n_6237)
);

INVx1_ASAP7_75t_L g6238 ( 
.A(n_5865),
.Y(n_6238)
);

OAI22xp33_ASAP7_75t_L g6239 ( 
.A1(n_5894),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_6239)
);

BUFx4_ASAP7_75t_SL g6240 ( 
.A(n_5913),
.Y(n_6240)
);

INVx2_ASAP7_75t_L g6241 ( 
.A(n_5907),
.Y(n_6241)
);

BUFx3_ASAP7_75t_L g6242 ( 
.A(n_5756),
.Y(n_6242)
);

HB1xp67_ASAP7_75t_L g6243 ( 
.A(n_5803),
.Y(n_6243)
);

NAND2x1p5_ASAP7_75t_L g6244 ( 
.A(n_5805),
.B(n_3381),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_5865),
.Y(n_6245)
);

OAI22xp33_ASAP7_75t_L g6246 ( 
.A1(n_5913),
.A2(n_92),
.B1(n_89),
.B2(n_91),
.Y(n_6246)
);

INVx1_ASAP7_75t_L g6247 ( 
.A(n_5883),
.Y(n_6247)
);

INVx2_ASAP7_75t_L g6248 ( 
.A(n_5914),
.Y(n_6248)
);

AOI22xp33_ASAP7_75t_L g6249 ( 
.A1(n_5839),
.A2(n_2227),
.B1(n_2966),
.B2(n_2964),
.Y(n_6249)
);

INVx3_ASAP7_75t_L g6250 ( 
.A(n_5827),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_5883),
.Y(n_6251)
);

AND2x4_ASAP7_75t_L g6252 ( 
.A(n_5749),
.B(n_91),
.Y(n_6252)
);

INVxp67_ASAP7_75t_L g6253 ( 
.A(n_5993),
.Y(n_6253)
);

CKINVDCx11_ASAP7_75t_R g6254 ( 
.A(n_5808),
.Y(n_6254)
);

AOI21x1_ASAP7_75t_L g6255 ( 
.A1(n_6005),
.A2(n_2688),
.B(n_2683),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_5936),
.Y(n_6256)
);

INVx2_ASAP7_75t_SL g6257 ( 
.A(n_5838),
.Y(n_6257)
);

HB1xp67_ASAP7_75t_L g6258 ( 
.A(n_5981),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_5936),
.Y(n_6259)
);

CKINVDCx11_ASAP7_75t_R g6260 ( 
.A(n_5808),
.Y(n_6260)
);

HB1xp67_ASAP7_75t_L g6261 ( 
.A(n_5803),
.Y(n_6261)
);

AND2x2_ASAP7_75t_L g6262 ( 
.A(n_5897),
.B(n_92),
.Y(n_6262)
);

CKINVDCx20_ASAP7_75t_R g6263 ( 
.A(n_5997),
.Y(n_6263)
);

OAI21x1_ASAP7_75t_L g6264 ( 
.A1(n_6001),
.A2(n_2775),
.B(n_2763),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_5874),
.Y(n_6265)
);

BUFx3_ASAP7_75t_L g6266 ( 
.A(n_5852),
.Y(n_6266)
);

INVx4_ASAP7_75t_L g6267 ( 
.A(n_5808),
.Y(n_6267)
);

CKINVDCx6p67_ASAP7_75t_R g6268 ( 
.A(n_5959),
.Y(n_6268)
);

CKINVDCx20_ASAP7_75t_R g6269 ( 
.A(n_5919),
.Y(n_6269)
);

INVx3_ASAP7_75t_L g6270 ( 
.A(n_6123),
.Y(n_6270)
);

NOR2xp33_ASAP7_75t_L g6271 ( 
.A(n_6155),
.B(n_5791),
.Y(n_6271)
);

INVx2_ASAP7_75t_L g6272 ( 
.A(n_6166),
.Y(n_6272)
);

AND2x4_ASAP7_75t_L g6273 ( 
.A(n_6177),
.B(n_5892),
.Y(n_6273)
);

HB1xp67_ASAP7_75t_L g6274 ( 
.A(n_6169),
.Y(n_6274)
);

HB1xp67_ASAP7_75t_L g6275 ( 
.A(n_6169),
.Y(n_6275)
);

INVx2_ASAP7_75t_L g6276 ( 
.A(n_6166),
.Y(n_6276)
);

INVx1_ASAP7_75t_L g6277 ( 
.A(n_6023),
.Y(n_6277)
);

INVx1_ASAP7_75t_L g6278 ( 
.A(n_6024),
.Y(n_6278)
);

INVx1_ASAP7_75t_L g6279 ( 
.A(n_6031),
.Y(n_6279)
);

AND2x2_ASAP7_75t_L g6280 ( 
.A(n_6191),
.B(n_5749),
.Y(n_6280)
);

HB1xp67_ASAP7_75t_SL g6281 ( 
.A(n_6152),
.Y(n_6281)
);

INVx3_ASAP7_75t_L g6282 ( 
.A(n_6123),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_6128),
.Y(n_6283)
);

INVx3_ASAP7_75t_L g6284 ( 
.A(n_6131),
.Y(n_6284)
);

OAI21xp5_ASAP7_75t_L g6285 ( 
.A1(n_6022),
.A2(n_5886),
.B(n_5829),
.Y(n_6285)
);

OAI21x1_ASAP7_75t_L g6286 ( 
.A1(n_6083),
.A2(n_5856),
.B(n_5766),
.Y(n_6286)
);

INVx2_ASAP7_75t_L g6287 ( 
.A(n_6166),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_6137),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_6138),
.Y(n_6289)
);

INVx2_ASAP7_75t_L g6290 ( 
.A(n_6186),
.Y(n_6290)
);

AND2x2_ASAP7_75t_L g6291 ( 
.A(n_6191),
.B(n_5827),
.Y(n_6291)
);

INVx2_ASAP7_75t_L g6292 ( 
.A(n_6186),
.Y(n_6292)
);

OA21x2_ASAP7_75t_L g6293 ( 
.A1(n_6072),
.A2(n_5767),
.B(n_5763),
.Y(n_6293)
);

OAI21xp5_ASAP7_75t_L g6294 ( 
.A1(n_6022),
.A2(n_5886),
.B(n_5829),
.Y(n_6294)
);

INVx1_ASAP7_75t_L g6295 ( 
.A(n_6143),
.Y(n_6295)
);

INVx1_ASAP7_75t_L g6296 ( 
.A(n_6144),
.Y(n_6296)
);

NOR2xp33_ASAP7_75t_L g6297 ( 
.A(n_6206),
.B(n_5772),
.Y(n_6297)
);

OA21x2_ASAP7_75t_L g6298 ( 
.A1(n_6072),
.A2(n_6103),
.B(n_6082),
.Y(n_6298)
);

INVx2_ASAP7_75t_SL g6299 ( 
.A(n_6071),
.Y(n_6299)
);

INVx1_ASAP7_75t_L g6300 ( 
.A(n_6067),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_6068),
.Y(n_6301)
);

A2O1A1Ixp33_ASAP7_75t_L g6302 ( 
.A1(n_6064),
.A2(n_5973),
.B(n_5995),
.C(n_5999),
.Y(n_6302)
);

BUFx3_ASAP7_75t_L g6303 ( 
.A(n_6162),
.Y(n_6303)
);

CKINVDCx10_ASAP7_75t_R g6304 ( 
.A(n_6202),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_6080),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_6093),
.Y(n_6306)
);

INVx2_ASAP7_75t_L g6307 ( 
.A(n_6186),
.Y(n_6307)
);

BUFx3_ASAP7_75t_L g6308 ( 
.A(n_6095),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_6097),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_6099),
.Y(n_6310)
);

NAND2xp5_ASAP7_75t_L g6311 ( 
.A(n_6253),
.B(n_6013),
.Y(n_6311)
);

INVx1_ASAP7_75t_L g6312 ( 
.A(n_6101),
.Y(n_6312)
);

BUFx3_ASAP7_75t_L g6313 ( 
.A(n_6084),
.Y(n_6313)
);

CKINVDCx6p67_ASAP7_75t_R g6314 ( 
.A(n_6028),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_6104),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_6108),
.Y(n_6316)
);

HB1xp67_ASAP7_75t_L g6317 ( 
.A(n_6034),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_6110),
.Y(n_6318)
);

BUFx3_ASAP7_75t_L g6319 ( 
.A(n_6084),
.Y(n_6319)
);

HB1xp67_ASAP7_75t_L g6320 ( 
.A(n_6236),
.Y(n_6320)
);

HB1xp67_ASAP7_75t_L g6321 ( 
.A(n_6236),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_6125),
.Y(n_6322)
);

INVx3_ASAP7_75t_L g6323 ( 
.A(n_6131),
.Y(n_6323)
);

OR2x6_ASAP7_75t_L g6324 ( 
.A(n_6132),
.B(n_5957),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_6126),
.Y(n_6325)
);

INVx1_ASAP7_75t_L g6326 ( 
.A(n_6127),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_6033),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_6037),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_6040),
.Y(n_6329)
);

INVx2_ASAP7_75t_L g6330 ( 
.A(n_6267),
.Y(n_6330)
);

INVx1_ASAP7_75t_SL g6331 ( 
.A(n_6120),
.Y(n_6331)
);

NAND2xp5_ASAP7_75t_L g6332 ( 
.A(n_6253),
.B(n_6005),
.Y(n_6332)
);

HB1xp67_ASAP7_75t_L g6333 ( 
.A(n_6258),
.Y(n_6333)
);

AOI221xp5_ASAP7_75t_L g6334 ( 
.A1(n_6044),
.A2(n_5760),
.B1(n_5999),
.B2(n_5972),
.C(n_5823),
.Y(n_6334)
);

INVx2_ASAP7_75t_L g6335 ( 
.A(n_6267),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_6043),
.Y(n_6336)
);

AOI21x1_ASAP7_75t_L g6337 ( 
.A1(n_6089),
.A2(n_6013),
.B(n_5963),
.Y(n_6337)
);

AO21x2_ASAP7_75t_L g6338 ( 
.A1(n_6192),
.A2(n_5815),
.B(n_5809),
.Y(n_6338)
);

INVx1_ASAP7_75t_L g6339 ( 
.A(n_6060),
.Y(n_6339)
);

OAI222xp33_ASAP7_75t_L g6340 ( 
.A1(n_6087),
.A2(n_6205),
.B1(n_6171),
.B2(n_6175),
.C1(n_6146),
.C2(n_6032),
.Y(n_6340)
);

BUFx3_ASAP7_75t_L g6341 ( 
.A(n_6071),
.Y(n_6341)
);

BUFx2_ASAP7_75t_L g6342 ( 
.A(n_6172),
.Y(n_6342)
);

AO21x1_ASAP7_75t_SL g6343 ( 
.A1(n_6219),
.A2(n_5919),
.B(n_5876),
.Y(n_6343)
);

OAI21x1_ASAP7_75t_L g6344 ( 
.A1(n_6201),
.A2(n_5798),
.B(n_5768),
.Y(n_6344)
);

OR2x6_ASAP7_75t_L g6345 ( 
.A(n_6028),
.B(n_5891),
.Y(n_6345)
);

AOI22xp33_ASAP7_75t_L g6346 ( 
.A1(n_6086),
.A2(n_5792),
.B1(n_5799),
.B2(n_5826),
.Y(n_6346)
);

INVx1_ASAP7_75t_L g6347 ( 
.A(n_6062),
.Y(n_6347)
);

AND2x4_ASAP7_75t_L g6348 ( 
.A(n_6207),
.B(n_5892),
.Y(n_6348)
);

OR2x6_ASAP7_75t_L g6349 ( 
.A(n_6107),
.B(n_5891),
.Y(n_6349)
);

OAI21xp5_ASAP7_75t_L g6350 ( 
.A1(n_6087),
.A2(n_5926),
.B(n_6000),
.Y(n_6350)
);

INVx1_ASAP7_75t_L g6351 ( 
.A(n_6157),
.Y(n_6351)
);

HB1xp67_ASAP7_75t_L g6352 ( 
.A(n_6258),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_6158),
.Y(n_6353)
);

OR2x2_ASAP7_75t_L g6354 ( 
.A(n_6026),
.B(n_5898),
.Y(n_6354)
);

INVx1_ASAP7_75t_L g6355 ( 
.A(n_6161),
.Y(n_6355)
);

OAI222xp33_ASAP7_75t_L g6356 ( 
.A1(n_6171),
.A2(n_6175),
.B1(n_6146),
.B2(n_6032),
.C1(n_6076),
.C2(n_6111),
.Y(n_6356)
);

INVx1_ASAP7_75t_L g6357 ( 
.A(n_6119),
.Y(n_6357)
);

OA21x2_ASAP7_75t_L g6358 ( 
.A1(n_6082),
.A2(n_6001),
.B(n_5748),
.Y(n_6358)
);

INVx2_ASAP7_75t_L g6359 ( 
.A(n_6021),
.Y(n_6359)
);

INVx1_ASAP7_75t_L g6360 ( 
.A(n_6124),
.Y(n_6360)
);

OA21x2_ASAP7_75t_L g6361 ( 
.A1(n_6187),
.A2(n_6019),
.B(n_6016),
.Y(n_6361)
);

HB1xp67_ASAP7_75t_L g6362 ( 
.A(n_6055),
.Y(n_6362)
);

INVx1_ASAP7_75t_L g6363 ( 
.A(n_6079),
.Y(n_6363)
);

OR2x6_ASAP7_75t_L g6364 ( 
.A(n_6107),
.B(n_5916),
.Y(n_6364)
);

INVx1_ASAP7_75t_L g6365 ( 
.A(n_6129),
.Y(n_6365)
);

INVx2_ASAP7_75t_L g6366 ( 
.A(n_6021),
.Y(n_6366)
);

INVx3_ASAP7_75t_L g6367 ( 
.A(n_6113),
.Y(n_6367)
);

OA21x2_ASAP7_75t_L g6368 ( 
.A1(n_6050),
.A2(n_6016),
.B(n_5884),
.Y(n_6368)
);

INVx1_ASAP7_75t_L g6369 ( 
.A(n_6164),
.Y(n_6369)
);

OAI21xp5_ASAP7_75t_L g6370 ( 
.A1(n_6188),
.A2(n_6011),
.B(n_5958),
.Y(n_6370)
);

INVx1_ASAP7_75t_L g6371 ( 
.A(n_6030),
.Y(n_6371)
);

INVx1_ASAP7_75t_L g6372 ( 
.A(n_6048),
.Y(n_6372)
);

HB1xp67_ASAP7_75t_L g6373 ( 
.A(n_6055),
.Y(n_6373)
);

HB1xp67_ASAP7_75t_L g6374 ( 
.A(n_6055),
.Y(n_6374)
);

CKINVDCx20_ASAP7_75t_R g6375 ( 
.A(n_6052),
.Y(n_6375)
);

INVx1_ASAP7_75t_L g6376 ( 
.A(n_6049),
.Y(n_6376)
);

INVx2_ASAP7_75t_SL g6377 ( 
.A(n_6098),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_6057),
.Y(n_6378)
);

INVx2_ASAP7_75t_L g6379 ( 
.A(n_6105),
.Y(n_6379)
);

HB1xp67_ASAP7_75t_L g6380 ( 
.A(n_6243),
.Y(n_6380)
);

HB1xp67_ASAP7_75t_L g6381 ( 
.A(n_6261),
.Y(n_6381)
);

INVx3_ASAP7_75t_L g6382 ( 
.A(n_6113),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_6228),
.Y(n_6383)
);

NOR2xp33_ASAP7_75t_L g6384 ( 
.A(n_6174),
.B(n_6152),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_6237),
.Y(n_6385)
);

OR2x2_ASAP7_75t_L g6386 ( 
.A(n_6039),
.B(n_5905),
.Y(n_6386)
);

INVx2_ASAP7_75t_L g6387 ( 
.A(n_6105),
.Y(n_6387)
);

AND2x2_ASAP7_75t_L g6388 ( 
.A(n_6250),
.B(n_5881),
.Y(n_6388)
);

OR2x6_ASAP7_75t_L g6389 ( 
.A(n_6069),
.B(n_6188),
.Y(n_6389)
);

OAI21x1_ASAP7_75t_L g6390 ( 
.A1(n_6235),
.A2(n_6244),
.B(n_6250),
.Y(n_6390)
);

INVx1_ASAP7_75t_SL g6391 ( 
.A(n_6120),
.Y(n_6391)
);

INVx2_ASAP7_75t_L g6392 ( 
.A(n_6230),
.Y(n_6392)
);

INVx2_ASAP7_75t_L g6393 ( 
.A(n_6163),
.Y(n_6393)
);

INVx2_ASAP7_75t_L g6394 ( 
.A(n_6182),
.Y(n_6394)
);

INVx3_ASAP7_75t_L g6395 ( 
.A(n_6106),
.Y(n_6395)
);

INVx2_ASAP7_75t_L g6396 ( 
.A(n_6185),
.Y(n_6396)
);

INVx1_ASAP7_75t_L g6397 ( 
.A(n_6238),
.Y(n_6397)
);

INVx1_ASAP7_75t_L g6398 ( 
.A(n_6245),
.Y(n_6398)
);

INVx2_ASAP7_75t_SL g6399 ( 
.A(n_6098),
.Y(n_6399)
);

INVx2_ASAP7_75t_SL g6400 ( 
.A(n_6038),
.Y(n_6400)
);

BUFx3_ASAP7_75t_L g6401 ( 
.A(n_6042),
.Y(n_6401)
);

INVx1_ASAP7_75t_L g6402 ( 
.A(n_6247),
.Y(n_6402)
);

INVx2_ASAP7_75t_L g6403 ( 
.A(n_6096),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_6251),
.Y(n_6404)
);

AOI22xp33_ASAP7_75t_L g6405 ( 
.A1(n_6075),
.A2(n_5792),
.B1(n_5799),
.B2(n_5958),
.Y(n_6405)
);

NAND2xp5_ASAP7_75t_L g6406 ( 
.A(n_6256),
.B(n_5977),
.Y(n_6406)
);

AND2x2_ASAP7_75t_L g6407 ( 
.A(n_6208),
.B(n_5881),
.Y(n_6407)
);

NAND2xp5_ASAP7_75t_L g6408 ( 
.A(n_6259),
.B(n_5977),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_6179),
.Y(n_6409)
);

BUFx2_ASAP7_75t_L g6410 ( 
.A(n_6145),
.Y(n_6410)
);

INVx2_ASAP7_75t_SL g6411 ( 
.A(n_6038),
.Y(n_6411)
);

INVx1_ASAP7_75t_L g6412 ( 
.A(n_6183),
.Y(n_6412)
);

HB1xp67_ASAP7_75t_L g6413 ( 
.A(n_6112),
.Y(n_6413)
);

INVxp67_ASAP7_75t_L g6414 ( 
.A(n_6145),
.Y(n_6414)
);

INVx2_ASAP7_75t_L g6415 ( 
.A(n_6096),
.Y(n_6415)
);

INVx2_ASAP7_75t_L g6416 ( 
.A(n_6115),
.Y(n_6416)
);

INVx1_ASAP7_75t_L g6417 ( 
.A(n_6140),
.Y(n_6417)
);

INVx1_ASAP7_75t_L g6418 ( 
.A(n_6061),
.Y(n_6418)
);

INVx1_ASAP7_75t_L g6419 ( 
.A(n_6073),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_6077),
.Y(n_6420)
);

BUFx2_ASAP7_75t_L g6421 ( 
.A(n_6173),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_6090),
.Y(n_6422)
);

NAND2xp5_ASAP7_75t_L g6423 ( 
.A(n_6041),
.B(n_6002),
.Y(n_6423)
);

BUFx2_ASAP7_75t_L g6424 ( 
.A(n_6173),
.Y(n_6424)
);

INVx1_ASAP7_75t_L g6425 ( 
.A(n_6091),
.Y(n_6425)
);

INVx2_ASAP7_75t_SL g6426 ( 
.A(n_6170),
.Y(n_6426)
);

INVx4_ASAP7_75t_L g6427 ( 
.A(n_6085),
.Y(n_6427)
);

AOI21x1_ASAP7_75t_L g6428 ( 
.A1(n_6214),
.A2(n_5965),
.B(n_5910),
.Y(n_6428)
);

BUFx3_ASAP7_75t_L g6429 ( 
.A(n_6150),
.Y(n_6429)
);

AND2x2_ASAP7_75t_L g6430 ( 
.A(n_6058),
.B(n_5915),
.Y(n_6430)
);

NAND2xp5_ASAP7_75t_L g6431 ( 
.A(n_6041),
.B(n_6209),
.Y(n_6431)
);

INVx5_ASAP7_75t_SL g6432 ( 
.A(n_6233),
.Y(n_6432)
);

INVx1_ASAP7_75t_L g6433 ( 
.A(n_6100),
.Y(n_6433)
);

OAI21x1_ASAP7_75t_L g6434 ( 
.A1(n_6059),
.A2(n_5833),
.B(n_5961),
.Y(n_6434)
);

HB1xp67_ASAP7_75t_L g6435 ( 
.A(n_6112),
.Y(n_6435)
);

INVx3_ASAP7_75t_L g6436 ( 
.A(n_6115),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_6190),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_6196),
.Y(n_6438)
);

AOI22xp33_ASAP7_75t_L g6439 ( 
.A1(n_6066),
.A2(n_5970),
.B1(n_5933),
.B2(n_5863),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_6081),
.Y(n_6440)
);

CKINVDCx11_ASAP7_75t_R g6441 ( 
.A(n_6199),
.Y(n_6441)
);

INVx2_ASAP7_75t_L g6442 ( 
.A(n_6170),
.Y(n_6442)
);

OR2x6_ASAP7_75t_L g6443 ( 
.A(n_6069),
.B(n_6053),
.Y(n_6443)
);

NAND2x1p5_ASAP7_75t_L g6444 ( 
.A(n_6176),
.B(n_5806),
.Y(n_6444)
);

INVx2_ASAP7_75t_L g6445 ( 
.A(n_6198),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_6197),
.Y(n_6446)
);

INVx1_ASAP7_75t_L g6447 ( 
.A(n_6203),
.Y(n_6447)
);

INVx2_ASAP7_75t_SL g6448 ( 
.A(n_6198),
.Y(n_6448)
);

AND2x2_ASAP7_75t_L g6449 ( 
.A(n_6058),
.B(n_5915),
.Y(n_6449)
);

OAI22xp5_ASAP7_75t_L g6450 ( 
.A1(n_6076),
.A2(n_5970),
.B1(n_5933),
.B2(n_5913),
.Y(n_6450)
);

OAI22xp5_ASAP7_75t_L g6451 ( 
.A1(n_6142),
.A2(n_5869),
.B1(n_5871),
.B2(n_5925),
.Y(n_6451)
);

OAI21xp5_ASAP7_75t_L g6452 ( 
.A1(n_6111),
.A2(n_5814),
.B(n_5844),
.Y(n_6452)
);

HB1xp67_ASAP7_75t_L g6453 ( 
.A(n_6029),
.Y(n_6453)
);

AO21x2_ASAP7_75t_L g6454 ( 
.A1(n_6211),
.A2(n_5964),
.B(n_5812),
.Y(n_6454)
);

INVx1_ASAP7_75t_L g6455 ( 
.A(n_6204),
.Y(n_6455)
);

NAND2xp5_ASAP7_75t_L g6456 ( 
.A(n_6041),
.B(n_6002),
.Y(n_6456)
);

AND2x2_ASAP7_75t_L g6457 ( 
.A(n_6121),
.B(n_5871),
.Y(n_6457)
);

AOI21x1_ASAP7_75t_L g6458 ( 
.A1(n_6262),
.A2(n_6017),
.B(n_5871),
.Y(n_6458)
);

HB1xp67_ASAP7_75t_L g6459 ( 
.A(n_6074),
.Y(n_6459)
);

INVx2_ASAP7_75t_L g6460 ( 
.A(n_6159),
.Y(n_6460)
);

AND2x2_ASAP7_75t_L g6461 ( 
.A(n_6121),
.B(n_6156),
.Y(n_6461)
);

INVx2_ASAP7_75t_L g6462 ( 
.A(n_6160),
.Y(n_6462)
);

HB1xp67_ASAP7_75t_L g6463 ( 
.A(n_6074),
.Y(n_6463)
);

INVx2_ASAP7_75t_L g6464 ( 
.A(n_6165),
.Y(n_6464)
);

OAI21x1_ASAP7_75t_L g6465 ( 
.A1(n_6027),
.A2(n_5988),
.B(n_5989),
.Y(n_6465)
);

NAND2xp5_ASAP7_75t_L g6466 ( 
.A(n_6209),
.B(n_6002),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_6065),
.Y(n_6467)
);

INVx1_ASAP7_75t_L g6468 ( 
.A(n_6184),
.Y(n_6468)
);

HB1xp67_ASAP7_75t_L g6469 ( 
.A(n_6224),
.Y(n_6469)
);

AOI21x1_ASAP7_75t_L g6470 ( 
.A1(n_6114),
.A2(n_6017),
.B(n_5998),
.Y(n_6470)
);

INVx2_ASAP7_75t_L g6471 ( 
.A(n_6225),
.Y(n_6471)
);

INVx1_ASAP7_75t_L g6472 ( 
.A(n_6176),
.Y(n_6472)
);

INVx3_ASAP7_75t_L g6473 ( 
.A(n_6156),
.Y(n_6473)
);

HB1xp67_ASAP7_75t_L g6474 ( 
.A(n_6092),
.Y(n_6474)
);

NAND2xp5_ASAP7_75t_L g6475 ( 
.A(n_6265),
.B(n_5764),
.Y(n_6475)
);

INVx1_ASAP7_75t_L g6476 ( 
.A(n_6210),
.Y(n_6476)
);

INVx2_ASAP7_75t_L g6477 ( 
.A(n_6227),
.Y(n_6477)
);

INVx1_ASAP7_75t_L g6478 ( 
.A(n_6213),
.Y(n_6478)
);

INVx1_ASAP7_75t_SL g6479 ( 
.A(n_6240),
.Y(n_6479)
);

INVx2_ASAP7_75t_L g6480 ( 
.A(n_6232),
.Y(n_6480)
);

INVx2_ASAP7_75t_L g6481 ( 
.A(n_6102),
.Y(n_6481)
);

NAND2xp5_ASAP7_75t_L g6482 ( 
.A(n_6200),
.B(n_5764),
.Y(n_6482)
);

CKINVDCx14_ASAP7_75t_R g6483 ( 
.A(n_6263),
.Y(n_6483)
);

INVx1_ASAP7_75t_L g6484 ( 
.A(n_6223),
.Y(n_6484)
);

INVx2_ASAP7_75t_L g6485 ( 
.A(n_6116),
.Y(n_6485)
);

OAI21x1_ASAP7_75t_L g6486 ( 
.A1(n_6109),
.A2(n_5988),
.B(n_5989),
.Y(n_6486)
);

BUFx6f_ASAP7_75t_L g6487 ( 
.A(n_6254),
.Y(n_6487)
);

INVx1_ASAP7_75t_L g6488 ( 
.A(n_6092),
.Y(n_6488)
);

INVx2_ASAP7_75t_L g6489 ( 
.A(n_6117),
.Y(n_6489)
);

BUFx2_ASAP7_75t_L g6490 ( 
.A(n_6135),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_6241),
.Y(n_6491)
);

INVx1_ASAP7_75t_L g6492 ( 
.A(n_6248),
.Y(n_6492)
);

INVx2_ASAP7_75t_L g6493 ( 
.A(n_6133),
.Y(n_6493)
);

OAI21x1_ASAP7_75t_L g6494 ( 
.A1(n_6215),
.A2(n_6014),
.B(n_6003),
.Y(n_6494)
);

CKINVDCx6p67_ASAP7_75t_R g6495 ( 
.A(n_6025),
.Y(n_6495)
);

AOI21x1_ASAP7_75t_L g6496 ( 
.A1(n_6063),
.A2(n_6216),
.B(n_6139),
.Y(n_6496)
);

INVx1_ASAP7_75t_L g6497 ( 
.A(n_6189),
.Y(n_6497)
);

AOI21x1_ASAP7_75t_L g6498 ( 
.A1(n_6051),
.A2(n_6017),
.B(n_5987),
.Y(n_6498)
);

INVx1_ASAP7_75t_L g6499 ( 
.A(n_6193),
.Y(n_6499)
);

INVx1_ASAP7_75t_L g6500 ( 
.A(n_6194),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_6257),
.Y(n_6501)
);

INVx2_ASAP7_75t_L g6502 ( 
.A(n_6147),
.Y(n_6502)
);

AOI33xp33_ASAP7_75t_L g6503 ( 
.A1(n_6334),
.A2(n_6118),
.A3(n_6200),
.B1(n_6036),
.B2(n_6136),
.B3(n_6234),
.Y(n_6503)
);

INVx3_ASAP7_75t_L g6504 ( 
.A(n_6487),
.Y(n_6504)
);

AO21x2_ASAP7_75t_L g6505 ( 
.A1(n_6320),
.A2(n_6094),
.B(n_6239),
.Y(n_6505)
);

OAI21x1_ASAP7_75t_L g6506 ( 
.A1(n_6496),
.A2(n_6217),
.B(n_6151),
.Y(n_6506)
);

AOI22xp5_ASAP7_75t_L g6507 ( 
.A1(n_6334),
.A2(n_6118),
.B1(n_6141),
.B2(n_6269),
.Y(n_6507)
);

AO22x1_ASAP7_75t_L g6508 ( 
.A1(n_6285),
.A2(n_6141),
.B1(n_6252),
.B2(n_6233),
.Y(n_6508)
);

AND2x2_ASAP7_75t_L g6509 ( 
.A(n_6461),
.B(n_6148),
.Y(n_6509)
);

NOR2xp33_ASAP7_75t_L g6510 ( 
.A(n_6479),
.B(n_6056),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_6274),
.Y(n_6511)
);

AND2x4_ASAP7_75t_L g6512 ( 
.A(n_6367),
.B(n_6266),
.Y(n_6512)
);

AOI22xp33_ASAP7_75t_L g6513 ( 
.A1(n_6285),
.A2(n_6069),
.B1(n_6218),
.B2(n_6130),
.Y(n_6513)
);

INVx1_ASAP7_75t_L g6514 ( 
.A(n_6274),
.Y(n_6514)
);

A2O1A1Ixp33_ASAP7_75t_L g6515 ( 
.A1(n_6294),
.A2(n_6136),
.B(n_6046),
.C(n_6134),
.Y(n_6515)
);

AOI22xp33_ASAP7_75t_L g6516 ( 
.A1(n_6294),
.A2(n_6178),
.B1(n_6054),
.B2(n_6035),
.Y(n_6516)
);

AO31x2_ASAP7_75t_L g6517 ( 
.A1(n_6423),
.A2(n_6222),
.A3(n_6149),
.B(n_6154),
.Y(n_6517)
);

AOI22xp5_ASAP7_75t_L g6518 ( 
.A1(n_6271),
.A2(n_6246),
.B1(n_6202),
.B2(n_6070),
.Y(n_6518)
);

OAI22xp5_ASAP7_75t_L g6519 ( 
.A1(n_6302),
.A2(n_6181),
.B1(n_6268),
.B2(n_6249),
.Y(n_6519)
);

INVx2_ASAP7_75t_SL g6520 ( 
.A(n_6304),
.Y(n_6520)
);

HB1xp67_ASAP7_75t_SL g6521 ( 
.A(n_6281),
.Y(n_6521)
);

INVx1_ASAP7_75t_L g6522 ( 
.A(n_6275),
.Y(n_6522)
);

INVx1_ASAP7_75t_L g6523 ( 
.A(n_6275),
.Y(n_6523)
);

NOR2xp33_ASAP7_75t_L g6524 ( 
.A(n_6479),
.B(n_6088),
.Y(n_6524)
);

AOI22xp33_ASAP7_75t_L g6525 ( 
.A1(n_6350),
.A2(n_6070),
.B1(n_6229),
.B2(n_6045),
.Y(n_6525)
);

AO221x2_ASAP7_75t_L g6526 ( 
.A1(n_6340),
.A2(n_6045),
.B1(n_6153),
.B2(n_6260),
.C(n_6252),
.Y(n_6526)
);

INVx4_ASAP7_75t_SL g6527 ( 
.A(n_6313),
.Y(n_6527)
);

OAI22xp5_ASAP7_75t_L g6528 ( 
.A1(n_6302),
.A2(n_6226),
.B1(n_6242),
.B2(n_6212),
.Y(n_6528)
);

AOI22xp33_ASAP7_75t_L g6529 ( 
.A1(n_6350),
.A2(n_6452),
.B1(n_6271),
.B2(n_6450),
.Y(n_6529)
);

OAI22xp5_ASAP7_75t_L g6530 ( 
.A1(n_6439),
.A2(n_6231),
.B1(n_6167),
.B2(n_6180),
.Y(n_6530)
);

OAI22xp5_ASAP7_75t_L g6531 ( 
.A1(n_6439),
.A2(n_6221),
.B1(n_6122),
.B2(n_6195),
.Y(n_6531)
);

INVx5_ASAP7_75t_L g6532 ( 
.A(n_6487),
.Y(n_6532)
);

OR2x6_ASAP7_75t_L g6533 ( 
.A(n_6377),
.B(n_5819),
.Y(n_6533)
);

INVx1_ASAP7_75t_L g6534 ( 
.A(n_6320),
.Y(n_6534)
);

AOI221xp5_ASAP7_75t_L g6535 ( 
.A1(n_6340),
.A2(n_6356),
.B1(n_6346),
.B2(n_6332),
.C(n_6311),
.Y(n_6535)
);

INVx2_ASAP7_75t_L g6536 ( 
.A(n_6367),
.Y(n_6536)
);

INVx1_ASAP7_75t_L g6537 ( 
.A(n_6321),
.Y(n_6537)
);

AOI21xp33_ASAP7_75t_SL g6538 ( 
.A1(n_6384),
.A2(n_6168),
.B(n_6078),
.Y(n_6538)
);

OAI22xp5_ASAP7_75t_L g6539 ( 
.A1(n_6450),
.A2(n_6255),
.B1(n_6220),
.B2(n_5969),
.Y(n_6539)
);

AOI221xp5_ASAP7_75t_L g6540 ( 
.A1(n_6356),
.A2(n_6012),
.B1(n_5969),
.B2(n_5819),
.C(n_5952),
.Y(n_6540)
);

NAND2xp5_ASAP7_75t_SL g6541 ( 
.A(n_6452),
.B(n_6047),
.Y(n_6541)
);

OAI22xp5_ASAP7_75t_L g6542 ( 
.A1(n_6389),
.A2(n_5969),
.B1(n_5819),
.B2(n_6007),
.Y(n_6542)
);

AOI22xp33_ASAP7_75t_SL g6543 ( 
.A1(n_6483),
.A2(n_5941),
.B1(n_6047),
.B2(n_6264),
.Y(n_6543)
);

OAI221xp5_ASAP7_75t_L g6544 ( 
.A1(n_6346),
.A2(n_6405),
.B1(n_6370),
.B2(n_6389),
.C(n_6443),
.Y(n_6544)
);

OAI22xp33_ASAP7_75t_L g6545 ( 
.A1(n_6389),
.A2(n_6014),
.B1(n_6003),
.B2(n_5941),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_6331),
.B(n_6047),
.Y(n_6546)
);

AOI22xp33_ASAP7_75t_L g6547 ( 
.A1(n_6467),
.A2(n_6392),
.B1(n_6382),
.B2(n_6297),
.Y(n_6547)
);

OAI22xp5_ASAP7_75t_L g6548 ( 
.A1(n_6405),
.A2(n_5941),
.B1(n_6047),
.B2(n_5937),
.Y(n_6548)
);

NAND3xp33_ASAP7_75t_L g6549 ( 
.A(n_6466),
.B(n_6047),
.C(n_93),
.Y(n_6549)
);

OAI22xp5_ASAP7_75t_L g6550 ( 
.A1(n_6414),
.A2(n_5948),
.B1(n_5962),
.B2(n_5984),
.Y(n_6550)
);

AO22x1_ASAP7_75t_L g6551 ( 
.A1(n_6370),
.A2(n_5948),
.B1(n_5928),
.B2(n_5962),
.Y(n_6551)
);

INVx1_ASAP7_75t_L g6552 ( 
.A(n_6321),
.Y(n_6552)
);

NAND3xp33_ASAP7_75t_L g6553 ( 
.A(n_6466),
.B(n_94),
.C(n_95),
.Y(n_6553)
);

OR2x2_ASAP7_75t_L g6554 ( 
.A(n_6342),
.B(n_5943),
.Y(n_6554)
);

OAI22xp5_ASAP7_75t_L g6555 ( 
.A1(n_6414),
.A2(n_5983),
.B1(n_5974),
.B2(n_5949),
.Y(n_6555)
);

AOI21xp33_ASAP7_75t_L g6556 ( 
.A1(n_6423),
.A2(n_5911),
.B(n_94),
.Y(n_6556)
);

AOI22xp33_ASAP7_75t_L g6557 ( 
.A1(n_6297),
.A2(n_5899),
.B1(n_2227),
.B2(n_2688),
.Y(n_6557)
);

OAI21x1_ASAP7_75t_L g6558 ( 
.A1(n_6444),
.A2(n_95),
.B(n_97),
.Y(n_6558)
);

AND2x2_ASAP7_75t_L g6559 ( 
.A(n_6430),
.B(n_97),
.Y(n_6559)
);

INVx1_ASAP7_75t_L g6560 ( 
.A(n_6333),
.Y(n_6560)
);

OAI21xp33_ASAP7_75t_SL g6561 ( 
.A1(n_6434),
.A2(n_98),
.B(n_99),
.Y(n_6561)
);

AND2x4_ASAP7_75t_L g6562 ( 
.A(n_6270),
.B(n_99),
.Y(n_6562)
);

AOI22xp33_ASAP7_75t_L g6563 ( 
.A1(n_6343),
.A2(n_2967),
.B1(n_2970),
.B2(n_2966),
.Y(n_6563)
);

AOI22xp5_ASAP7_75t_L g6564 ( 
.A1(n_6443),
.A2(n_6399),
.B1(n_6472),
.B2(n_6349),
.Y(n_6564)
);

OAI22xp33_ASAP7_75t_L g6565 ( 
.A1(n_6443),
.A2(n_6421),
.B1(n_6424),
.B2(n_6410),
.Y(n_6565)
);

INVx1_ASAP7_75t_L g6566 ( 
.A(n_6333),
.Y(n_6566)
);

BUFx3_ASAP7_75t_L g6567 ( 
.A(n_6429),
.Y(n_6567)
);

NAND2xp5_ASAP7_75t_L g6568 ( 
.A(n_6331),
.B(n_6391),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_6352),
.Y(n_6569)
);

AO222x2_ASAP7_75t_L g6570 ( 
.A1(n_6281),
.A2(n_104),
.B1(n_106),
.B2(n_101),
.C1(n_102),
.C2(n_105),
.Y(n_6570)
);

AOI22xp33_ASAP7_75t_L g6571 ( 
.A1(n_6499),
.A2(n_2967),
.B1(n_2970),
.B2(n_2966),
.Y(n_6571)
);

AOI221xp5_ASAP7_75t_L g6572 ( 
.A1(n_6311),
.A2(n_105),
.B1(n_101),
.B2(n_102),
.C(n_106),
.Y(n_6572)
);

NOR2xp67_ASAP7_75t_L g6573 ( 
.A(n_6395),
.B(n_108),
.Y(n_6573)
);

OAI211xp5_ASAP7_75t_L g6574 ( 
.A1(n_6482),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_6574)
);

INVx2_ASAP7_75t_L g6575 ( 
.A(n_6436),
.Y(n_6575)
);

AOI22xp33_ASAP7_75t_SL g6576 ( 
.A1(n_6432),
.A2(n_114),
.B1(n_110),
.B2(n_113),
.Y(n_6576)
);

OAI21x1_ASAP7_75t_L g6577 ( 
.A1(n_6444),
.A2(n_114),
.B(n_115),
.Y(n_6577)
);

AOI22xp33_ASAP7_75t_L g6578 ( 
.A1(n_6491),
.A2(n_2970),
.B1(n_2967),
.B2(n_3421),
.Y(n_6578)
);

INVx2_ASAP7_75t_L g6579 ( 
.A(n_6436),
.Y(n_6579)
);

AND2x2_ASAP7_75t_L g6580 ( 
.A(n_6449),
.B(n_116),
.Y(n_6580)
);

OAI21x1_ASAP7_75t_L g6581 ( 
.A1(n_6390),
.A2(n_116),
.B(n_117),
.Y(n_6581)
);

OAI22xp5_ASAP7_75t_SL g6582 ( 
.A1(n_6324),
.A2(n_120),
.B1(n_117),
.B2(n_118),
.Y(n_6582)
);

INVx2_ASAP7_75t_L g6583 ( 
.A(n_6270),
.Y(n_6583)
);

A2O1A1Ixp33_ASAP7_75t_L g6584 ( 
.A1(n_6456),
.A2(n_6391),
.B(n_6482),
.C(n_6411),
.Y(n_6584)
);

AND2x4_ASAP7_75t_L g6585 ( 
.A(n_6282),
.B(n_118),
.Y(n_6585)
);

INVx4_ASAP7_75t_L g6586 ( 
.A(n_6319),
.Y(n_6586)
);

OAI221xp5_ASAP7_75t_L g6587 ( 
.A1(n_6345),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.C(n_123),
.Y(n_6587)
);

AOI22xp33_ASAP7_75t_L g6588 ( 
.A1(n_6492),
.A2(n_2970),
.B1(n_2967),
.B2(n_3421),
.Y(n_6588)
);

OAI22xp5_ASAP7_75t_L g6589 ( 
.A1(n_6324),
.A2(n_126),
.B1(n_121),
.B2(n_125),
.Y(n_6589)
);

OR2x6_ASAP7_75t_L g6590 ( 
.A(n_6345),
.B(n_127),
.Y(n_6590)
);

AOI221xp5_ASAP7_75t_L g6591 ( 
.A1(n_6332),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.C(n_131),
.Y(n_6591)
);

NOR2xp33_ASAP7_75t_L g6592 ( 
.A(n_6400),
.B(n_129),
.Y(n_6592)
);

OAI211xp5_ASAP7_75t_L g6593 ( 
.A1(n_6362),
.A2(n_134),
.B(n_132),
.C(n_133),
.Y(n_6593)
);

OR2x2_ASAP7_75t_L g6594 ( 
.A(n_6363),
.B(n_136),
.Y(n_6594)
);

AOI221xp5_ASAP7_75t_L g6595 ( 
.A1(n_6417),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.C(n_139),
.Y(n_6595)
);

AOI221xp5_ASAP7_75t_L g6596 ( 
.A1(n_6431),
.A2(n_142),
.B1(n_139),
.B2(n_141),
.C(n_143),
.Y(n_6596)
);

AOI222xp33_ASAP7_75t_L g6597 ( 
.A1(n_6365),
.A2(n_145),
.B1(n_147),
.B2(n_141),
.C1(n_144),
.C2(n_146),
.Y(n_6597)
);

HB1xp67_ASAP7_75t_L g6598 ( 
.A(n_6380),
.Y(n_6598)
);

AOI222xp33_ASAP7_75t_L g6599 ( 
.A1(n_6406),
.A2(n_149),
.B1(n_151),
.B2(n_144),
.C1(n_148),
.C2(n_150),
.Y(n_6599)
);

BUFx2_ASAP7_75t_L g6600 ( 
.A(n_6324),
.Y(n_6600)
);

AOI21xp5_ASAP7_75t_L g6601 ( 
.A1(n_6406),
.A2(n_150),
.B(n_152),
.Y(n_6601)
);

OAI221xp5_ASAP7_75t_L g6602 ( 
.A1(n_6345),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.C(n_155),
.Y(n_6602)
);

AOI222xp33_ASAP7_75t_L g6603 ( 
.A1(n_6408),
.A2(n_6369),
.B1(n_6451),
.B2(n_6381),
.C1(n_6380),
.C2(n_6431),
.Y(n_6603)
);

AO21x2_ASAP7_75t_L g6604 ( 
.A1(n_6352),
.A2(n_154),
.B(n_156),
.Y(n_6604)
);

AOI22xp33_ASAP7_75t_L g6605 ( 
.A1(n_6440),
.A2(n_2970),
.B1(n_2967),
.B2(n_3421),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_6277),
.Y(n_6606)
);

AOI22xp33_ASAP7_75t_SL g6607 ( 
.A1(n_6432),
.A2(n_6451),
.B1(n_6362),
.B2(n_6374),
.Y(n_6607)
);

OAI211xp5_ASAP7_75t_L g6608 ( 
.A1(n_6373),
.A2(n_158),
.B(n_156),
.C(n_157),
.Y(n_6608)
);

AND2x2_ASAP7_75t_L g6609 ( 
.A(n_6291),
.B(n_157),
.Y(n_6609)
);

AND2x4_ASAP7_75t_L g6610 ( 
.A(n_6282),
.B(n_159),
.Y(n_6610)
);

OAI22xp5_ASAP7_75t_L g6611 ( 
.A1(n_6426),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_6611)
);

AND2x2_ASAP7_75t_L g6612 ( 
.A(n_6388),
.B(n_163),
.Y(n_6612)
);

OR2x6_ASAP7_75t_L g6613 ( 
.A(n_6349),
.B(n_164),
.Y(n_6613)
);

OAI22xp33_ASAP7_75t_L g6614 ( 
.A1(n_6473),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_6278),
.Y(n_6615)
);

HB1xp67_ASAP7_75t_L g6616 ( 
.A(n_6381),
.Y(n_6616)
);

INVx2_ASAP7_75t_L g6617 ( 
.A(n_6284),
.Y(n_6617)
);

OAI22xp33_ASAP7_75t_L g6618 ( 
.A1(n_6473),
.A2(n_169),
.B1(n_165),
.B2(n_168),
.Y(n_6618)
);

HB1xp67_ASAP7_75t_L g6619 ( 
.A(n_6317),
.Y(n_6619)
);

AOI22xp33_ASAP7_75t_SL g6620 ( 
.A1(n_6432),
.A2(n_172),
.B1(n_169),
.B2(n_170),
.Y(n_6620)
);

AOI22xp33_ASAP7_75t_L g6621 ( 
.A1(n_6349),
.A2(n_3421),
.B1(n_3290),
.B2(n_3286),
.Y(n_6621)
);

INVx4_ASAP7_75t_SL g6622 ( 
.A(n_6341),
.Y(n_6622)
);

AND2x2_ASAP7_75t_L g6623 ( 
.A(n_6407),
.B(n_172),
.Y(n_6623)
);

INVx2_ASAP7_75t_L g6624 ( 
.A(n_6284),
.Y(n_6624)
);

INVx1_ASAP7_75t_L g6625 ( 
.A(n_6279),
.Y(n_6625)
);

AND2x2_ASAP7_75t_L g6626 ( 
.A(n_6280),
.B(n_173),
.Y(n_6626)
);

AOI22xp33_ASAP7_75t_L g6627 ( 
.A1(n_6457),
.A2(n_3290),
.B1(n_3286),
.B2(n_1325),
.Y(n_6627)
);

AND2x2_ASAP7_75t_L g6628 ( 
.A(n_6442),
.B(n_174),
.Y(n_6628)
);

OAI211xp5_ASAP7_75t_L g6629 ( 
.A1(n_6373),
.A2(n_181),
.B(n_175),
.C(n_178),
.Y(n_6629)
);

INVx2_ASAP7_75t_L g6630 ( 
.A(n_6323),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_6445),
.B(n_175),
.Y(n_6631)
);

INVx2_ASAP7_75t_L g6632 ( 
.A(n_6323),
.Y(n_6632)
);

CKINVDCx5p33_ASAP7_75t_R g6633 ( 
.A(n_6441),
.Y(n_6633)
);

INVx2_ASAP7_75t_L g6634 ( 
.A(n_6308),
.Y(n_6634)
);

INVx1_ASAP7_75t_L g6635 ( 
.A(n_6327),
.Y(n_6635)
);

INVx2_ASAP7_75t_L g6636 ( 
.A(n_6490),
.Y(n_6636)
);

AOI22xp33_ASAP7_75t_L g6637 ( 
.A1(n_6314),
.A2(n_3290),
.B1(n_1325),
.B2(n_1337),
.Y(n_6637)
);

INVx4_ASAP7_75t_L g6638 ( 
.A(n_6495),
.Y(n_6638)
);

INVx2_ASAP7_75t_L g6639 ( 
.A(n_6272),
.Y(n_6639)
);

BUFx3_ASAP7_75t_L g6640 ( 
.A(n_6303),
.Y(n_6640)
);

NAND2xp5_ASAP7_75t_L g6641 ( 
.A(n_6276),
.B(n_181),
.Y(n_6641)
);

INVx2_ASAP7_75t_L g6642 ( 
.A(n_6287),
.Y(n_6642)
);

AO21x2_ASAP7_75t_L g6643 ( 
.A1(n_6317),
.A2(n_182),
.B(n_184),
.Y(n_6643)
);

OAI22xp5_ASAP7_75t_L g6644 ( 
.A1(n_6448),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_6644)
);

OAI22xp33_ASAP7_75t_L g6645 ( 
.A1(n_6364),
.A2(n_188),
.B1(n_185),
.B2(n_187),
.Y(n_6645)
);

NAND2xp5_ASAP7_75t_L g6646 ( 
.A(n_6290),
.B(n_188),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6328),
.Y(n_6647)
);

AOI22xp33_ASAP7_75t_L g6648 ( 
.A1(n_6330),
.A2(n_1325),
.B1(n_1337),
.B2(n_1250),
.Y(n_6648)
);

INVx2_ASAP7_75t_L g6649 ( 
.A(n_6292),
.Y(n_6649)
);

INVx2_ASAP7_75t_L g6650 ( 
.A(n_6307),
.Y(n_6650)
);

INVx2_ASAP7_75t_L g6651 ( 
.A(n_6335),
.Y(n_6651)
);

INVx3_ASAP7_75t_L g6652 ( 
.A(n_6364),
.Y(n_6652)
);

OAI221xp5_ASAP7_75t_L g6653 ( 
.A1(n_6299),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.C(n_192),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_6329),
.Y(n_6654)
);

INVx1_ASAP7_75t_L g6655 ( 
.A(n_6336),
.Y(n_6655)
);

OAI22xp5_ASAP7_75t_L g6656 ( 
.A1(n_6364),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_6656)
);

AOI21xp5_ASAP7_75t_L g6657 ( 
.A1(n_6408),
.A2(n_193),
.B(n_194),
.Y(n_6657)
);

OAI33xp33_ASAP7_75t_L g6658 ( 
.A1(n_6488),
.A2(n_196),
.A3(n_198),
.B1(n_193),
.B2(n_195),
.B3(n_197),
.Y(n_6658)
);

AOI22xp33_ASAP7_75t_L g6659 ( 
.A1(n_6393),
.A2(n_1325),
.B1(n_1337),
.B2(n_1250),
.Y(n_6659)
);

A2O1A1Ixp33_ASAP7_75t_L g6660 ( 
.A1(n_6374),
.A2(n_200),
.B(n_196),
.C(n_199),
.Y(n_6660)
);

AOI22xp5_ASAP7_75t_L g6661 ( 
.A1(n_6501),
.A2(n_202),
.B1(n_199),
.B2(n_201),
.Y(n_6661)
);

NAND2xp5_ASAP7_75t_L g6662 ( 
.A(n_6337),
.B(n_203),
.Y(n_6662)
);

AOI22xp33_ASAP7_75t_L g6663 ( 
.A1(n_6394),
.A2(n_6396),
.B1(n_6404),
.B2(n_6402),
.Y(n_6663)
);

AOI22xp33_ASAP7_75t_L g6664 ( 
.A1(n_6500),
.A2(n_1337),
.B1(n_1341),
.B2(n_1250),
.Y(n_6664)
);

OAI22xp33_ASAP7_75t_L g6665 ( 
.A1(n_6395),
.A2(n_207),
.B1(n_204),
.B2(n_206),
.Y(n_6665)
);

INVx1_ASAP7_75t_L g6666 ( 
.A(n_6339),
.Y(n_6666)
);

AOI22xp33_ASAP7_75t_SL g6667 ( 
.A1(n_6338),
.A2(n_210),
.B1(n_206),
.B2(n_207),
.Y(n_6667)
);

CKINVDCx6p67_ASAP7_75t_R g6668 ( 
.A(n_6401),
.Y(n_6668)
);

AND2x4_ASAP7_75t_L g6669 ( 
.A(n_6403),
.B(n_210),
.Y(n_6669)
);

OAI22xp5_ASAP7_75t_L g6670 ( 
.A1(n_6354),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_6670)
);

AOI22xp33_ASAP7_75t_SL g6671 ( 
.A1(n_6338),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_6671)
);

AOI22xp33_ASAP7_75t_SL g6672 ( 
.A1(n_6453),
.A2(n_217),
.B1(n_214),
.B2(n_216),
.Y(n_6672)
);

AOI22xp33_ASAP7_75t_L g6673 ( 
.A1(n_6397),
.A2(n_1397),
.B1(n_1416),
.B2(n_1341),
.Y(n_6673)
);

AOI22xp33_ASAP7_75t_L g6674 ( 
.A1(n_6398),
.A2(n_1397),
.B1(n_1416),
.B2(n_1341),
.Y(n_6674)
);

OAI22xp5_ASAP7_75t_L g6675 ( 
.A1(n_6386),
.A2(n_220),
.B1(n_214),
.B2(n_217),
.Y(n_6675)
);

AOI221xp5_ASAP7_75t_L g6676 ( 
.A1(n_6453),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.C(n_224),
.Y(n_6676)
);

AOI22xp33_ASAP7_75t_L g6677 ( 
.A1(n_6383),
.A2(n_6385),
.B1(n_6476),
.B2(n_6468),
.Y(n_6677)
);

OR2x2_ASAP7_75t_L g6678 ( 
.A(n_6478),
.B(n_221),
.Y(n_6678)
);

INVx1_ASAP7_75t_L g6679 ( 
.A(n_6347),
.Y(n_6679)
);

AOI221xp5_ASAP7_75t_L g6680 ( 
.A1(n_6474),
.A2(n_227),
.B1(n_222),
.B2(n_226),
.C(n_230),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_6283),
.Y(n_6681)
);

INVx1_ASAP7_75t_L g6682 ( 
.A(n_6288),
.Y(n_6682)
);

OAI211xp5_ASAP7_75t_L g6683 ( 
.A1(n_6474),
.A2(n_231),
.B(n_226),
.C(n_230),
.Y(n_6683)
);

INVx3_ASAP7_75t_L g6684 ( 
.A(n_6348),
.Y(n_6684)
);

AOI21xp5_ASAP7_75t_L g6685 ( 
.A1(n_6375),
.A2(n_232),
.B(n_233),
.Y(n_6685)
);

AOI22xp33_ASAP7_75t_L g6686 ( 
.A1(n_6484),
.A2(n_1397),
.B1(n_1416),
.B2(n_1341),
.Y(n_6686)
);

NAND2xp5_ASAP7_75t_L g6687 ( 
.A(n_6289),
.B(n_234),
.Y(n_6687)
);

AOI22xp33_ASAP7_75t_L g6688 ( 
.A1(n_6497),
.A2(n_1397),
.B1(n_1416),
.B2(n_1341),
.Y(n_6688)
);

HB1xp67_ASAP7_75t_L g6689 ( 
.A(n_6469),
.Y(n_6689)
);

AOI222xp33_ASAP7_75t_L g6690 ( 
.A1(n_6413),
.A2(n_237),
.B1(n_239),
.B2(n_235),
.C1(n_236),
.C2(n_238),
.Y(n_6690)
);

BUFx6f_ASAP7_75t_L g6691 ( 
.A(n_6427),
.Y(n_6691)
);

INVx2_ASAP7_75t_L g6692 ( 
.A(n_6415),
.Y(n_6692)
);

BUFx2_ASAP7_75t_L g6693 ( 
.A(n_6416),
.Y(n_6693)
);

AOI222xp33_ASAP7_75t_L g6694 ( 
.A1(n_6413),
.A2(n_237),
.B1(n_240),
.B2(n_235),
.C1(n_236),
.C2(n_238),
.Y(n_6694)
);

OAI22xp5_ASAP7_75t_L g6695 ( 
.A1(n_6458),
.A2(n_243),
.B1(n_240),
.B2(n_241),
.Y(n_6695)
);

OAI211xp5_ASAP7_75t_SL g6696 ( 
.A1(n_6475),
.A2(n_245),
.B(n_241),
.C(n_244),
.Y(n_6696)
);

OAI211xp5_ASAP7_75t_L g6697 ( 
.A1(n_6459),
.A2(n_249),
.B(n_245),
.C(n_246),
.Y(n_6697)
);

OAI22xp5_ASAP7_75t_L g6698 ( 
.A1(n_6359),
.A2(n_253),
.B1(n_246),
.B2(n_250),
.Y(n_6698)
);

INVx1_ASAP7_75t_L g6699 ( 
.A(n_6295),
.Y(n_6699)
);

AOI22xp5_ASAP7_75t_L g6700 ( 
.A1(n_6296),
.A2(n_256),
.B1(n_253),
.B2(n_254),
.Y(n_6700)
);

AOI221xp5_ASAP7_75t_L g6701 ( 
.A1(n_6459),
.A2(n_258),
.B1(n_254),
.B2(n_257),
.C(n_259),
.Y(n_6701)
);

AND2x2_ASAP7_75t_SL g6702 ( 
.A(n_6361),
.B(n_257),
.Y(n_6702)
);

AND2x2_ASAP7_75t_L g6703 ( 
.A(n_6366),
.B(n_260),
.Y(n_6703)
);

AOI22xp5_ASAP7_75t_L g6704 ( 
.A1(n_6300),
.A2(n_264),
.B1(n_261),
.B2(n_263),
.Y(n_6704)
);

AOI22xp33_ASAP7_75t_L g6705 ( 
.A1(n_6379),
.A2(n_1416),
.B1(n_1422),
.B2(n_1397),
.Y(n_6705)
);

AOI22xp33_ASAP7_75t_L g6706 ( 
.A1(n_6387),
.A2(n_1422),
.B1(n_2792),
.B2(n_2775),
.Y(n_6706)
);

BUFx3_ASAP7_75t_L g6707 ( 
.A(n_6273),
.Y(n_6707)
);

AND2x2_ASAP7_75t_L g6708 ( 
.A(n_6481),
.B(n_263),
.Y(n_6708)
);

AOI22xp33_ASAP7_75t_L g6709 ( 
.A1(n_6485),
.A2(n_6493),
.B1(n_6502),
.B2(n_6489),
.Y(n_6709)
);

BUFx4f_ASAP7_75t_L g6710 ( 
.A(n_6361),
.Y(n_6710)
);

OAI22xp33_ASAP7_75t_L g6711 ( 
.A1(n_6428),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_6711)
);

HB1xp67_ASAP7_75t_L g6712 ( 
.A(n_6469),
.Y(n_6712)
);

INVx5_ASAP7_75t_SL g6713 ( 
.A(n_6454),
.Y(n_6713)
);

NAND3xp33_ASAP7_75t_L g6714 ( 
.A(n_6293),
.B(n_265),
.C(n_266),
.Y(n_6714)
);

AOI22xp33_ASAP7_75t_SL g6715 ( 
.A1(n_6293),
.A2(n_270),
.B1(n_267),
.B2(n_269),
.Y(n_6715)
);

HB1xp67_ASAP7_75t_L g6716 ( 
.A(n_6298),
.Y(n_6716)
);

AO21x2_ASAP7_75t_L g6717 ( 
.A1(n_6435),
.A2(n_269),
.B(n_271),
.Y(n_6717)
);

AOI22xp33_ASAP7_75t_SL g6718 ( 
.A1(n_6298),
.A2(n_6454),
.B1(n_6435),
.B2(n_6463),
.Y(n_6718)
);

OAI22xp5_ASAP7_75t_L g6719 ( 
.A1(n_6301),
.A2(n_276),
.B1(n_273),
.B2(n_274),
.Y(n_6719)
);

NAND3xp33_ASAP7_75t_L g6720 ( 
.A(n_6358),
.B(n_273),
.C(n_274),
.Y(n_6720)
);

INVx1_ASAP7_75t_L g6721 ( 
.A(n_6598),
.Y(n_6721)
);

NAND2xp5_ASAP7_75t_L g6722 ( 
.A(n_6535),
.B(n_6305),
.Y(n_6722)
);

INVx1_ASAP7_75t_L g6723 ( 
.A(n_6616),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_6619),
.Y(n_6724)
);

AND2x2_ASAP7_75t_L g6725 ( 
.A(n_6509),
.B(n_6512),
.Y(n_6725)
);

INVx2_ASAP7_75t_L g6726 ( 
.A(n_6504),
.Y(n_6726)
);

INVx2_ASAP7_75t_L g6727 ( 
.A(n_6504),
.Y(n_6727)
);

AND2x4_ASAP7_75t_L g6728 ( 
.A(n_6512),
.B(n_6306),
.Y(n_6728)
);

NOR2x1_ASAP7_75t_SL g6729 ( 
.A(n_6590),
.B(n_6470),
.Y(n_6729)
);

HB1xp67_ASAP7_75t_L g6730 ( 
.A(n_6716),
.Y(n_6730)
);

INVx1_ASAP7_75t_L g6731 ( 
.A(n_6689),
.Y(n_6731)
);

AND2x2_ASAP7_75t_L g6732 ( 
.A(n_6510),
.B(n_6409),
.Y(n_6732)
);

INVx1_ASAP7_75t_L g6733 ( 
.A(n_6712),
.Y(n_6733)
);

NAND2xp5_ASAP7_75t_L g6734 ( 
.A(n_6511),
.B(n_6309),
.Y(n_6734)
);

INVx1_ASAP7_75t_L g6735 ( 
.A(n_6566),
.Y(n_6735)
);

NAND2x1_ASAP7_75t_L g6736 ( 
.A(n_6533),
.B(n_6310),
.Y(n_6736)
);

NAND2xp5_ASAP7_75t_L g6737 ( 
.A(n_6514),
.B(n_6312),
.Y(n_6737)
);

INVx1_ASAP7_75t_L g6738 ( 
.A(n_6566),
.Y(n_6738)
);

AND2x2_ASAP7_75t_L g6739 ( 
.A(n_6634),
.B(n_6412),
.Y(n_6739)
);

HB1xp67_ASAP7_75t_L g6740 ( 
.A(n_6643),
.Y(n_6740)
);

OR2x2_ASAP7_75t_L g6741 ( 
.A(n_6568),
.B(n_6357),
.Y(n_6741)
);

INVx1_ASAP7_75t_L g6742 ( 
.A(n_6569),
.Y(n_6742)
);

AND2x2_ASAP7_75t_L g6743 ( 
.A(n_6636),
.B(n_6437),
.Y(n_6743)
);

INVx2_ASAP7_75t_L g6744 ( 
.A(n_6567),
.Y(n_6744)
);

AND2x2_ASAP7_75t_L g6745 ( 
.A(n_6652),
.B(n_6438),
.Y(n_6745)
);

INVx1_ASAP7_75t_L g6746 ( 
.A(n_6569),
.Y(n_6746)
);

HB1xp67_ASAP7_75t_L g6747 ( 
.A(n_6643),
.Y(n_6747)
);

HB1xp67_ASAP7_75t_L g6748 ( 
.A(n_6717),
.Y(n_6748)
);

NAND3xp33_ASAP7_75t_L g6749 ( 
.A(n_6599),
.B(n_6463),
.C(n_6358),
.Y(n_6749)
);

NAND2xp5_ASAP7_75t_L g6750 ( 
.A(n_6522),
.B(n_6315),
.Y(n_6750)
);

INVxp67_ASAP7_75t_L g6751 ( 
.A(n_6521),
.Y(n_6751)
);

INVx1_ASAP7_75t_L g6752 ( 
.A(n_6523),
.Y(n_6752)
);

AND2x2_ASAP7_75t_L g6753 ( 
.A(n_6652),
.B(n_6638),
.Y(n_6753)
);

INVx2_ASAP7_75t_L g6754 ( 
.A(n_6684),
.Y(n_6754)
);

NOR2xp33_ASAP7_75t_L g6755 ( 
.A(n_6532),
.B(n_6316),
.Y(n_6755)
);

INVxp67_ASAP7_75t_L g6756 ( 
.A(n_6604),
.Y(n_6756)
);

INVx1_ASAP7_75t_L g6757 ( 
.A(n_6534),
.Y(n_6757)
);

INVx1_ASAP7_75t_L g6758 ( 
.A(n_6537),
.Y(n_6758)
);

NAND2x1p5_ASAP7_75t_L g6759 ( 
.A(n_6581),
.B(n_6344),
.Y(n_6759)
);

INVx2_ASAP7_75t_L g6760 ( 
.A(n_6713),
.Y(n_6760)
);

INVx1_ASAP7_75t_L g6761 ( 
.A(n_6552),
.Y(n_6761)
);

NAND2x1_ASAP7_75t_L g6762 ( 
.A(n_6600),
.B(n_6318),
.Y(n_6762)
);

AND2x2_ASAP7_75t_L g6763 ( 
.A(n_6638),
.B(n_6622),
.Y(n_6763)
);

HB1xp67_ASAP7_75t_L g6764 ( 
.A(n_6717),
.Y(n_6764)
);

AND2x2_ASAP7_75t_L g6765 ( 
.A(n_6622),
.B(n_6446),
.Y(n_6765)
);

INVx3_ASAP7_75t_L g6766 ( 
.A(n_6586),
.Y(n_6766)
);

INVx3_ASAP7_75t_L g6767 ( 
.A(n_6586),
.Y(n_6767)
);

AND2x2_ASAP7_75t_L g6768 ( 
.A(n_6640),
.B(n_6447),
.Y(n_6768)
);

AND2x2_ASAP7_75t_L g6769 ( 
.A(n_6547),
.B(n_6455),
.Y(n_6769)
);

HB1xp67_ASAP7_75t_L g6770 ( 
.A(n_6604),
.Y(n_6770)
);

AND2x2_ASAP7_75t_L g6771 ( 
.A(n_6564),
.B(n_6360),
.Y(n_6771)
);

AND2x2_ASAP7_75t_L g6772 ( 
.A(n_6668),
.B(n_6371),
.Y(n_6772)
);

AND2x2_ASAP7_75t_L g6773 ( 
.A(n_6693),
.B(n_6372),
.Y(n_6773)
);

NOR2x1_ASAP7_75t_L g6774 ( 
.A(n_6573),
.B(n_6322),
.Y(n_6774)
);

INVx2_ASAP7_75t_SL g6775 ( 
.A(n_6532),
.Y(n_6775)
);

BUFx2_ASAP7_75t_L g6776 ( 
.A(n_6590),
.Y(n_6776)
);

AND2x2_ASAP7_75t_L g6777 ( 
.A(n_6536),
.B(n_6376),
.Y(n_6777)
);

AND2x2_ASAP7_75t_L g6778 ( 
.A(n_6583),
.B(n_6378),
.Y(n_6778)
);

INVx2_ASAP7_75t_L g6779 ( 
.A(n_6532),
.Y(n_6779)
);

AND2x2_ASAP7_75t_L g6780 ( 
.A(n_6617),
.B(n_6418),
.Y(n_6780)
);

AND2x2_ASAP7_75t_L g6781 ( 
.A(n_6624),
.B(n_6419),
.Y(n_6781)
);

AND2x2_ASAP7_75t_L g6782 ( 
.A(n_6630),
.B(n_6420),
.Y(n_6782)
);

INVx3_ASAP7_75t_L g6783 ( 
.A(n_6691),
.Y(n_6783)
);

INVx2_ASAP7_75t_L g6784 ( 
.A(n_6691),
.Y(n_6784)
);

INVx1_ASAP7_75t_L g6785 ( 
.A(n_6560),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_6654),
.Y(n_6786)
);

BUFx3_ASAP7_75t_L g6787 ( 
.A(n_6520),
.Y(n_6787)
);

AND2x2_ASAP7_75t_L g6788 ( 
.A(n_6632),
.B(n_6422),
.Y(n_6788)
);

AND2x2_ASAP7_75t_L g6789 ( 
.A(n_6651),
.B(n_6425),
.Y(n_6789)
);

AND2x4_ASAP7_75t_L g6790 ( 
.A(n_6613),
.B(n_6527),
.Y(n_6790)
);

NAND2xp5_ASAP7_75t_L g6791 ( 
.A(n_6529),
.B(n_6325),
.Y(n_6791)
);

NAND2xp5_ASAP7_75t_L g6792 ( 
.A(n_6516),
.B(n_6326),
.Y(n_6792)
);

INVx1_ASAP7_75t_L g6793 ( 
.A(n_6654),
.Y(n_6793)
);

NOR2x1_ASAP7_75t_L g6794 ( 
.A(n_6613),
.B(n_6351),
.Y(n_6794)
);

INVx1_ASAP7_75t_L g6795 ( 
.A(n_6606),
.Y(n_6795)
);

BUFx3_ASAP7_75t_L g6796 ( 
.A(n_6633),
.Y(n_6796)
);

AND2x2_ASAP7_75t_L g6797 ( 
.A(n_6527),
.B(n_6433),
.Y(n_6797)
);

NAND2xp5_ASAP7_75t_L g6798 ( 
.A(n_6601),
.B(n_6353),
.Y(n_6798)
);

NAND2xp5_ASAP7_75t_L g6799 ( 
.A(n_6657),
.B(n_6355),
.Y(n_6799)
);

AND2x2_ASAP7_75t_L g6800 ( 
.A(n_6639),
.B(n_6498),
.Y(n_6800)
);

INVx2_ASAP7_75t_L g6801 ( 
.A(n_6707),
.Y(n_6801)
);

AND2x2_ASAP7_75t_L g6802 ( 
.A(n_6642),
.B(n_6460),
.Y(n_6802)
);

AO21x2_ASAP7_75t_L g6803 ( 
.A1(n_6541),
.A2(n_6464),
.B(n_6462),
.Y(n_6803)
);

HB1xp67_ASAP7_75t_L g6804 ( 
.A(n_6505),
.Y(n_6804)
);

HB1xp67_ASAP7_75t_L g6805 ( 
.A(n_6505),
.Y(n_6805)
);

INVx1_ASAP7_75t_L g6806 ( 
.A(n_6615),
.Y(n_6806)
);

OR2x2_ASAP7_75t_L g6807 ( 
.A(n_6692),
.B(n_6475),
.Y(n_6807)
);

INVx1_ASAP7_75t_L g6808 ( 
.A(n_6625),
.Y(n_6808)
);

HB1xp67_ASAP7_75t_L g6809 ( 
.A(n_6720),
.Y(n_6809)
);

BUFx3_ASAP7_75t_L g6810 ( 
.A(n_6562),
.Y(n_6810)
);

INVx1_ASAP7_75t_L g6811 ( 
.A(n_6635),
.Y(n_6811)
);

OAI21xp33_ASAP7_75t_L g6812 ( 
.A1(n_6503),
.A2(n_6486),
.B(n_6477),
.Y(n_6812)
);

INVx1_ASAP7_75t_L g6813 ( 
.A(n_6647),
.Y(n_6813)
);

INVx2_ASAP7_75t_L g6814 ( 
.A(n_6575),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_6579),
.Y(n_6815)
);

AND2x2_ASAP7_75t_L g6816 ( 
.A(n_6649),
.B(n_6471),
.Y(n_6816)
);

AND2x2_ASAP7_75t_L g6817 ( 
.A(n_6650),
.B(n_6480),
.Y(n_6817)
);

BUFx3_ASAP7_75t_L g6818 ( 
.A(n_6562),
.Y(n_6818)
);

INVx1_ASAP7_75t_L g6819 ( 
.A(n_6655),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_6666),
.Y(n_6820)
);

INVx2_ASAP7_75t_L g6821 ( 
.A(n_6713),
.Y(n_6821)
);

INVx2_ASAP7_75t_L g6822 ( 
.A(n_6702),
.Y(n_6822)
);

INVx2_ASAP7_75t_L g6823 ( 
.A(n_6669),
.Y(n_6823)
);

INVx2_ASAP7_75t_L g6824 ( 
.A(n_6669),
.Y(n_6824)
);

INVx1_ASAP7_75t_L g6825 ( 
.A(n_6679),
.Y(n_6825)
);

AND2x2_ASAP7_75t_L g6826 ( 
.A(n_6524),
.B(n_6368),
.Y(n_6826)
);

INVx2_ASAP7_75t_L g6827 ( 
.A(n_6506),
.Y(n_6827)
);

BUFx3_ASAP7_75t_L g6828 ( 
.A(n_6585),
.Y(n_6828)
);

AND2x2_ASAP7_75t_L g6829 ( 
.A(n_6526),
.B(n_6368),
.Y(n_6829)
);

AND2x4_ASAP7_75t_L g6830 ( 
.A(n_6585),
.B(n_6286),
.Y(n_6830)
);

OR2x2_ASAP7_75t_L g6831 ( 
.A(n_6584),
.B(n_6465),
.Y(n_6831)
);

INVx2_ASAP7_75t_L g6832 ( 
.A(n_6610),
.Y(n_6832)
);

AND2x4_ASAP7_75t_L g6833 ( 
.A(n_6610),
.B(n_6494),
.Y(n_6833)
);

AND2x2_ASAP7_75t_L g6834 ( 
.A(n_6526),
.B(n_277),
.Y(n_6834)
);

NAND2xp5_ASAP7_75t_L g6835 ( 
.A(n_6681),
.B(n_277),
.Y(n_6835)
);

INVx1_ASAP7_75t_L g6836 ( 
.A(n_6682),
.Y(n_6836)
);

AND2x2_ASAP7_75t_SL g6837 ( 
.A(n_6710),
.B(n_278),
.Y(n_6837)
);

INVx2_ASAP7_75t_L g6838 ( 
.A(n_6517),
.Y(n_6838)
);

INVx1_ASAP7_75t_L g6839 ( 
.A(n_6699),
.Y(n_6839)
);

INVx2_ASAP7_75t_L g6840 ( 
.A(n_6517),
.Y(n_6840)
);

AND2x2_ASAP7_75t_L g6841 ( 
.A(n_6607),
.B(n_279),
.Y(n_6841)
);

INVx3_ASAP7_75t_L g6842 ( 
.A(n_6517),
.Y(n_6842)
);

AND2x2_ASAP7_75t_L g6843 ( 
.A(n_6626),
.B(n_6559),
.Y(n_6843)
);

INVx2_ASAP7_75t_L g6844 ( 
.A(n_6710),
.Y(n_6844)
);

INVx1_ASAP7_75t_L g6845 ( 
.A(n_6678),
.Y(n_6845)
);

NOR2xp33_ASAP7_75t_L g6846 ( 
.A(n_6570),
.B(n_6538),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_6594),
.Y(n_6847)
);

INVx5_ASAP7_75t_L g6848 ( 
.A(n_6628),
.Y(n_6848)
);

HB1xp67_ASAP7_75t_L g6849 ( 
.A(n_6714),
.Y(n_6849)
);

OR2x2_ASAP7_75t_L g6850 ( 
.A(n_6531),
.B(n_280),
.Y(n_6850)
);

INVxp67_ASAP7_75t_L g6851 ( 
.A(n_6549),
.Y(n_6851)
);

BUFx6f_ASAP7_75t_L g6852 ( 
.A(n_6631),
.Y(n_6852)
);

HB1xp67_ASAP7_75t_L g6853 ( 
.A(n_6558),
.Y(n_6853)
);

INVx1_ASAP7_75t_L g6854 ( 
.A(n_6687),
.Y(n_6854)
);

NOR2x1_ASAP7_75t_SL g6855 ( 
.A(n_6528),
.B(n_280),
.Y(n_6855)
);

AND2x2_ASAP7_75t_L g6856 ( 
.A(n_6580),
.B(n_281),
.Y(n_6856)
);

INVx8_ASAP7_75t_L g6857 ( 
.A(n_6708),
.Y(n_6857)
);

BUFx2_ASAP7_75t_L g6858 ( 
.A(n_6561),
.Y(n_6858)
);

AND2x2_ASAP7_75t_L g6859 ( 
.A(n_6609),
.B(n_281),
.Y(n_6859)
);

HB1xp67_ASAP7_75t_L g6860 ( 
.A(n_6577),
.Y(n_6860)
);

AND2x2_ASAP7_75t_L g6861 ( 
.A(n_6612),
.B(n_282),
.Y(n_6861)
);

AND2x2_ASAP7_75t_L g6862 ( 
.A(n_6530),
.B(n_282),
.Y(n_6862)
);

AND2x4_ASAP7_75t_L g6863 ( 
.A(n_6703),
.B(n_283),
.Y(n_6863)
);

INVx1_ASAP7_75t_L g6864 ( 
.A(n_6641),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_6646),
.Y(n_6865)
);

BUFx6f_ASAP7_75t_L g6866 ( 
.A(n_6623),
.Y(n_6866)
);

AND2x2_ASAP7_75t_L g6867 ( 
.A(n_6508),
.B(n_284),
.Y(n_6867)
);

AND2x4_ASAP7_75t_L g6868 ( 
.A(n_6546),
.B(n_285),
.Y(n_6868)
);

AND2x4_ASAP7_75t_L g6869 ( 
.A(n_6507),
.B(n_286),
.Y(n_6869)
);

AND2x2_ASAP7_75t_L g6870 ( 
.A(n_6709),
.B(n_6525),
.Y(n_6870)
);

OR2x2_ASAP7_75t_L g6871 ( 
.A(n_6662),
.B(n_289),
.Y(n_6871)
);

AND2x2_ASAP7_75t_L g6872 ( 
.A(n_6513),
.B(n_289),
.Y(n_6872)
);

INVx2_ASAP7_75t_L g6873 ( 
.A(n_6554),
.Y(n_6873)
);

INVxp67_ASAP7_75t_L g6874 ( 
.A(n_6553),
.Y(n_6874)
);

INVx1_ASAP7_75t_L g6875 ( 
.A(n_6677),
.Y(n_6875)
);

HB1xp67_ASAP7_75t_L g6876 ( 
.A(n_6695),
.Y(n_6876)
);

AND2x2_ASAP7_75t_L g6877 ( 
.A(n_6518),
.B(n_290),
.Y(n_6877)
);

INVx1_ASAP7_75t_L g6878 ( 
.A(n_6574),
.Y(n_6878)
);

HB1xp67_ASAP7_75t_L g6879 ( 
.A(n_6582),
.Y(n_6879)
);

HB1xp67_ASAP7_75t_L g6880 ( 
.A(n_6542),
.Y(n_6880)
);

NAND2xp5_ASAP7_75t_L g6881 ( 
.A(n_6603),
.B(n_290),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_6683),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_6719),
.Y(n_6883)
);

AOI22xp33_ASAP7_75t_SL g6884 ( 
.A1(n_6544),
.A2(n_296),
.B1(n_293),
.B2(n_295),
.Y(n_6884)
);

INVx1_ASAP7_75t_L g6885 ( 
.A(n_6670),
.Y(n_6885)
);

INVx2_ASAP7_75t_L g6886 ( 
.A(n_6551),
.Y(n_6886)
);

INVxp67_ASAP7_75t_SL g6887 ( 
.A(n_6718),
.Y(n_6887)
);

AND2x2_ASAP7_75t_L g6888 ( 
.A(n_6543),
.B(n_293),
.Y(n_6888)
);

AND2x4_ASAP7_75t_L g6889 ( 
.A(n_6515),
.B(n_295),
.Y(n_6889)
);

OR2x2_ASAP7_75t_L g6890 ( 
.A(n_6663),
.B(n_297),
.Y(n_6890)
);

NAND2xp5_ASAP7_75t_L g6891 ( 
.A(n_6667),
.B(n_297),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_6675),
.Y(n_6892)
);

NAND2xp5_ASAP7_75t_L g6893 ( 
.A(n_6887),
.B(n_6690),
.Y(n_6893)
);

AND2x2_ASAP7_75t_L g6894 ( 
.A(n_6787),
.B(n_6592),
.Y(n_6894)
);

OR2x2_ASAP7_75t_L g6895 ( 
.A(n_6822),
.B(n_6519),
.Y(n_6895)
);

AOI22xp33_ASAP7_75t_SL g6896 ( 
.A1(n_6889),
.A2(n_6608),
.B1(n_6629),
.B2(n_6593),
.Y(n_6896)
);

NOR2xp33_ASAP7_75t_L g6897 ( 
.A(n_6751),
.B(n_6565),
.Y(n_6897)
);

INVx2_ASAP7_75t_L g6898 ( 
.A(n_6790),
.Y(n_6898)
);

BUFx3_ASAP7_75t_L g6899 ( 
.A(n_6790),
.Y(n_6899)
);

INVx1_ASAP7_75t_L g6900 ( 
.A(n_6730),
.Y(n_6900)
);

AND2x2_ASAP7_75t_L g6901 ( 
.A(n_6763),
.B(n_6563),
.Y(n_6901)
);

BUFx2_ASAP7_75t_SL g6902 ( 
.A(n_6775),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6730),
.Y(n_6903)
);

AND2x2_ASAP7_75t_L g6904 ( 
.A(n_6753),
.B(n_6539),
.Y(n_6904)
);

OAI222xp33_ASAP7_75t_L g6905 ( 
.A1(n_6887),
.A2(n_6671),
.B1(n_6715),
.B2(n_6711),
.C1(n_6602),
.C2(n_6587),
.Y(n_6905)
);

AND2x2_ASAP7_75t_L g6906 ( 
.A(n_6766),
.B(n_6548),
.Y(n_6906)
);

INVx1_ASAP7_75t_L g6907 ( 
.A(n_6748),
.Y(n_6907)
);

BUFx6f_ASAP7_75t_L g6908 ( 
.A(n_6796),
.Y(n_6908)
);

AND2x2_ASAP7_75t_L g6909 ( 
.A(n_6766),
.B(n_6540),
.Y(n_6909)
);

INVxp67_ASAP7_75t_SL g6910 ( 
.A(n_6804),
.Y(n_6910)
);

AND2x2_ASAP7_75t_L g6911 ( 
.A(n_6767),
.B(n_6685),
.Y(n_6911)
);

INVx1_ASAP7_75t_L g6912 ( 
.A(n_6748),
.Y(n_6912)
);

AND2x4_ASAP7_75t_SL g6913 ( 
.A(n_6767),
.B(n_6661),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_6764),
.Y(n_6914)
);

INVx2_ASAP7_75t_L g6915 ( 
.A(n_6810),
.Y(n_6915)
);

AOI222xp33_ASAP7_75t_L g6916 ( 
.A1(n_6846),
.A2(n_6676),
.B1(n_6591),
.B2(n_6572),
.C1(n_6596),
.C2(n_6680),
.Y(n_6916)
);

NOR2xp67_ASAP7_75t_L g6917 ( 
.A(n_6751),
.B(n_6697),
.Y(n_6917)
);

INVx1_ASAP7_75t_L g6918 ( 
.A(n_6764),
.Y(n_6918)
);

INVx2_ASAP7_75t_SL g6919 ( 
.A(n_6810),
.Y(n_6919)
);

OR2x2_ASAP7_75t_L g6920 ( 
.A(n_6822),
.B(n_6589),
.Y(n_6920)
);

HB1xp67_ASAP7_75t_L g6921 ( 
.A(n_6774),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6770),
.Y(n_6922)
);

AOI22xp33_ASAP7_75t_L g6923 ( 
.A1(n_6889),
.A2(n_6696),
.B1(n_6595),
.B2(n_6701),
.Y(n_6923)
);

HB1xp67_ASAP7_75t_L g6924 ( 
.A(n_6804),
.Y(n_6924)
);

NAND2xp5_ASAP7_75t_L g6925 ( 
.A(n_6805),
.B(n_6694),
.Y(n_6925)
);

AND2x2_ASAP7_75t_L g6926 ( 
.A(n_6725),
.B(n_6744),
.Y(n_6926)
);

OR2x2_ASAP7_75t_L g6927 ( 
.A(n_6791),
.B(n_6656),
.Y(n_6927)
);

INVx2_ASAP7_75t_L g6928 ( 
.A(n_6818),
.Y(n_6928)
);

AND2x2_ASAP7_75t_L g6929 ( 
.A(n_6776),
.B(n_6621),
.Y(n_6929)
);

INVx2_ASAP7_75t_L g6930 ( 
.A(n_6818),
.Y(n_6930)
);

INVx1_ASAP7_75t_L g6931 ( 
.A(n_6740),
.Y(n_6931)
);

AND2x2_ASAP7_75t_L g6932 ( 
.A(n_6843),
.B(n_6576),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_6740),
.Y(n_6933)
);

BUFx2_ASAP7_75t_L g6934 ( 
.A(n_6828),
.Y(n_6934)
);

INVx1_ASAP7_75t_L g6935 ( 
.A(n_6747),
.Y(n_6935)
);

AND2x2_ASAP7_75t_L g6936 ( 
.A(n_6848),
.B(n_6620),
.Y(n_6936)
);

INVx2_ASAP7_75t_SL g6937 ( 
.A(n_6736),
.Y(n_6937)
);

INVx1_ASAP7_75t_L g6938 ( 
.A(n_6747),
.Y(n_6938)
);

AND2x2_ASAP7_75t_L g6939 ( 
.A(n_6848),
.B(n_6672),
.Y(n_6939)
);

AND2x4_ASAP7_75t_L g6940 ( 
.A(n_6779),
.B(n_6660),
.Y(n_6940)
);

HB1xp67_ASAP7_75t_L g6941 ( 
.A(n_6805),
.Y(n_6941)
);

AOI22xp33_ASAP7_75t_L g6942 ( 
.A1(n_6846),
.A2(n_6884),
.B1(n_6870),
.B2(n_6876),
.Y(n_6942)
);

INVx2_ASAP7_75t_SL g6943 ( 
.A(n_6848),
.Y(n_6943)
);

AOI22xp33_ASAP7_75t_L g6944 ( 
.A1(n_6884),
.A2(n_6658),
.B1(n_6597),
.B2(n_6556),
.Y(n_6944)
);

INVx1_ASAP7_75t_SL g6945 ( 
.A(n_6837),
.Y(n_6945)
);

HB1xp67_ASAP7_75t_L g6946 ( 
.A(n_6756),
.Y(n_6946)
);

INVx1_ASAP7_75t_L g6947 ( 
.A(n_6735),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_6738),
.Y(n_6948)
);

INVx1_ASAP7_75t_L g6949 ( 
.A(n_6742),
.Y(n_6949)
);

INVx1_ASAP7_75t_L g6950 ( 
.A(n_6746),
.Y(n_6950)
);

INVx2_ASAP7_75t_L g6951 ( 
.A(n_6866),
.Y(n_6951)
);

AND2x2_ASAP7_75t_L g6952 ( 
.A(n_6848),
.B(n_6698),
.Y(n_6952)
);

INVxp67_ASAP7_75t_L g6953 ( 
.A(n_6879),
.Y(n_6953)
);

AND2x2_ASAP7_75t_L g6954 ( 
.A(n_6726),
.B(n_6700),
.Y(n_6954)
);

OR2x2_ASAP7_75t_L g6955 ( 
.A(n_6791),
.B(n_6849),
.Y(n_6955)
);

BUFx3_ASAP7_75t_L g6956 ( 
.A(n_6852),
.Y(n_6956)
);

INVx1_ASAP7_75t_SL g6957 ( 
.A(n_6837),
.Y(n_6957)
);

OR2x2_ASAP7_75t_L g6958 ( 
.A(n_6849),
.B(n_6665),
.Y(n_6958)
);

AND2x2_ASAP7_75t_L g6959 ( 
.A(n_6727),
.B(n_6832),
.Y(n_6959)
);

INVx2_ASAP7_75t_L g6960 ( 
.A(n_6866),
.Y(n_6960)
);

OR2x2_ASAP7_75t_L g6961 ( 
.A(n_6823),
.B(n_6645),
.Y(n_6961)
);

AND2x2_ASAP7_75t_L g6962 ( 
.A(n_6772),
.B(n_6704),
.Y(n_6962)
);

AND2x2_ASAP7_75t_L g6963 ( 
.A(n_6824),
.B(n_6578),
.Y(n_6963)
);

NAND2xp5_ASAP7_75t_L g6964 ( 
.A(n_6809),
.B(n_6614),
.Y(n_6964)
);

AND2x2_ASAP7_75t_L g6965 ( 
.A(n_6866),
.B(n_6588),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6721),
.Y(n_6966)
);

INVx2_ASAP7_75t_L g6967 ( 
.A(n_6852),
.Y(n_6967)
);

INVx2_ASAP7_75t_L g6968 ( 
.A(n_6852),
.Y(n_6968)
);

NOR2xp33_ASAP7_75t_L g6969 ( 
.A(n_6851),
.B(n_6783),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6723),
.Y(n_6970)
);

NOR2xp67_ASAP7_75t_L g6971 ( 
.A(n_6783),
.B(n_6550),
.Y(n_6971)
);

OR2x2_ASAP7_75t_SL g6972 ( 
.A(n_6879),
.B(n_6618),
.Y(n_6972)
);

INVxp67_ASAP7_75t_SL g6973 ( 
.A(n_6756),
.Y(n_6973)
);

INVx1_ASAP7_75t_L g6974 ( 
.A(n_6724),
.Y(n_6974)
);

CKINVDCx16_ASAP7_75t_R g6975 ( 
.A(n_6834),
.Y(n_6975)
);

AND2x2_ASAP7_75t_L g6976 ( 
.A(n_6784),
.B(n_6605),
.Y(n_6976)
);

AND2x4_ASAP7_75t_L g6977 ( 
.A(n_6794),
.B(n_6571),
.Y(n_6977)
);

OR2x2_ASAP7_75t_L g6978 ( 
.A(n_6809),
.B(n_6611),
.Y(n_6978)
);

INVx1_ASAP7_75t_L g6979 ( 
.A(n_6731),
.Y(n_6979)
);

INVx1_ASAP7_75t_L g6980 ( 
.A(n_6733),
.Y(n_6980)
);

AND2x4_ASAP7_75t_L g6981 ( 
.A(n_6797),
.B(n_6706),
.Y(n_6981)
);

NAND2xp5_ASAP7_75t_L g6982 ( 
.A(n_6881),
.B(n_6644),
.Y(n_6982)
);

AND2x2_ASAP7_75t_L g6983 ( 
.A(n_6732),
.B(n_6627),
.Y(n_6983)
);

OAI22xp5_ASAP7_75t_L g6984 ( 
.A1(n_6749),
.A2(n_6653),
.B1(n_6545),
.B2(n_6659),
.Y(n_6984)
);

INVx1_ASAP7_75t_L g6985 ( 
.A(n_6786),
.Y(n_6985)
);

NAND2xp5_ASAP7_75t_L g6986 ( 
.A(n_6881),
.B(n_6673),
.Y(n_6986)
);

NAND2xp5_ASAP7_75t_L g6987 ( 
.A(n_6878),
.B(n_6674),
.Y(n_6987)
);

INVx2_ASAP7_75t_L g6988 ( 
.A(n_6754),
.Y(n_6988)
);

AND2x2_ASAP7_75t_L g6989 ( 
.A(n_6855),
.B(n_6555),
.Y(n_6989)
);

BUFx3_ASAP7_75t_L g6990 ( 
.A(n_6857),
.Y(n_6990)
);

BUFx2_ASAP7_75t_L g6991 ( 
.A(n_6754),
.Y(n_6991)
);

OR2x2_ASAP7_75t_L g6992 ( 
.A(n_6851),
.B(n_6705),
.Y(n_6992)
);

BUFx5_ASAP7_75t_L g6993 ( 
.A(n_6867),
.Y(n_6993)
);

HB1xp67_ASAP7_75t_L g6994 ( 
.A(n_6876),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6793),
.Y(n_6995)
);

AND2x2_ASAP7_75t_L g6996 ( 
.A(n_6768),
.B(n_6648),
.Y(n_6996)
);

NAND2xp5_ASAP7_75t_L g6997 ( 
.A(n_6874),
.B(n_6882),
.Y(n_6997)
);

BUFx2_ASAP7_75t_L g6998 ( 
.A(n_6765),
.Y(n_6998)
);

NAND2xp5_ASAP7_75t_L g6999 ( 
.A(n_6874),
.B(n_6664),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6845),
.Y(n_7000)
);

NAND2xp5_ASAP7_75t_L g7001 ( 
.A(n_6869),
.B(n_6858),
.Y(n_7001)
);

HB1xp67_ASAP7_75t_L g7002 ( 
.A(n_6853),
.Y(n_7002)
);

NOR3xp33_ASAP7_75t_L g7003 ( 
.A(n_6841),
.B(n_298),
.C(n_300),
.Y(n_7003)
);

NAND2xp33_ASAP7_75t_SL g7004 ( 
.A(n_6829),
.B(n_6637),
.Y(n_7004)
);

AND2x2_ASAP7_75t_L g7005 ( 
.A(n_6801),
.B(n_6686),
.Y(n_7005)
);

AND2x2_ASAP7_75t_L g7006 ( 
.A(n_6771),
.B(n_6688),
.Y(n_7006)
);

NAND2xp5_ASAP7_75t_L g7007 ( 
.A(n_6869),
.B(n_6885),
.Y(n_7007)
);

AND2x2_ASAP7_75t_L g7008 ( 
.A(n_6769),
.B(n_6557),
.Y(n_7008)
);

INVx1_ASAP7_75t_L g7009 ( 
.A(n_6847),
.Y(n_7009)
);

INVx2_ASAP7_75t_L g7010 ( 
.A(n_6762),
.Y(n_7010)
);

INVx1_ASAP7_75t_L g7011 ( 
.A(n_6752),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6757),
.Y(n_7012)
);

NAND2xp5_ASAP7_75t_L g7013 ( 
.A(n_6892),
.B(n_300),
.Y(n_7013)
);

INVx1_ASAP7_75t_L g7014 ( 
.A(n_6758),
.Y(n_7014)
);

INVx1_ASAP7_75t_L g7015 ( 
.A(n_6761),
.Y(n_7015)
);

AOI22xp33_ASAP7_75t_L g7016 ( 
.A1(n_6875),
.A2(n_6749),
.B1(n_6722),
.B2(n_6792),
.Y(n_7016)
);

INVx2_ASAP7_75t_L g7017 ( 
.A(n_6857),
.Y(n_7017)
);

AND2x2_ASAP7_75t_L g7018 ( 
.A(n_6880),
.B(n_301),
.Y(n_7018)
);

INVx1_ASAP7_75t_L g7019 ( 
.A(n_6785),
.Y(n_7019)
);

AOI22xp33_ASAP7_75t_L g7020 ( 
.A1(n_6722),
.A2(n_1422),
.B1(n_2925),
.B2(n_2792),
.Y(n_7020)
);

HB1xp67_ASAP7_75t_L g7021 ( 
.A(n_6853),
.Y(n_7021)
);

NOR2xp33_ASAP7_75t_L g7022 ( 
.A(n_6871),
.B(n_302),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_6734),
.Y(n_7023)
);

OR2x2_ASAP7_75t_L g7024 ( 
.A(n_6883),
.B(n_302),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6924),
.Y(n_7025)
);

INVx3_ASAP7_75t_L g7026 ( 
.A(n_6899),
.Y(n_7026)
);

AND2x2_ASAP7_75t_L g7027 ( 
.A(n_6894),
.B(n_6739),
.Y(n_7027)
);

OR2x2_ASAP7_75t_L g7028 ( 
.A(n_6945),
.B(n_6798),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6924),
.Y(n_7029)
);

OR2x2_ASAP7_75t_L g7030 ( 
.A(n_6945),
.B(n_6798),
.Y(n_7030)
);

AND2x2_ASAP7_75t_L g7031 ( 
.A(n_6898),
.B(n_6728),
.Y(n_7031)
);

INVx2_ASAP7_75t_L g7032 ( 
.A(n_6943),
.Y(n_7032)
);

AND2x4_ASAP7_75t_L g7033 ( 
.A(n_6937),
.B(n_6728),
.Y(n_7033)
);

OR2x2_ASAP7_75t_L g7034 ( 
.A(n_6957),
.B(n_6799),
.Y(n_7034)
);

AND2x2_ASAP7_75t_L g7035 ( 
.A(n_6998),
.B(n_6926),
.Y(n_7035)
);

HB1xp67_ASAP7_75t_L g7036 ( 
.A(n_6941),
.Y(n_7036)
);

INVxp67_ASAP7_75t_L g7037 ( 
.A(n_6994),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6941),
.Y(n_7038)
);

INVx2_ASAP7_75t_L g7039 ( 
.A(n_6908),
.Y(n_7039)
);

INVx1_ASAP7_75t_L g7040 ( 
.A(n_6910),
.Y(n_7040)
);

NAND2xp5_ASAP7_75t_L g7041 ( 
.A(n_6942),
.B(n_6792),
.Y(n_7041)
);

INVx2_ASAP7_75t_L g7042 ( 
.A(n_6908),
.Y(n_7042)
);

INVx1_ASAP7_75t_L g7043 ( 
.A(n_6910),
.Y(n_7043)
);

INVx5_ASAP7_75t_SL g7044 ( 
.A(n_6908),
.Y(n_7044)
);

INVx1_ASAP7_75t_L g7045 ( 
.A(n_6946),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_6900),
.Y(n_7046)
);

INVx1_ASAP7_75t_L g7047 ( 
.A(n_6903),
.Y(n_7047)
);

OR2x2_ASAP7_75t_L g7048 ( 
.A(n_6957),
.B(n_6799),
.Y(n_7048)
);

AND2x2_ASAP7_75t_L g7049 ( 
.A(n_6911),
.B(n_6888),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_7002),
.Y(n_7050)
);

AND2x2_ASAP7_75t_L g7051 ( 
.A(n_6904),
.B(n_6773),
.Y(n_7051)
);

INVx2_ASAP7_75t_L g7052 ( 
.A(n_6934),
.Y(n_7052)
);

AOI22xp33_ASAP7_75t_SL g7053 ( 
.A1(n_6893),
.A2(n_6729),
.B1(n_6872),
.B2(n_6860),
.Y(n_7053)
);

HB1xp67_ASAP7_75t_L g7054 ( 
.A(n_6994),
.Y(n_7054)
);

NAND2xp5_ASAP7_75t_L g7055 ( 
.A(n_7016),
.B(n_6864),
.Y(n_7055)
);

HB1xp67_ASAP7_75t_L g7056 ( 
.A(n_7002),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_7021),
.Y(n_7057)
);

INVx2_ASAP7_75t_L g7058 ( 
.A(n_6956),
.Y(n_7058)
);

OR2x2_ASAP7_75t_L g7059 ( 
.A(n_7001),
.B(n_6741),
.Y(n_7059)
);

AO21x2_ASAP7_75t_L g7060 ( 
.A1(n_6973),
.A2(n_6844),
.B(n_6821),
.Y(n_7060)
);

INVx1_ASAP7_75t_L g7061 ( 
.A(n_7021),
.Y(n_7061)
);

NAND2xp5_ASAP7_75t_L g7062 ( 
.A(n_6893),
.B(n_6865),
.Y(n_7062)
);

INVxp67_ASAP7_75t_SL g7063 ( 
.A(n_6921),
.Y(n_7063)
);

INVx1_ASAP7_75t_L g7064 ( 
.A(n_6973),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_6991),
.Y(n_7065)
);

INVx2_ASAP7_75t_SL g7066 ( 
.A(n_6990),
.Y(n_7066)
);

NAND2xp5_ASAP7_75t_L g7067 ( 
.A(n_6925),
.B(n_6854),
.Y(n_7067)
);

INVx1_ASAP7_75t_L g7068 ( 
.A(n_6907),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_6912),
.Y(n_7069)
);

AND2x2_ASAP7_75t_L g7070 ( 
.A(n_6936),
.B(n_6860),
.Y(n_7070)
);

INVx3_ASAP7_75t_L g7071 ( 
.A(n_7010),
.Y(n_7071)
);

BUFx2_ASAP7_75t_L g7072 ( 
.A(n_6953),
.Y(n_7072)
);

INVx2_ASAP7_75t_L g7073 ( 
.A(n_6919),
.Y(n_7073)
);

HB1xp67_ASAP7_75t_L g7074 ( 
.A(n_6953),
.Y(n_7074)
);

OR2x2_ASAP7_75t_L g7075 ( 
.A(n_7001),
.B(n_6814),
.Y(n_7075)
);

NOR2xp33_ASAP7_75t_SL g7076 ( 
.A(n_6955),
.B(n_6890),
.Y(n_7076)
);

AND2x2_ASAP7_75t_L g7077 ( 
.A(n_6915),
.B(n_6815),
.Y(n_7077)
);

AND2x2_ASAP7_75t_L g7078 ( 
.A(n_6928),
.B(n_6743),
.Y(n_7078)
);

INVx1_ASAP7_75t_L g7079 ( 
.A(n_6914),
.Y(n_7079)
);

OR2x2_ASAP7_75t_L g7080 ( 
.A(n_6972),
.B(n_6850),
.Y(n_7080)
);

AND2x2_ASAP7_75t_L g7081 ( 
.A(n_6930),
.B(n_6745),
.Y(n_7081)
);

INVxp67_ASAP7_75t_L g7082 ( 
.A(n_6902),
.Y(n_7082)
);

OR2x2_ASAP7_75t_L g7083 ( 
.A(n_7007),
.B(n_6734),
.Y(n_7083)
);

AND2x2_ASAP7_75t_L g7084 ( 
.A(n_7017),
.B(n_6877),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_6918),
.Y(n_7085)
);

BUFx3_ASAP7_75t_L g7086 ( 
.A(n_6967),
.Y(n_7086)
);

INVxp67_ASAP7_75t_L g7087 ( 
.A(n_6939),
.Y(n_7087)
);

INVx2_ASAP7_75t_L g7088 ( 
.A(n_6951),
.Y(n_7088)
);

INVx2_ASAP7_75t_SL g7089 ( 
.A(n_6960),
.Y(n_7089)
);

INVx2_ASAP7_75t_L g7090 ( 
.A(n_6993),
.Y(n_7090)
);

HB1xp67_ASAP7_75t_L g7091 ( 
.A(n_6917),
.Y(n_7091)
);

INVx2_ASAP7_75t_SL g7092 ( 
.A(n_6968),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6922),
.Y(n_7093)
);

AND2x2_ASAP7_75t_L g7094 ( 
.A(n_6952),
.B(n_6862),
.Y(n_7094)
);

HB1xp67_ASAP7_75t_L g7095 ( 
.A(n_6931),
.Y(n_7095)
);

BUFx2_ASAP7_75t_L g7096 ( 
.A(n_6993),
.Y(n_7096)
);

BUFx2_ASAP7_75t_L g7097 ( 
.A(n_6993),
.Y(n_7097)
);

INVx2_ASAP7_75t_L g7098 ( 
.A(n_6959),
.Y(n_7098)
);

NAND2xp5_ASAP7_75t_L g7099 ( 
.A(n_6925),
.B(n_6868),
.Y(n_7099)
);

OR2x2_ASAP7_75t_L g7100 ( 
.A(n_7007),
.B(n_6737),
.Y(n_7100)
);

OR2x2_ASAP7_75t_L g7101 ( 
.A(n_6920),
.B(n_6737),
.Y(n_7101)
);

HB1xp67_ASAP7_75t_L g7102 ( 
.A(n_6933),
.Y(n_7102)
);

INVx1_ASAP7_75t_L g7103 ( 
.A(n_6935),
.Y(n_7103)
);

AND2x2_ASAP7_75t_L g7104 ( 
.A(n_6940),
.B(n_6868),
.Y(n_7104)
);

OR2x2_ASAP7_75t_L g7105 ( 
.A(n_6978),
.B(n_6750),
.Y(n_7105)
);

BUFx3_ASAP7_75t_L g7106 ( 
.A(n_6940),
.Y(n_7106)
);

INVxp67_ASAP7_75t_L g7107 ( 
.A(n_6897),
.Y(n_7107)
);

NAND2xp5_ASAP7_75t_L g7108 ( 
.A(n_6923),
.B(n_6795),
.Y(n_7108)
);

INVx3_ASAP7_75t_SL g7109 ( 
.A(n_7024),
.Y(n_7109)
);

AND2x2_ASAP7_75t_L g7110 ( 
.A(n_6975),
.B(n_6755),
.Y(n_7110)
);

AND2x2_ASAP7_75t_L g7111 ( 
.A(n_6913),
.B(n_6778),
.Y(n_7111)
);

AND2x2_ASAP7_75t_L g7112 ( 
.A(n_6932),
.B(n_6780),
.Y(n_7112)
);

INVx3_ASAP7_75t_L g7113 ( 
.A(n_6988),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_6938),
.Y(n_7114)
);

AND2x2_ASAP7_75t_L g7115 ( 
.A(n_6909),
.B(n_6781),
.Y(n_7115)
);

INVxp67_ASAP7_75t_SL g7116 ( 
.A(n_7003),
.Y(n_7116)
);

AND2x2_ASAP7_75t_L g7117 ( 
.A(n_6906),
.B(n_6782),
.Y(n_7117)
);

AND2x2_ASAP7_75t_L g7118 ( 
.A(n_6954),
.B(n_6788),
.Y(n_7118)
);

INVx1_ASAP7_75t_L g7119 ( 
.A(n_6966),
.Y(n_7119)
);

HB1xp67_ASAP7_75t_L g7120 ( 
.A(n_7018),
.Y(n_7120)
);

AND2x4_ASAP7_75t_L g7121 ( 
.A(n_6970),
.B(n_6844),
.Y(n_7121)
);

AND2x4_ASAP7_75t_L g7122 ( 
.A(n_6974),
.B(n_6979),
.Y(n_7122)
);

AND2x2_ASAP7_75t_L g7123 ( 
.A(n_6969),
.B(n_6826),
.Y(n_7123)
);

BUFx6f_ASAP7_75t_L g7124 ( 
.A(n_7022),
.Y(n_7124)
);

INVx1_ASAP7_75t_L g7125 ( 
.A(n_6980),
.Y(n_7125)
);

INVx2_ASAP7_75t_L g7126 ( 
.A(n_6961),
.Y(n_7126)
);

AND2x2_ASAP7_75t_L g7127 ( 
.A(n_6962),
.B(n_6789),
.Y(n_7127)
);

INVx1_ASAP7_75t_L g7128 ( 
.A(n_6947),
.Y(n_7128)
);

BUFx6f_ASAP7_75t_L g7129 ( 
.A(n_7013),
.Y(n_7129)
);

AND2x2_ASAP7_75t_L g7130 ( 
.A(n_6901),
.B(n_6777),
.Y(n_7130)
);

NAND2xp5_ASAP7_75t_L g7131 ( 
.A(n_6916),
.B(n_6896),
.Y(n_7131)
);

BUFx2_ASAP7_75t_L g7132 ( 
.A(n_6989),
.Y(n_7132)
);

INVx3_ASAP7_75t_L g7133 ( 
.A(n_6948),
.Y(n_7133)
);

INVx1_ASAP7_75t_SL g7134 ( 
.A(n_6958),
.Y(n_7134)
);

BUFx2_ASAP7_75t_L g7135 ( 
.A(n_6977),
.Y(n_7135)
);

INVx1_ASAP7_75t_L g7136 ( 
.A(n_6949),
.Y(n_7136)
);

NAND2x1_ASAP7_75t_L g7137 ( 
.A(n_6977),
.B(n_6830),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_6950),
.Y(n_7138)
);

NOR2xp33_ASAP7_75t_L g7139 ( 
.A(n_6997),
.B(n_6835),
.Y(n_7139)
);

INVx2_ASAP7_75t_L g7140 ( 
.A(n_6976),
.Y(n_7140)
);

OR2x2_ASAP7_75t_L g7141 ( 
.A(n_6997),
.B(n_6750),
.Y(n_7141)
);

HB1xp67_ASAP7_75t_L g7142 ( 
.A(n_6964),
.Y(n_7142)
);

INVx1_ASAP7_75t_L g7143 ( 
.A(n_6985),
.Y(n_7143)
);

AND2x4_ASAP7_75t_L g7144 ( 
.A(n_7000),
.B(n_6760),
.Y(n_7144)
);

INVx1_ASAP7_75t_SL g7145 ( 
.A(n_6895),
.Y(n_7145)
);

HB1xp67_ASAP7_75t_L g7146 ( 
.A(n_6964),
.Y(n_7146)
);

HB1xp67_ASAP7_75t_L g7147 ( 
.A(n_6927),
.Y(n_7147)
);

INVx1_ASAP7_75t_L g7148 ( 
.A(n_6995),
.Y(n_7148)
);

INVxp67_ASAP7_75t_L g7149 ( 
.A(n_7013),
.Y(n_7149)
);

OR2x2_ASAP7_75t_L g7150 ( 
.A(n_7134),
.B(n_6982),
.Y(n_7150)
);

AND2x2_ASAP7_75t_L g7151 ( 
.A(n_7110),
.B(n_6929),
.Y(n_7151)
);

INVx1_ASAP7_75t_L g7152 ( 
.A(n_7054),
.Y(n_7152)
);

BUFx2_ASAP7_75t_L g7153 ( 
.A(n_7106),
.Y(n_7153)
);

INVxp67_ASAP7_75t_SL g7154 ( 
.A(n_7054),
.Y(n_7154)
);

INVx2_ASAP7_75t_L g7155 ( 
.A(n_7096),
.Y(n_7155)
);

AND2x2_ASAP7_75t_L g7156 ( 
.A(n_7035),
.B(n_6963),
.Y(n_7156)
);

AND2x2_ASAP7_75t_L g7157 ( 
.A(n_7051),
.B(n_6996),
.Y(n_7157)
);

AND2x4_ASAP7_75t_L g7158 ( 
.A(n_7033),
.B(n_7009),
.Y(n_7158)
);

OAI22xp5_ASAP7_75t_L g7159 ( 
.A1(n_7053),
.A2(n_6944),
.B1(n_6891),
.B2(n_6984),
.Y(n_7159)
);

INVx2_ASAP7_75t_L g7160 ( 
.A(n_7097),
.Y(n_7160)
);

INVx2_ASAP7_75t_L g7161 ( 
.A(n_7044),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_7056),
.Y(n_7162)
);

INVx2_ASAP7_75t_SL g7163 ( 
.A(n_7033),
.Y(n_7163)
);

INVx1_ASAP7_75t_L g7164 ( 
.A(n_7056),
.Y(n_7164)
);

AND2x2_ASAP7_75t_L g7165 ( 
.A(n_7026),
.B(n_6965),
.Y(n_7165)
);

NOR2xp67_ASAP7_75t_L g7166 ( 
.A(n_7036),
.B(n_6842),
.Y(n_7166)
);

NAND2xp5_ASAP7_75t_L g7167 ( 
.A(n_7082),
.B(n_7091),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_7036),
.Y(n_7168)
);

NOR2x1_ASAP7_75t_SL g7169 ( 
.A(n_7060),
.B(n_6803),
.Y(n_7169)
);

INVx2_ASAP7_75t_L g7170 ( 
.A(n_7044),
.Y(n_7170)
);

INVx1_ASAP7_75t_L g7171 ( 
.A(n_7095),
.Y(n_7171)
);

AND2x2_ASAP7_75t_L g7172 ( 
.A(n_7026),
.B(n_7005),
.Y(n_7172)
);

OR2x2_ASAP7_75t_L g7173 ( 
.A(n_7080),
.B(n_6992),
.Y(n_7173)
);

AND2x2_ASAP7_75t_L g7174 ( 
.A(n_7104),
.B(n_6981),
.Y(n_7174)
);

NOR2xp33_ASAP7_75t_L g7175 ( 
.A(n_7082),
.B(n_7107),
.Y(n_7175)
);

NOR2xp33_ASAP7_75t_L g7176 ( 
.A(n_7107),
.B(n_6905),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_7095),
.Y(n_7177)
);

INVx1_ASAP7_75t_L g7178 ( 
.A(n_7102),
.Y(n_7178)
);

INVx1_ASAP7_75t_L g7179 ( 
.A(n_7102),
.Y(n_7179)
);

INVx1_ASAP7_75t_L g7180 ( 
.A(n_7074),
.Y(n_7180)
);

OR2x2_ASAP7_75t_L g7181 ( 
.A(n_7145),
.B(n_6987),
.Y(n_7181)
);

INVx1_ASAP7_75t_L g7182 ( 
.A(n_7074),
.Y(n_7182)
);

INVx2_ASAP7_75t_L g7183 ( 
.A(n_7044),
.Y(n_7183)
);

OR2x2_ASAP7_75t_L g7184 ( 
.A(n_7145),
.B(n_6987),
.Y(n_7184)
);

INVx1_ASAP7_75t_L g7185 ( 
.A(n_7072),
.Y(n_7185)
);

AND2x2_ASAP7_75t_L g7186 ( 
.A(n_7094),
.B(n_6981),
.Y(n_7186)
);

HB1xp67_ASAP7_75t_L g7187 ( 
.A(n_7060),
.Y(n_7187)
);

NOR2x1_ASAP7_75t_L g7188 ( 
.A(n_7040),
.B(n_6835),
.Y(n_7188)
);

NOR2x1_ASAP7_75t_L g7189 ( 
.A(n_7043),
.B(n_6891),
.Y(n_7189)
);

INVx1_ASAP7_75t_L g7190 ( 
.A(n_7050),
.Y(n_7190)
);

AND2x2_ASAP7_75t_L g7191 ( 
.A(n_7031),
.B(n_6983),
.Y(n_7191)
);

AND2x4_ASAP7_75t_L g7192 ( 
.A(n_7111),
.B(n_7011),
.Y(n_7192)
);

NOR2x1_ASAP7_75t_L g7193 ( 
.A(n_7064),
.B(n_6905),
.Y(n_7193)
);

NAND2xp5_ASAP7_75t_L g7194 ( 
.A(n_7091),
.B(n_7003),
.Y(n_7194)
);

INVx2_ASAP7_75t_L g7195 ( 
.A(n_7137),
.Y(n_7195)
);

INVx2_ASAP7_75t_L g7196 ( 
.A(n_7071),
.Y(n_7196)
);

INVx1_ASAP7_75t_L g7197 ( 
.A(n_7057),
.Y(n_7197)
);

AND2x2_ASAP7_75t_L g7198 ( 
.A(n_7132),
.B(n_7006),
.Y(n_7198)
);

AND2x2_ASAP7_75t_L g7199 ( 
.A(n_7115),
.B(n_7117),
.Y(n_7199)
);

NAND2xp5_ASAP7_75t_L g7200 ( 
.A(n_7131),
.B(n_6916),
.Y(n_7200)
);

OR2x2_ASAP7_75t_L g7201 ( 
.A(n_7135),
.B(n_6999),
.Y(n_7201)
);

OAI21xp5_ASAP7_75t_SL g7202 ( 
.A1(n_7053),
.A2(n_6984),
.B(n_6986),
.Y(n_7202)
);

INVx2_ASAP7_75t_L g7203 ( 
.A(n_7071),
.Y(n_7203)
);

INVx4_ASAP7_75t_L g7204 ( 
.A(n_7039),
.Y(n_7204)
);

AND2x2_ASAP7_75t_L g7205 ( 
.A(n_7127),
.B(n_6863),
.Y(n_7205)
);

INVxp33_ASAP7_75t_SL g7206 ( 
.A(n_7147),
.Y(n_7206)
);

NAND2xp5_ASAP7_75t_L g7207 ( 
.A(n_7131),
.B(n_7023),
.Y(n_7207)
);

INVxp67_ASAP7_75t_L g7208 ( 
.A(n_7147),
.Y(n_7208)
);

AND2x2_ASAP7_75t_L g7209 ( 
.A(n_7112),
.B(n_6863),
.Y(n_7209)
);

CKINVDCx16_ASAP7_75t_R g7210 ( 
.A(n_7076),
.Y(n_7210)
);

AND2x2_ASAP7_75t_L g7211 ( 
.A(n_7027),
.B(n_6859),
.Y(n_7211)
);

INVx1_ASAP7_75t_L g7212 ( 
.A(n_7061),
.Y(n_7212)
);

INVx1_ASAP7_75t_L g7213 ( 
.A(n_7037),
.Y(n_7213)
);

INVx2_ASAP7_75t_L g7214 ( 
.A(n_7090),
.Y(n_7214)
);

OR2x6_ASAP7_75t_L g7215 ( 
.A(n_7037),
.B(n_6986),
.Y(n_7215)
);

NOR3xp33_ASAP7_75t_L g7216 ( 
.A(n_7041),
.B(n_6999),
.C(n_7004),
.Y(n_7216)
);

INVx1_ASAP7_75t_L g7217 ( 
.A(n_7025),
.Y(n_7217)
);

INVx1_ASAP7_75t_L g7218 ( 
.A(n_7029),
.Y(n_7218)
);

AND2x2_ASAP7_75t_L g7219 ( 
.A(n_7087),
.B(n_6861),
.Y(n_7219)
);

NAND2xp5_ASAP7_75t_L g7220 ( 
.A(n_7116),
.B(n_7063),
.Y(n_7220)
);

NAND2xp5_ASAP7_75t_L g7221 ( 
.A(n_7070),
.B(n_7008),
.Y(n_7221)
);

AND2x2_ASAP7_75t_L g7222 ( 
.A(n_7087),
.B(n_6856),
.Y(n_7222)
);

NAND2xp5_ASAP7_75t_L g7223 ( 
.A(n_7049),
.B(n_7120),
.Y(n_7223)
);

AND2x2_ASAP7_75t_L g7224 ( 
.A(n_7130),
.B(n_6760),
.Y(n_7224)
);

AND2x2_ASAP7_75t_L g7225 ( 
.A(n_7118),
.B(n_6821),
.Y(n_7225)
);

AND2x4_ASAP7_75t_L g7226 ( 
.A(n_7052),
.B(n_7012),
.Y(n_7226)
);

NAND2xp5_ASAP7_75t_L g7227 ( 
.A(n_7116),
.B(n_7014),
.Y(n_7227)
);

INVx1_ASAP7_75t_L g7228 ( 
.A(n_7038),
.Y(n_7228)
);

NOR3xp33_ASAP7_75t_L g7229 ( 
.A(n_7041),
.B(n_6812),
.C(n_7015),
.Y(n_7229)
);

INVx3_ASAP7_75t_L g7230 ( 
.A(n_7113),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_7045),
.Y(n_7231)
);

AND2x2_ASAP7_75t_L g7232 ( 
.A(n_7081),
.B(n_6833),
.Y(n_7232)
);

AND2x2_ASAP7_75t_L g7233 ( 
.A(n_7073),
.B(n_6833),
.Y(n_7233)
);

AND2x2_ASAP7_75t_L g7234 ( 
.A(n_7078),
.B(n_7019),
.Y(n_7234)
);

NAND2xp5_ASAP7_75t_L g7235 ( 
.A(n_7123),
.B(n_6806),
.Y(n_7235)
);

AND2x2_ASAP7_75t_L g7236 ( 
.A(n_7109),
.B(n_6802),
.Y(n_7236)
);

NAND2xp5_ASAP7_75t_L g7237 ( 
.A(n_7063),
.B(n_6808),
.Y(n_7237)
);

NAND2xp5_ASAP7_75t_L g7238 ( 
.A(n_7142),
.B(n_6811),
.Y(n_7238)
);

AND2x2_ASAP7_75t_L g7239 ( 
.A(n_7126),
.B(n_6816),
.Y(n_7239)
);

AND2x2_ASAP7_75t_L g7240 ( 
.A(n_7084),
.B(n_6817),
.Y(n_7240)
);

INVxp67_ASAP7_75t_L g7241 ( 
.A(n_7076),
.Y(n_7241)
);

INVx2_ASAP7_75t_L g7242 ( 
.A(n_7086),
.Y(n_7242)
);

NAND2xp5_ASAP7_75t_SL g7243 ( 
.A(n_7129),
.B(n_6971),
.Y(n_7243)
);

OR2x2_ASAP7_75t_L g7244 ( 
.A(n_7028),
.B(n_6813),
.Y(n_7244)
);

INVx1_ASAP7_75t_L g7245 ( 
.A(n_7065),
.Y(n_7245)
);

OR2x2_ASAP7_75t_L g7246 ( 
.A(n_7030),
.B(n_6819),
.Y(n_7246)
);

INVx1_ASAP7_75t_L g7247 ( 
.A(n_7075),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_L g7248 ( 
.A(n_7142),
.B(n_6820),
.Y(n_7248)
);

INVx1_ASAP7_75t_L g7249 ( 
.A(n_7113),
.Y(n_7249)
);

INVx2_ASAP7_75t_L g7250 ( 
.A(n_7032),
.Y(n_7250)
);

NAND2xp5_ASAP7_75t_L g7251 ( 
.A(n_7146),
.B(n_6825),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_7133),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_7133),
.Y(n_7253)
);

NAND2xp5_ASAP7_75t_L g7254 ( 
.A(n_7144),
.B(n_6836),
.Y(n_7254)
);

OR2x2_ASAP7_75t_L g7255 ( 
.A(n_7034),
.B(n_7048),
.Y(n_7255)
);

AND2x2_ASAP7_75t_L g7256 ( 
.A(n_7042),
.B(n_6839),
.Y(n_7256)
);

NAND2xp5_ASAP7_75t_L g7257 ( 
.A(n_7144),
.B(n_6838),
.Y(n_7257)
);

NAND2xp5_ASAP7_75t_SL g7258 ( 
.A(n_7129),
.B(n_6831),
.Y(n_7258)
);

AND2x2_ASAP7_75t_L g7259 ( 
.A(n_7151),
.B(n_7066),
.Y(n_7259)
);

AND2x2_ASAP7_75t_L g7260 ( 
.A(n_7186),
.B(n_7058),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_7187),
.Y(n_7261)
);

OR2x2_ASAP7_75t_L g7262 ( 
.A(n_7210),
.B(n_7099),
.Y(n_7262)
);

OAI22xp5_ASAP7_75t_L g7263 ( 
.A1(n_7193),
.A2(n_7055),
.B1(n_7108),
.B2(n_7105),
.Y(n_7263)
);

INVx2_ASAP7_75t_L g7264 ( 
.A(n_7163),
.Y(n_7264)
);

INVx1_ASAP7_75t_L g7265 ( 
.A(n_7166),
.Y(n_7265)
);

AND2x2_ASAP7_75t_L g7266 ( 
.A(n_7199),
.B(n_7098),
.Y(n_7266)
);

INVx1_ASAP7_75t_L g7267 ( 
.A(n_7166),
.Y(n_7267)
);

NAND2xp5_ASAP7_75t_L g7268 ( 
.A(n_7193),
.B(n_7202),
.Y(n_7268)
);

NAND2xp5_ASAP7_75t_L g7269 ( 
.A(n_7202),
.B(n_7089),
.Y(n_7269)
);

AND2x2_ASAP7_75t_L g7270 ( 
.A(n_7174),
.B(n_7077),
.Y(n_7270)
);

NAND2xp5_ASAP7_75t_L g7271 ( 
.A(n_7154),
.B(n_7092),
.Y(n_7271)
);

AND2x2_ASAP7_75t_L g7272 ( 
.A(n_7156),
.B(n_7140),
.Y(n_7272)
);

NOR2xp67_ASAP7_75t_L g7273 ( 
.A(n_7208),
.B(n_7059),
.Y(n_7273)
);

INVx2_ASAP7_75t_L g7274 ( 
.A(n_7230),
.Y(n_7274)
);

HB1xp67_ASAP7_75t_L g7275 ( 
.A(n_7215),
.Y(n_7275)
);

INVx1_ASAP7_75t_L g7276 ( 
.A(n_7152),
.Y(n_7276)
);

BUFx3_ASAP7_75t_L g7277 ( 
.A(n_7153),
.Y(n_7277)
);

AND2x2_ASAP7_75t_L g7278 ( 
.A(n_7209),
.B(n_7088),
.Y(n_7278)
);

INVx1_ASAP7_75t_L g7279 ( 
.A(n_7162),
.Y(n_7279)
);

AND2x2_ASAP7_75t_L g7280 ( 
.A(n_7157),
.B(n_7124),
.Y(n_7280)
);

INVx1_ASAP7_75t_L g7281 ( 
.A(n_7164),
.Y(n_7281)
);

NOR4xp25_ASAP7_75t_SL g7282 ( 
.A(n_7243),
.B(n_7069),
.C(n_7079),
.D(n_7068),
.Y(n_7282)
);

AND2x2_ASAP7_75t_L g7283 ( 
.A(n_7224),
.B(n_7124),
.Y(n_7283)
);

AND2x2_ASAP7_75t_L g7284 ( 
.A(n_7165),
.B(n_7225),
.Y(n_7284)
);

AND2x2_ASAP7_75t_L g7285 ( 
.A(n_7236),
.B(n_7124),
.Y(n_7285)
);

AND2x2_ASAP7_75t_L g7286 ( 
.A(n_7205),
.B(n_7129),
.Y(n_7286)
);

AND2x2_ASAP7_75t_L g7287 ( 
.A(n_7232),
.B(n_7121),
.Y(n_7287)
);

AND2x2_ASAP7_75t_L g7288 ( 
.A(n_7198),
.B(n_7121),
.Y(n_7288)
);

INVx1_ASAP7_75t_L g7289 ( 
.A(n_7168),
.Y(n_7289)
);

NOR2xp33_ASAP7_75t_L g7290 ( 
.A(n_7206),
.B(n_7099),
.Y(n_7290)
);

INVx1_ASAP7_75t_L g7291 ( 
.A(n_7167),
.Y(n_7291)
);

INVx1_ASAP7_75t_L g7292 ( 
.A(n_7171),
.Y(n_7292)
);

NAND2xp5_ASAP7_75t_L g7293 ( 
.A(n_7215),
.B(n_7159),
.Y(n_7293)
);

BUFx6f_ASAP7_75t_SL g7294 ( 
.A(n_7215),
.Y(n_7294)
);

INVx1_ASAP7_75t_L g7295 ( 
.A(n_7177),
.Y(n_7295)
);

AND2x2_ASAP7_75t_L g7296 ( 
.A(n_7191),
.B(n_7101),
.Y(n_7296)
);

NAND2xp5_ASAP7_75t_L g7297 ( 
.A(n_7159),
.B(n_7122),
.Y(n_7297)
);

NOR2xp33_ASAP7_75t_L g7298 ( 
.A(n_7241),
.B(n_7083),
.Y(n_7298)
);

AND2x2_ASAP7_75t_L g7299 ( 
.A(n_7219),
.B(n_7149),
.Y(n_7299)
);

OR2x2_ASAP7_75t_L g7300 ( 
.A(n_7150),
.B(n_7100),
.Y(n_7300)
);

NAND2xp5_ASAP7_75t_L g7301 ( 
.A(n_7176),
.B(n_7122),
.Y(n_7301)
);

AND2x2_ASAP7_75t_L g7302 ( 
.A(n_7222),
.B(n_7149),
.Y(n_7302)
);

INVx1_ASAP7_75t_L g7303 ( 
.A(n_7178),
.Y(n_7303)
);

NAND2xp5_ASAP7_75t_L g7304 ( 
.A(n_7189),
.B(n_7046),
.Y(n_7304)
);

BUFx2_ASAP7_75t_L g7305 ( 
.A(n_7158),
.Y(n_7305)
);

AOI22xp5_ASAP7_75t_L g7306 ( 
.A1(n_7216),
.A2(n_7108),
.B1(n_7055),
.B2(n_7139),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_7179),
.Y(n_7307)
);

AND2x2_ASAP7_75t_L g7308 ( 
.A(n_7211),
.B(n_7047),
.Y(n_7308)
);

INVx2_ASAP7_75t_L g7309 ( 
.A(n_7230),
.Y(n_7309)
);

AND2x2_ASAP7_75t_L g7310 ( 
.A(n_7172),
.B(n_7141),
.Y(n_7310)
);

INVx1_ASAP7_75t_L g7311 ( 
.A(n_7180),
.Y(n_7311)
);

INVx1_ASAP7_75t_L g7312 ( 
.A(n_7182),
.Y(n_7312)
);

OR2x2_ASAP7_75t_L g7313 ( 
.A(n_7173),
.B(n_7067),
.Y(n_7313)
);

INVx2_ASAP7_75t_L g7314 ( 
.A(n_7158),
.Y(n_7314)
);

OAI21xp33_ASAP7_75t_L g7315 ( 
.A1(n_7200),
.A2(n_7062),
.B(n_7119),
.Y(n_7315)
);

INVx1_ASAP7_75t_L g7316 ( 
.A(n_7223),
.Y(n_7316)
);

NAND2xp5_ASAP7_75t_L g7317 ( 
.A(n_7189),
.B(n_7085),
.Y(n_7317)
);

NOR2xp33_ASAP7_75t_L g7318 ( 
.A(n_7200),
.B(n_7062),
.Y(n_7318)
);

INVx1_ASAP7_75t_L g7319 ( 
.A(n_7257),
.Y(n_7319)
);

INVx1_ASAP7_75t_L g7320 ( 
.A(n_7257),
.Y(n_7320)
);

INVx2_ASAP7_75t_L g7321 ( 
.A(n_7169),
.Y(n_7321)
);

AND2x2_ASAP7_75t_L g7322 ( 
.A(n_7233),
.B(n_7240),
.Y(n_7322)
);

INVx2_ASAP7_75t_L g7323 ( 
.A(n_7195),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_7254),
.Y(n_7324)
);

HB1xp67_ASAP7_75t_L g7325 ( 
.A(n_7220),
.Y(n_7325)
);

INVx1_ASAP7_75t_L g7326 ( 
.A(n_7254),
.Y(n_7326)
);

INVx1_ASAP7_75t_L g7327 ( 
.A(n_7185),
.Y(n_7327)
);

INVx3_ASAP7_75t_L g7328 ( 
.A(n_7204),
.Y(n_7328)
);

NAND2xp5_ASAP7_75t_L g7329 ( 
.A(n_7175),
.B(n_7093),
.Y(n_7329)
);

BUFx6f_ASAP7_75t_L g7330 ( 
.A(n_7161),
.Y(n_7330)
);

AND2x4_ASAP7_75t_L g7331 ( 
.A(n_7170),
.B(n_7125),
.Y(n_7331)
);

INVx2_ASAP7_75t_L g7332 ( 
.A(n_7183),
.Y(n_7332)
);

AND2x2_ASAP7_75t_L g7333 ( 
.A(n_7242),
.B(n_7103),
.Y(n_7333)
);

NOR2xp33_ASAP7_75t_L g7334 ( 
.A(n_7220),
.B(n_7114),
.Y(n_7334)
);

INVx1_ASAP7_75t_L g7335 ( 
.A(n_7237),
.Y(n_7335)
);

INVx2_ASAP7_75t_SL g7336 ( 
.A(n_7192),
.Y(n_7336)
);

AND2x2_ASAP7_75t_L g7337 ( 
.A(n_7239),
.B(n_7128),
.Y(n_7337)
);

INVx1_ASAP7_75t_L g7338 ( 
.A(n_7237),
.Y(n_7338)
);

NAND3xp33_ASAP7_75t_L g7339 ( 
.A(n_7194),
.B(n_7138),
.C(n_7136),
.Y(n_7339)
);

NAND2x1p5_ASAP7_75t_L g7340 ( 
.A(n_7204),
.B(n_7143),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_7305),
.Y(n_7341)
);

INVx3_ASAP7_75t_L g7342 ( 
.A(n_7328),
.Y(n_7342)
);

HB1xp67_ASAP7_75t_L g7343 ( 
.A(n_7275),
.Y(n_7343)
);

AND2x2_ASAP7_75t_L g7344 ( 
.A(n_7284),
.B(n_7192),
.Y(n_7344)
);

AOI22xp5_ASAP7_75t_L g7345 ( 
.A1(n_7263),
.A2(n_7229),
.B1(n_7258),
.B2(n_7207),
.Y(n_7345)
);

OR2x2_ASAP7_75t_L g7346 ( 
.A(n_7336),
.B(n_7255),
.Y(n_7346)
);

NAND2xp33_ASAP7_75t_SL g7347 ( 
.A(n_7294),
.B(n_7181),
.Y(n_7347)
);

AND2x4_ASAP7_75t_L g7348 ( 
.A(n_7288),
.B(n_7196),
.Y(n_7348)
);

INVx1_ASAP7_75t_L g7349 ( 
.A(n_7275),
.Y(n_7349)
);

NAND2xp5_ASAP7_75t_L g7350 ( 
.A(n_7263),
.B(n_7268),
.Y(n_7350)
);

OR2x2_ASAP7_75t_L g7351 ( 
.A(n_7269),
.B(n_7221),
.Y(n_7351)
);

INVx1_ASAP7_75t_L g7352 ( 
.A(n_7294),
.Y(n_7352)
);

INVx1_ASAP7_75t_L g7353 ( 
.A(n_7265),
.Y(n_7353)
);

INVx1_ASAP7_75t_L g7354 ( 
.A(n_7267),
.Y(n_7354)
);

OR2x2_ASAP7_75t_L g7355 ( 
.A(n_7269),
.B(n_7201),
.Y(n_7355)
);

NOR3xp33_ASAP7_75t_L g7356 ( 
.A(n_7268),
.B(n_7247),
.C(n_7207),
.Y(n_7356)
);

AND2x2_ASAP7_75t_L g7357 ( 
.A(n_7259),
.B(n_7250),
.Y(n_7357)
);

INVx1_ASAP7_75t_L g7358 ( 
.A(n_7271),
.Y(n_7358)
);

AND2x4_ASAP7_75t_L g7359 ( 
.A(n_7277),
.B(n_7203),
.Y(n_7359)
);

OR2x2_ASAP7_75t_L g7360 ( 
.A(n_7262),
.B(n_7184),
.Y(n_7360)
);

AND2x2_ASAP7_75t_L g7361 ( 
.A(n_7283),
.B(n_7234),
.Y(n_7361)
);

AND2x2_ASAP7_75t_L g7362 ( 
.A(n_7287),
.B(n_7256),
.Y(n_7362)
);

INVxp67_ASAP7_75t_L g7363 ( 
.A(n_7290),
.Y(n_7363)
);

AND2x2_ASAP7_75t_L g7364 ( 
.A(n_7270),
.B(n_7245),
.Y(n_7364)
);

OR2x2_ASAP7_75t_L g7365 ( 
.A(n_7314),
.B(n_7235),
.Y(n_7365)
);

NOR2xp33_ASAP7_75t_L g7366 ( 
.A(n_7330),
.B(n_7244),
.Y(n_7366)
);

AND2x2_ASAP7_75t_L g7367 ( 
.A(n_7280),
.B(n_7226),
.Y(n_7367)
);

AOI211xp5_ASAP7_75t_SL g7368 ( 
.A1(n_7318),
.A2(n_7213),
.B(n_7227),
.C(n_7252),
.Y(n_7368)
);

AND2x2_ASAP7_75t_L g7369 ( 
.A(n_7260),
.B(n_7249),
.Y(n_7369)
);

NAND4xp75_ASAP7_75t_L g7370 ( 
.A(n_7273),
.B(n_7188),
.C(n_7253),
.D(n_7227),
.Y(n_7370)
);

NAND2xp5_ASAP7_75t_L g7371 ( 
.A(n_7318),
.B(n_7188),
.Y(n_7371)
);

AND2x2_ASAP7_75t_L g7372 ( 
.A(n_7272),
.B(n_7296),
.Y(n_7372)
);

INVx1_ASAP7_75t_L g7373 ( 
.A(n_7325),
.Y(n_7373)
);

BUFx2_ASAP7_75t_L g7374 ( 
.A(n_7340),
.Y(n_7374)
);

INVx2_ASAP7_75t_SL g7375 ( 
.A(n_7286),
.Y(n_7375)
);

INVx2_ASAP7_75t_L g7376 ( 
.A(n_7340),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_7310),
.Y(n_7377)
);

NAND2x1p5_ASAP7_75t_L g7378 ( 
.A(n_7285),
.B(n_7155),
.Y(n_7378)
);

AND2x4_ASAP7_75t_L g7379 ( 
.A(n_7264),
.B(n_7160),
.Y(n_7379)
);

AND2x2_ASAP7_75t_L g7380 ( 
.A(n_7322),
.B(n_7231),
.Y(n_7380)
);

AND2x4_ASAP7_75t_L g7381 ( 
.A(n_7274),
.B(n_7190),
.Y(n_7381)
);

OR2x2_ASAP7_75t_L g7382 ( 
.A(n_7297),
.B(n_7246),
.Y(n_7382)
);

INVx1_ASAP7_75t_L g7383 ( 
.A(n_7321),
.Y(n_7383)
);

OAI211xp5_ASAP7_75t_SL g7384 ( 
.A1(n_7306),
.A2(n_7248),
.B(n_7251),
.C(n_7238),
.Y(n_7384)
);

INVx1_ASAP7_75t_L g7385 ( 
.A(n_7321),
.Y(n_7385)
);

INVx1_ASAP7_75t_L g7386 ( 
.A(n_7308),
.Y(n_7386)
);

AND2x2_ASAP7_75t_L g7387 ( 
.A(n_7266),
.B(n_7197),
.Y(n_7387)
);

NAND4xp25_ASAP7_75t_L g7388 ( 
.A(n_7293),
.B(n_7212),
.C(n_7218),
.D(n_7217),
.Y(n_7388)
);

AND2x2_ASAP7_75t_L g7389 ( 
.A(n_7278),
.B(n_7228),
.Y(n_7389)
);

AND2x4_ASAP7_75t_L g7390 ( 
.A(n_7309),
.B(n_7214),
.Y(n_7390)
);

INVx1_ASAP7_75t_SL g7391 ( 
.A(n_7304),
.Y(n_7391)
);

INVx1_ASAP7_75t_L g7392 ( 
.A(n_7299),
.Y(n_7392)
);

AND2x2_ASAP7_75t_L g7393 ( 
.A(n_7302),
.B(n_7148),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_7304),
.Y(n_7394)
);

INVx1_ASAP7_75t_L g7395 ( 
.A(n_7317),
.Y(n_7395)
);

AND2x2_ASAP7_75t_L g7396 ( 
.A(n_7332),
.B(n_7238),
.Y(n_7396)
);

NAND4xp25_ASAP7_75t_L g7397 ( 
.A(n_7293),
.B(n_7251),
.C(n_7248),
.D(n_7020),
.Y(n_7397)
);

AND2x2_ASAP7_75t_L g7398 ( 
.A(n_7333),
.B(n_6800),
.Y(n_7398)
);

INVx3_ASAP7_75t_L g7399 ( 
.A(n_7330),
.Y(n_7399)
);

NAND2xp5_ASAP7_75t_L g7400 ( 
.A(n_7331),
.B(n_6840),
.Y(n_7400)
);

OAI33xp33_ASAP7_75t_L g7401 ( 
.A1(n_7297),
.A2(n_6807),
.A3(n_6886),
.B1(n_6827),
.B2(n_6873),
.B3(n_6803),
.Y(n_7401)
);

INVx1_ASAP7_75t_L g7402 ( 
.A(n_7317),
.Y(n_7402)
);

BUFx3_ASAP7_75t_L g7403 ( 
.A(n_7323),
.Y(n_7403)
);

AND2x2_ASAP7_75t_L g7404 ( 
.A(n_7337),
.B(n_6759),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_7261),
.Y(n_7405)
);

INVx1_ASAP7_75t_SL g7406 ( 
.A(n_7300),
.Y(n_7406)
);

OAI22xp5_ASAP7_75t_L g7407 ( 
.A1(n_7345),
.A2(n_7313),
.B1(n_7301),
.B2(n_7282),
.Y(n_7407)
);

OAI322xp33_ASAP7_75t_L g7408 ( 
.A1(n_7345),
.A2(n_7334),
.A3(n_7301),
.B1(n_7329),
.B2(n_7338),
.C1(n_7335),
.C2(n_7298),
.Y(n_7408)
);

OAI22xp33_ASAP7_75t_SL g7409 ( 
.A1(n_7350),
.A2(n_7276),
.B1(n_7281),
.B2(n_7279),
.Y(n_7409)
);

AOI21x1_ASAP7_75t_L g7410 ( 
.A1(n_7350),
.A2(n_7289),
.B(n_7329),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_7346),
.Y(n_7411)
);

INVxp67_ASAP7_75t_L g7412 ( 
.A(n_7374),
.Y(n_7412)
);

OAI322xp33_ASAP7_75t_L g7413 ( 
.A1(n_7371),
.A2(n_7334),
.A3(n_7298),
.B1(n_7312),
.B2(n_7311),
.C1(n_7327),
.C2(n_7339),
.Y(n_7413)
);

AND2x2_ASAP7_75t_L g7414 ( 
.A(n_7372),
.B(n_7316),
.Y(n_7414)
);

NAND2xp5_ASAP7_75t_L g7415 ( 
.A(n_7344),
.B(n_7331),
.Y(n_7415)
);

OAI32xp33_ASAP7_75t_L g7416 ( 
.A1(n_7371),
.A2(n_7315),
.A3(n_7339),
.B1(n_7303),
.B2(n_7307),
.Y(n_7416)
);

INVx2_ASAP7_75t_L g7417 ( 
.A(n_7399),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_7343),
.Y(n_7418)
);

INVx1_ASAP7_75t_L g7419 ( 
.A(n_7399),
.Y(n_7419)
);

AOI22xp5_ASAP7_75t_L g7420 ( 
.A1(n_7375),
.A2(n_7291),
.B1(n_7295),
.B2(n_7292),
.Y(n_7420)
);

INVx1_ASAP7_75t_SL g7421 ( 
.A(n_7406),
.Y(n_7421)
);

AOI221xp5_ASAP7_75t_L g7422 ( 
.A1(n_7356),
.A2(n_7326),
.B1(n_7324),
.B2(n_7319),
.C(n_7320),
.Y(n_7422)
);

OR2x2_ASAP7_75t_L g7423 ( 
.A(n_7341),
.B(n_7282),
.Y(n_7423)
);

INVx1_ASAP7_75t_SL g7424 ( 
.A(n_7367),
.Y(n_7424)
);

INVx3_ASAP7_75t_L g7425 ( 
.A(n_7342),
.Y(n_7425)
);

INVx1_ASAP7_75t_L g7426 ( 
.A(n_7342),
.Y(n_7426)
);

OR2x2_ASAP7_75t_L g7427 ( 
.A(n_7360),
.B(n_308),
.Y(n_7427)
);

OAI33xp33_ASAP7_75t_L g7428 ( 
.A1(n_7384),
.A2(n_313),
.A3(n_317),
.B1(n_311),
.B2(n_312),
.B3(n_315),
.Y(n_7428)
);

INVx1_ASAP7_75t_L g7429 ( 
.A(n_7380),
.Y(n_7429)
);

NAND3xp33_ASAP7_75t_L g7430 ( 
.A(n_7368),
.B(n_313),
.C(n_315),
.Y(n_7430)
);

INVx2_ASAP7_75t_L g7431 ( 
.A(n_7378),
.Y(n_7431)
);

OR2x2_ASAP7_75t_L g7432 ( 
.A(n_7382),
.B(n_317),
.Y(n_7432)
);

INVx1_ASAP7_75t_L g7433 ( 
.A(n_7359),
.Y(n_7433)
);

AND2x2_ASAP7_75t_L g7434 ( 
.A(n_7361),
.B(n_318),
.Y(n_7434)
);

OAI32xp33_ASAP7_75t_L g7435 ( 
.A1(n_7391),
.A2(n_324),
.A3(n_319),
.B1(n_322),
.B2(n_325),
.Y(n_7435)
);

INVx1_ASAP7_75t_L g7436 ( 
.A(n_7359),
.Y(n_7436)
);

OR2x2_ASAP7_75t_L g7437 ( 
.A(n_7355),
.B(n_325),
.Y(n_7437)
);

INVx1_ASAP7_75t_L g7438 ( 
.A(n_7364),
.Y(n_7438)
);

INVx2_ASAP7_75t_L g7439 ( 
.A(n_7348),
.Y(n_7439)
);

INVx1_ASAP7_75t_L g7440 ( 
.A(n_7370),
.Y(n_7440)
);

NAND2xp5_ASAP7_75t_L g7441 ( 
.A(n_7362),
.B(n_326),
.Y(n_7441)
);

INVxp67_ASAP7_75t_L g7442 ( 
.A(n_7366),
.Y(n_7442)
);

OR2x2_ASAP7_75t_L g7443 ( 
.A(n_7377),
.B(n_327),
.Y(n_7443)
);

NAND2x1p5_ASAP7_75t_L g7444 ( 
.A(n_7357),
.B(n_328),
.Y(n_7444)
);

NAND2x1_ASAP7_75t_L g7445 ( 
.A(n_7373),
.B(n_329),
.Y(n_7445)
);

OR2x2_ASAP7_75t_L g7446 ( 
.A(n_7351),
.B(n_329),
.Y(n_7446)
);

AND2x2_ASAP7_75t_L g7447 ( 
.A(n_7369),
.B(n_330),
.Y(n_7447)
);

INVx2_ASAP7_75t_SL g7448 ( 
.A(n_7376),
.Y(n_7448)
);

NAND2x1p5_ASAP7_75t_L g7449 ( 
.A(n_7379),
.B(n_7403),
.Y(n_7449)
);

INVx2_ASAP7_75t_L g7450 ( 
.A(n_7379),
.Y(n_7450)
);

OAI31xp33_ASAP7_75t_L g7451 ( 
.A1(n_7384),
.A2(n_335),
.A3(n_330),
.B(n_331),
.Y(n_7451)
);

AOI22xp5_ASAP7_75t_L g7452 ( 
.A1(n_7363),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_7452)
);

NAND2xp5_ASAP7_75t_L g7453 ( 
.A(n_7349),
.B(n_336),
.Y(n_7453)
);

OR2x2_ASAP7_75t_L g7454 ( 
.A(n_7365),
.B(n_339),
.Y(n_7454)
);

INVx1_ASAP7_75t_L g7455 ( 
.A(n_7387),
.Y(n_7455)
);

OR2x2_ASAP7_75t_L g7456 ( 
.A(n_7386),
.B(n_339),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_7389),
.Y(n_7457)
);

NAND2xp5_ASAP7_75t_L g7458 ( 
.A(n_7398),
.B(n_7368),
.Y(n_7458)
);

NOR2xp33_ASAP7_75t_L g7459 ( 
.A(n_7392),
.B(n_340),
.Y(n_7459)
);

OAI33xp33_ASAP7_75t_L g7460 ( 
.A1(n_7383),
.A2(n_341),
.A3(n_343),
.B1(n_344),
.B2(n_345),
.B3(n_346),
.Y(n_7460)
);

NAND3xp33_ASAP7_75t_L g7461 ( 
.A(n_7347),
.B(n_343),
.C(n_345),
.Y(n_7461)
);

INVx1_ASAP7_75t_L g7462 ( 
.A(n_7449),
.Y(n_7462)
);

INVxp67_ASAP7_75t_L g7463 ( 
.A(n_7415),
.Y(n_7463)
);

INVx2_ASAP7_75t_L g7464 ( 
.A(n_7425),
.Y(n_7464)
);

INVx1_ASAP7_75t_L g7465 ( 
.A(n_7425),
.Y(n_7465)
);

NAND2xp5_ASAP7_75t_L g7466 ( 
.A(n_7424),
.B(n_7391),
.Y(n_7466)
);

NAND2xp5_ASAP7_75t_L g7467 ( 
.A(n_7421),
.B(n_7390),
.Y(n_7467)
);

NAND2xp5_ASAP7_75t_L g7468 ( 
.A(n_7433),
.B(n_7390),
.Y(n_7468)
);

INVx3_ASAP7_75t_L g7469 ( 
.A(n_7450),
.Y(n_7469)
);

NOR2x1_ASAP7_75t_L g7470 ( 
.A(n_7430),
.B(n_7388),
.Y(n_7470)
);

CKINVDCx5p33_ASAP7_75t_R g7471 ( 
.A(n_7431),
.Y(n_7471)
);

INVx3_ASAP7_75t_L g7472 ( 
.A(n_7439),
.Y(n_7472)
);

AND3x1_ASAP7_75t_L g7473 ( 
.A(n_7451),
.B(n_7396),
.C(n_7352),
.Y(n_7473)
);

INVx1_ASAP7_75t_L g7474 ( 
.A(n_7436),
.Y(n_7474)
);

INVx1_ASAP7_75t_L g7475 ( 
.A(n_7444),
.Y(n_7475)
);

NAND2xp5_ASAP7_75t_L g7476 ( 
.A(n_7434),
.B(n_7381),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_7445),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_7447),
.Y(n_7478)
);

NAND2xp5_ASAP7_75t_L g7479 ( 
.A(n_7411),
.B(n_7385),
.Y(n_7479)
);

OR2x2_ASAP7_75t_L g7480 ( 
.A(n_7458),
.B(n_7388),
.Y(n_7480)
);

AND2x4_ASAP7_75t_L g7481 ( 
.A(n_7426),
.B(n_7393),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_7418),
.Y(n_7482)
);

AND2x2_ASAP7_75t_SL g7483 ( 
.A(n_7414),
.B(n_7404),
.Y(n_7483)
);

OR2x2_ASAP7_75t_L g7484 ( 
.A(n_7427),
.B(n_7358),
.Y(n_7484)
);

HB1xp67_ASAP7_75t_L g7485 ( 
.A(n_7412),
.Y(n_7485)
);

OR2x2_ASAP7_75t_L g7486 ( 
.A(n_7429),
.B(n_7397),
.Y(n_7486)
);

AND2x2_ASAP7_75t_L g7487 ( 
.A(n_7438),
.B(n_7353),
.Y(n_7487)
);

AND2x2_ASAP7_75t_L g7488 ( 
.A(n_7455),
.B(n_7354),
.Y(n_7488)
);

INVx1_ASAP7_75t_L g7489 ( 
.A(n_7432),
.Y(n_7489)
);

BUFx2_ASAP7_75t_L g7490 ( 
.A(n_7417),
.Y(n_7490)
);

AND2x2_ASAP7_75t_L g7491 ( 
.A(n_7457),
.B(n_7405),
.Y(n_7491)
);

INVx1_ASAP7_75t_L g7492 ( 
.A(n_7437),
.Y(n_7492)
);

NAND2xp5_ASAP7_75t_L g7493 ( 
.A(n_7448),
.B(n_7394),
.Y(n_7493)
);

AOI211xp5_ASAP7_75t_L g7494 ( 
.A1(n_7407),
.A2(n_7402),
.B(n_7395),
.C(n_7397),
.Y(n_7494)
);

INVxp67_ASAP7_75t_L g7495 ( 
.A(n_7459),
.Y(n_7495)
);

NOR2x1_ASAP7_75t_L g7496 ( 
.A(n_7408),
.B(n_7400),
.Y(n_7496)
);

NAND2xp5_ASAP7_75t_L g7497 ( 
.A(n_7419),
.B(n_7400),
.Y(n_7497)
);

INVx2_ASAP7_75t_L g7498 ( 
.A(n_7454),
.Y(n_7498)
);

INVx1_ASAP7_75t_L g7499 ( 
.A(n_7441),
.Y(n_7499)
);

HB1xp67_ASAP7_75t_L g7500 ( 
.A(n_7410),
.Y(n_7500)
);

INVx1_ASAP7_75t_SL g7501 ( 
.A(n_7423),
.Y(n_7501)
);

INVx2_ASAP7_75t_L g7502 ( 
.A(n_7443),
.Y(n_7502)
);

INVx1_ASAP7_75t_L g7503 ( 
.A(n_7446),
.Y(n_7503)
);

INVx2_ASAP7_75t_L g7504 ( 
.A(n_7483),
.Y(n_7504)
);

INVx1_ASAP7_75t_L g7505 ( 
.A(n_7466),
.Y(n_7505)
);

AND2x4_ASAP7_75t_L g7506 ( 
.A(n_7477),
.B(n_7442),
.Y(n_7506)
);

INVx1_ASAP7_75t_L g7507 ( 
.A(n_7467),
.Y(n_7507)
);

NAND2xp5_ASAP7_75t_L g7508 ( 
.A(n_7500),
.B(n_7440),
.Y(n_7508)
);

INVx1_ASAP7_75t_L g7509 ( 
.A(n_7467),
.Y(n_7509)
);

HB1xp67_ASAP7_75t_L g7510 ( 
.A(n_7481),
.Y(n_7510)
);

OR2x2_ASAP7_75t_L g7511 ( 
.A(n_7476),
.B(n_7461),
.Y(n_7511)
);

OR2x2_ASAP7_75t_L g7512 ( 
.A(n_7468),
.B(n_7453),
.Y(n_7512)
);

INVx1_ASAP7_75t_L g7513 ( 
.A(n_7485),
.Y(n_7513)
);

INVx2_ASAP7_75t_L g7514 ( 
.A(n_7469),
.Y(n_7514)
);

NOR2xp33_ASAP7_75t_L g7515 ( 
.A(n_7469),
.B(n_7413),
.Y(n_7515)
);

OAI22x1_ASAP7_75t_L g7516 ( 
.A1(n_7481),
.A2(n_7420),
.B1(n_7440),
.B2(n_7452),
.Y(n_7516)
);

INVx2_ASAP7_75t_L g7517 ( 
.A(n_7472),
.Y(n_7517)
);

BUFx3_ASAP7_75t_L g7518 ( 
.A(n_7472),
.Y(n_7518)
);

NAND2xp5_ASAP7_75t_L g7519 ( 
.A(n_7465),
.B(n_7422),
.Y(n_7519)
);

INVx2_ASAP7_75t_SL g7520 ( 
.A(n_7464),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_7490),
.Y(n_7521)
);

AND3x1_ASAP7_75t_L g7522 ( 
.A(n_7496),
.B(n_7409),
.C(n_7416),
.Y(n_7522)
);

AOI21xp5_ASAP7_75t_L g7523 ( 
.A1(n_7479),
.A2(n_7416),
.B(n_7401),
.Y(n_7523)
);

AND2x4_ASAP7_75t_L g7524 ( 
.A(n_7475),
.B(n_7456),
.Y(n_7524)
);

INVx1_ASAP7_75t_SL g7525 ( 
.A(n_7484),
.Y(n_7525)
);

INVx1_ASAP7_75t_L g7526 ( 
.A(n_7487),
.Y(n_7526)
);

INVx1_ASAP7_75t_SL g7527 ( 
.A(n_7488),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_7510),
.Y(n_7528)
);

AOI322xp5_ASAP7_75t_L g7529 ( 
.A1(n_7515),
.A2(n_7470),
.A3(n_7501),
.B1(n_7462),
.B2(n_7463),
.C1(n_7474),
.C2(n_7482),
.Y(n_7529)
);

OAI22xp5_ASAP7_75t_L g7530 ( 
.A1(n_7522),
.A2(n_7471),
.B1(n_7480),
.B2(n_7473),
.Y(n_7530)
);

O2A1O1Ixp33_ASAP7_75t_L g7531 ( 
.A1(n_7523),
.A2(n_7494),
.B(n_7435),
.C(n_7493),
.Y(n_7531)
);

OAI321xp33_ASAP7_75t_L g7532 ( 
.A1(n_7519),
.A2(n_7494),
.A3(n_7497),
.B1(n_7486),
.B2(n_7495),
.C(n_7478),
.Y(n_7532)
);

AOI21x1_ASAP7_75t_L g7533 ( 
.A1(n_7516),
.A2(n_7491),
.B(n_7489),
.Y(n_7533)
);

A2O1A1Ixp33_ASAP7_75t_L g7534 ( 
.A1(n_7518),
.A2(n_7492),
.B(n_7503),
.C(n_7498),
.Y(n_7534)
);

NAND2xp5_ASAP7_75t_L g7535 ( 
.A(n_7527),
.B(n_7502),
.Y(n_7535)
);

INVxp67_ASAP7_75t_L g7536 ( 
.A(n_7522),
.Y(n_7536)
);

INVx2_ASAP7_75t_L g7537 ( 
.A(n_7514),
.Y(n_7537)
);

AND2x4_ASAP7_75t_L g7538 ( 
.A(n_7517),
.B(n_7473),
.Y(n_7538)
);

OAI221xp5_ASAP7_75t_SL g7539 ( 
.A1(n_7527),
.A2(n_7499),
.B1(n_7428),
.B2(n_7460),
.C(n_7435),
.Y(n_7539)
);

OAI222xp33_ASAP7_75t_L g7540 ( 
.A1(n_7525),
.A2(n_7521),
.B1(n_7513),
.B2(n_7504),
.C1(n_7507),
.C2(n_7509),
.Y(n_7540)
);

NAND2xp5_ASAP7_75t_L g7541 ( 
.A(n_7506),
.B(n_7520),
.Y(n_7541)
);

NAND2xp5_ASAP7_75t_L g7542 ( 
.A(n_7506),
.B(n_346),
.Y(n_7542)
);

NAND2xp5_ASAP7_75t_L g7543 ( 
.A(n_7524),
.B(n_348),
.Y(n_7543)
);

AOI22xp33_ASAP7_75t_L g7544 ( 
.A1(n_7505),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_7544)
);

INVx1_ASAP7_75t_L g7545 ( 
.A(n_7511),
.Y(n_7545)
);

AND2x4_ASAP7_75t_L g7546 ( 
.A(n_7524),
.B(n_351),
.Y(n_7546)
);

AOI22xp5_ASAP7_75t_L g7547 ( 
.A1(n_7526),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_7547)
);

AOI221xp5_ASAP7_75t_L g7548 ( 
.A1(n_7508),
.A2(n_356),
.B1(n_352),
.B2(n_355),
.C(n_358),
.Y(n_7548)
);

NAND2xp5_ASAP7_75t_L g7549 ( 
.A(n_7546),
.B(n_7519),
.Y(n_7549)
);

OAI221xp5_ASAP7_75t_L g7550 ( 
.A1(n_7536),
.A2(n_7512),
.B1(n_359),
.B2(n_355),
.C(n_356),
.Y(n_7550)
);

O2A1O1Ixp33_ASAP7_75t_L g7551 ( 
.A1(n_7530),
.A2(n_362),
.B(n_360),
.C(n_361),
.Y(n_7551)
);

NAND2xp33_ASAP7_75t_SL g7552 ( 
.A(n_7541),
.B(n_361),
.Y(n_7552)
);

INVx1_ASAP7_75t_L g7553 ( 
.A(n_7533),
.Y(n_7553)
);

INVx1_ASAP7_75t_SL g7554 ( 
.A(n_7538),
.Y(n_7554)
);

NAND2xp5_ASAP7_75t_L g7555 ( 
.A(n_7546),
.B(n_362),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_7543),
.Y(n_7556)
);

AOI221xp5_ASAP7_75t_L g7557 ( 
.A1(n_7531),
.A2(n_368),
.B1(n_364),
.B2(n_366),
.C(n_369),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_7542),
.Y(n_7558)
);

INVx1_ASAP7_75t_L g7559 ( 
.A(n_7535),
.Y(n_7559)
);

INVx2_ASAP7_75t_L g7560 ( 
.A(n_7537),
.Y(n_7560)
);

INVx1_ASAP7_75t_L g7561 ( 
.A(n_7545),
.Y(n_7561)
);

AND2x4_ASAP7_75t_L g7562 ( 
.A(n_7534),
.B(n_7547),
.Y(n_7562)
);

AOI332xp33_ASAP7_75t_L g7563 ( 
.A1(n_7540),
.A2(n_375),
.A3(n_376),
.B1(n_377),
.B2(n_378),
.B3(n_379),
.C1(n_380),
.C2(n_381),
.Y(n_7563)
);

AO22x1_ASAP7_75t_L g7564 ( 
.A1(n_7532),
.A2(n_7529),
.B1(n_7539),
.B2(n_7548),
.Y(n_7564)
);

OR2x2_ASAP7_75t_L g7565 ( 
.A(n_7544),
.B(n_375),
.Y(n_7565)
);

AND2x4_ASAP7_75t_L g7566 ( 
.A(n_7528),
.B(n_377),
.Y(n_7566)
);

NAND3xp33_ASAP7_75t_SL g7567 ( 
.A(n_7531),
.B(n_378),
.C(n_379),
.Y(n_7567)
);

AOI22xp5_ASAP7_75t_L g7568 ( 
.A1(n_7528),
.A2(n_389),
.B1(n_382),
.B2(n_388),
.Y(n_7568)
);

NAND2xp5_ASAP7_75t_L g7569 ( 
.A(n_7546),
.B(n_389),
.Y(n_7569)
);

OAI21xp5_ASAP7_75t_L g7570 ( 
.A1(n_7536),
.A2(n_390),
.B(n_391),
.Y(n_7570)
);

OAI22xp5_ASAP7_75t_L g7571 ( 
.A1(n_7553),
.A2(n_396),
.B1(n_392),
.B2(n_395),
.Y(n_7571)
);

XNOR2xp5_ASAP7_75t_L g7572 ( 
.A(n_7564),
.B(n_395),
.Y(n_7572)
);

NAND2xp5_ASAP7_75t_L g7573 ( 
.A(n_7554),
.B(n_396),
.Y(n_7573)
);

INVx1_ASAP7_75t_SL g7574 ( 
.A(n_7552),
.Y(n_7574)
);

NOR2xp33_ASAP7_75t_L g7575 ( 
.A(n_7567),
.B(n_397),
.Y(n_7575)
);

INVx1_ASAP7_75t_L g7576 ( 
.A(n_7566),
.Y(n_7576)
);

NAND2xp5_ASAP7_75t_L g7577 ( 
.A(n_7557),
.B(n_399),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_7555),
.Y(n_7578)
);

NAND2xp5_ASAP7_75t_L g7579 ( 
.A(n_7561),
.B(n_7559),
.Y(n_7579)
);

INVx2_ASAP7_75t_L g7580 ( 
.A(n_7560),
.Y(n_7580)
);

AND2x2_ASAP7_75t_L g7581 ( 
.A(n_7562),
.B(n_400),
.Y(n_7581)
);

HB1xp67_ASAP7_75t_L g7582 ( 
.A(n_7569),
.Y(n_7582)
);

AND2x2_ASAP7_75t_L g7583 ( 
.A(n_7570),
.B(n_401),
.Y(n_7583)
);

INVx1_ASAP7_75t_L g7584 ( 
.A(n_7549),
.Y(n_7584)
);

INVx1_ASAP7_75t_L g7585 ( 
.A(n_7565),
.Y(n_7585)
);

AOI22xp33_ASAP7_75t_L g7586 ( 
.A1(n_7558),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_7586)
);

AND2x2_ASAP7_75t_L g7587 ( 
.A(n_7556),
.B(n_404),
.Y(n_7587)
);

NAND2xp5_ASAP7_75t_L g7588 ( 
.A(n_7568),
.B(n_405),
.Y(n_7588)
);

AND2x2_ASAP7_75t_L g7589 ( 
.A(n_7551),
.B(n_408),
.Y(n_7589)
);

AOI221xp5_ASAP7_75t_L g7590 ( 
.A1(n_7550),
.A2(n_410),
.B1(n_412),
.B2(n_413),
.C(n_414),
.Y(n_7590)
);

INVx1_ASAP7_75t_L g7591 ( 
.A(n_7563),
.Y(n_7591)
);

AND2x2_ASAP7_75t_L g7592 ( 
.A(n_7581),
.B(n_415),
.Y(n_7592)
);

INVx1_ASAP7_75t_L g7593 ( 
.A(n_7572),
.Y(n_7593)
);

NAND2xp5_ASAP7_75t_L g7594 ( 
.A(n_7587),
.B(n_416),
.Y(n_7594)
);

NAND2xp5_ASAP7_75t_L g7595 ( 
.A(n_7576),
.B(n_418),
.Y(n_7595)
);

INVx1_ASAP7_75t_L g7596 ( 
.A(n_7573),
.Y(n_7596)
);

NOR2xp33_ASAP7_75t_L g7597 ( 
.A(n_7591),
.B(n_7574),
.Y(n_7597)
);

AND2x2_ASAP7_75t_L g7598 ( 
.A(n_7580),
.B(n_420),
.Y(n_7598)
);

NOR2x1_ASAP7_75t_L g7599 ( 
.A(n_7571),
.B(n_423),
.Y(n_7599)
);

INVx1_ASAP7_75t_SL g7600 ( 
.A(n_7589),
.Y(n_7600)
);

AOI21xp5_ASAP7_75t_L g7601 ( 
.A1(n_7579),
.A2(n_7577),
.B(n_7575),
.Y(n_7601)
);

INVx1_ASAP7_75t_L g7602 ( 
.A(n_7583),
.Y(n_7602)
);

AOI322xp5_ASAP7_75t_L g7603 ( 
.A1(n_7584),
.A2(n_424),
.A3(n_425),
.B1(n_427),
.B2(n_428),
.C1(n_429),
.C2(n_430),
.Y(n_7603)
);

OAI21xp5_ASAP7_75t_L g7604 ( 
.A1(n_7588),
.A2(n_424),
.B(n_425),
.Y(n_7604)
);

NAND2xp5_ASAP7_75t_L g7605 ( 
.A(n_7590),
.B(n_427),
.Y(n_7605)
);

NAND2xp5_ASAP7_75t_L g7606 ( 
.A(n_7586),
.B(n_431),
.Y(n_7606)
);

NOR2xp33_ASAP7_75t_L g7607 ( 
.A(n_7585),
.B(n_7582),
.Y(n_7607)
);

INVx1_ASAP7_75t_L g7608 ( 
.A(n_7578),
.Y(n_7608)
);

NAND2xp5_ASAP7_75t_L g7609 ( 
.A(n_7592),
.B(n_433),
.Y(n_7609)
);

OAI21xp5_ASAP7_75t_L g7610 ( 
.A1(n_7597),
.A2(n_434),
.B(n_435),
.Y(n_7610)
);

AOI211x1_ASAP7_75t_L g7611 ( 
.A1(n_7601),
.A2(n_438),
.B(n_435),
.C(n_437),
.Y(n_7611)
);

AOI21xp5_ASAP7_75t_L g7612 ( 
.A1(n_7605),
.A2(n_443),
.B(n_444),
.Y(n_7612)
);

NOR2x1_ASAP7_75t_L g7613 ( 
.A(n_7599),
.B(n_443),
.Y(n_7613)
);

NOR2x1_ASAP7_75t_L g7614 ( 
.A(n_7595),
.B(n_7594),
.Y(n_7614)
);

AOI211x1_ASAP7_75t_L g7615 ( 
.A1(n_7606),
.A2(n_449),
.B(n_447),
.C(n_448),
.Y(n_7615)
);

INVx1_ASAP7_75t_L g7616 ( 
.A(n_7598),
.Y(n_7616)
);

AOI21xp5_ASAP7_75t_L g7617 ( 
.A1(n_7607),
.A2(n_448),
.B(n_449),
.Y(n_7617)
);

NOR3xp33_ASAP7_75t_L g7618 ( 
.A(n_7593),
.B(n_452),
.C(n_453),
.Y(n_7618)
);

AOI21xp5_ASAP7_75t_L g7619 ( 
.A1(n_7604),
.A2(n_453),
.B(n_454),
.Y(n_7619)
);

AOI21xp5_ASAP7_75t_L g7620 ( 
.A1(n_7608),
.A2(n_455),
.B(n_456),
.Y(n_7620)
);

NOR4xp25_ASAP7_75t_L g7621 ( 
.A(n_7600),
.B(n_460),
.C(n_458),
.D(n_459),
.Y(n_7621)
);

INVx2_ASAP7_75t_L g7622 ( 
.A(n_7602),
.Y(n_7622)
);

AND2x2_ASAP7_75t_L g7623 ( 
.A(n_7596),
.B(n_467),
.Y(n_7623)
);

INVx1_ASAP7_75t_L g7624 ( 
.A(n_7609),
.Y(n_7624)
);

INVx2_ASAP7_75t_L g7625 ( 
.A(n_7623),
.Y(n_7625)
);

OAI21xp33_ASAP7_75t_L g7626 ( 
.A1(n_7622),
.A2(n_7603),
.B(n_468),
.Y(n_7626)
);

NOR2xp67_ASAP7_75t_L g7627 ( 
.A(n_7620),
.B(n_477),
.Y(n_7627)
);

OAI211xp5_ASAP7_75t_SL g7628 ( 
.A1(n_7614),
.A2(n_478),
.B(n_479),
.C(n_480),
.Y(n_7628)
);

AOI21xp33_ASAP7_75t_L g7629 ( 
.A1(n_7616),
.A2(n_479),
.B(n_480),
.Y(n_7629)
);

OAI211xp5_ASAP7_75t_SL g7630 ( 
.A1(n_7612),
.A2(n_482),
.B(n_484),
.C(n_485),
.Y(n_7630)
);

INVx1_ASAP7_75t_L g7631 ( 
.A(n_7611),
.Y(n_7631)
);

AOI211xp5_ASAP7_75t_L g7632 ( 
.A1(n_7621),
.A2(n_7619),
.B(n_7610),
.C(n_7617),
.Y(n_7632)
);

A2O1A1Ixp33_ASAP7_75t_L g7633 ( 
.A1(n_7618),
.A2(n_486),
.B(n_487),
.C(n_488),
.Y(n_7633)
);

INVx1_ASAP7_75t_L g7634 ( 
.A(n_7615),
.Y(n_7634)
);

BUFx2_ASAP7_75t_L g7635 ( 
.A(n_7613),
.Y(n_7635)
);

HB1xp67_ASAP7_75t_L g7636 ( 
.A(n_7627),
.Y(n_7636)
);

AOI22xp5_ASAP7_75t_L g7637 ( 
.A1(n_7628),
.A2(n_500),
.B1(n_502),
.B2(n_503),
.Y(n_7637)
);

AOI221xp5_ASAP7_75t_L g7638 ( 
.A1(n_7630),
.A2(n_507),
.B1(n_508),
.B2(n_509),
.C(n_510),
.Y(n_7638)
);

A2O1A1Ixp33_ASAP7_75t_SL g7639 ( 
.A1(n_7624),
.A2(n_508),
.B(n_509),
.C(n_510),
.Y(n_7639)
);

AOI221xp5_ASAP7_75t_L g7640 ( 
.A1(n_7631),
.A2(n_511),
.B1(n_512),
.B2(n_513),
.C(n_515),
.Y(n_7640)
);

AOI221xp5_ASAP7_75t_L g7641 ( 
.A1(n_7634),
.A2(n_511),
.B1(n_512),
.B2(n_515),
.C(n_517),
.Y(n_7641)
);

A2O1A1Ixp33_ASAP7_75t_SL g7642 ( 
.A1(n_7625),
.A2(n_518),
.B(n_521),
.C(n_522),
.Y(n_7642)
);

OAI221xp5_ASAP7_75t_SL g7643 ( 
.A1(n_7632),
.A2(n_524),
.B1(n_525),
.B2(n_526),
.C(n_527),
.Y(n_7643)
);

AOI21xp5_ASAP7_75t_L g7644 ( 
.A1(n_7635),
.A2(n_528),
.B(n_529),
.Y(n_7644)
);

INVx1_ASAP7_75t_L g7645 ( 
.A(n_7633),
.Y(n_7645)
);

AOI211xp5_ASAP7_75t_L g7646 ( 
.A1(n_7629),
.A2(n_532),
.B(n_533),
.C(n_534),
.Y(n_7646)
);

OAI211xp5_ASAP7_75t_L g7647 ( 
.A1(n_7626),
.A2(n_537),
.B(n_539),
.C(n_540),
.Y(n_7647)
);

AOI222xp33_ASAP7_75t_L g7648 ( 
.A1(n_7626),
.A2(n_544),
.B1(n_545),
.B2(n_547),
.C1(n_548),
.C2(n_549),
.Y(n_7648)
);

NAND4xp75_ASAP7_75t_L g7649 ( 
.A(n_7645),
.B(n_553),
.C(n_555),
.D(n_556),
.Y(n_7649)
);

NAND2xp5_ASAP7_75t_L g7650 ( 
.A(n_7644),
.B(n_555),
.Y(n_7650)
);

NAND2xp5_ASAP7_75t_L g7651 ( 
.A(n_7648),
.B(n_558),
.Y(n_7651)
);

NAND2xp5_ASAP7_75t_L g7652 ( 
.A(n_7637),
.B(n_559),
.Y(n_7652)
);

NOR3xp33_ASAP7_75t_L g7653 ( 
.A(n_7647),
.B(n_559),
.C(n_560),
.Y(n_7653)
);

NAND4xp75_ASAP7_75t_L g7654 ( 
.A(n_7638),
.B(n_564),
.C(n_565),
.D(n_566),
.Y(n_7654)
);

INVx1_ASAP7_75t_L g7655 ( 
.A(n_7636),
.Y(n_7655)
);

NAND2xp5_ASAP7_75t_SL g7656 ( 
.A(n_7646),
.B(n_568),
.Y(n_7656)
);

NOR3xp33_ASAP7_75t_L g7657 ( 
.A(n_7643),
.B(n_569),
.C(n_570),
.Y(n_7657)
);

NOR3xp33_ASAP7_75t_L g7658 ( 
.A(n_7639),
.B(n_571),
.C(n_573),
.Y(n_7658)
);

AOI221x1_ASAP7_75t_L g7659 ( 
.A1(n_7655),
.A2(n_7642),
.B1(n_7641),
.B2(n_7640),
.C(n_575),
.Y(n_7659)
);

NAND3xp33_ASAP7_75t_SL g7660 ( 
.A(n_7658),
.B(n_576),
.C(n_577),
.Y(n_7660)
);

OAI221xp5_ASAP7_75t_SL g7661 ( 
.A1(n_7653),
.A2(n_7657),
.B1(n_7651),
.B2(n_7652),
.C(n_7650),
.Y(n_7661)
);

AOI221xp5_ASAP7_75t_L g7662 ( 
.A1(n_7656),
.A2(n_585),
.B1(n_586),
.B2(n_587),
.C(n_588),
.Y(n_7662)
);

NOR2x1_ASAP7_75t_L g7663 ( 
.A(n_7649),
.B(n_586),
.Y(n_7663)
);

NAND5xp2_ASAP7_75t_L g7664 ( 
.A(n_7654),
.B(n_587),
.C(n_588),
.D(n_589),
.E(n_590),
.Y(n_7664)
);

NAND4xp75_ASAP7_75t_L g7665 ( 
.A(n_7663),
.B(n_593),
.C(n_594),
.D(n_595),
.Y(n_7665)
);

XOR2xp5_ASAP7_75t_L g7666 ( 
.A(n_7660),
.B(n_598),
.Y(n_7666)
);

AND5x1_ASAP7_75t_L g7667 ( 
.A(n_7666),
.B(n_7662),
.C(n_7661),
.D(n_7659),
.E(n_7664),
.Y(n_7667)
);

NOR2xp33_ASAP7_75t_L g7668 ( 
.A(n_7665),
.B(n_600),
.Y(n_7668)
);

OAI21xp33_ASAP7_75t_L g7669 ( 
.A1(n_7667),
.A2(n_601),
.B(n_603),
.Y(n_7669)
);

NAND5xp2_ASAP7_75t_L g7670 ( 
.A(n_7668),
.B(n_608),
.C(n_609),
.D(n_610),
.E(n_611),
.Y(n_7670)
);

NAND4xp25_ASAP7_75t_L g7671 ( 
.A(n_7669),
.B(n_610),
.C(n_611),
.D(n_614),
.Y(n_7671)
);

INVxp67_ASAP7_75t_L g7672 ( 
.A(n_7670),
.Y(n_7672)
);

NAND2xp5_ASAP7_75t_L g7673 ( 
.A(n_7669),
.B(n_617),
.Y(n_7673)
);

AOI22xp5_ASAP7_75t_L g7674 ( 
.A1(n_7671),
.A2(n_618),
.B1(n_621),
.B2(n_622),
.Y(n_7674)
);

BUFx2_ASAP7_75t_L g7675 ( 
.A(n_7673),
.Y(n_7675)
);

AND2x4_ASAP7_75t_L g7676 ( 
.A(n_7675),
.B(n_7672),
.Y(n_7676)
);

INVx1_ASAP7_75t_L g7677 ( 
.A(n_7674),
.Y(n_7677)
);

INVx2_ASAP7_75t_L g7678 ( 
.A(n_7676),
.Y(n_7678)
);

NAND2x1p5_ASAP7_75t_L g7679 ( 
.A(n_7676),
.B(n_2116),
.Y(n_7679)
);

NAND2xp5_ASAP7_75t_L g7680 ( 
.A(n_7677),
.B(n_626),
.Y(n_7680)
);

INVx1_ASAP7_75t_L g7681 ( 
.A(n_7679),
.Y(n_7681)
);

INVx1_ASAP7_75t_L g7682 ( 
.A(n_7678),
.Y(n_7682)
);

NOR2x1p5_ASAP7_75t_L g7683 ( 
.A(n_7681),
.B(n_7680),
.Y(n_7683)
);

OR2x6_ASAP7_75t_L g7684 ( 
.A(n_7682),
.B(n_2115),
.Y(n_7684)
);

INVx2_ASAP7_75t_L g7685 ( 
.A(n_7684),
.Y(n_7685)
);

AOI22xp33_ASAP7_75t_L g7686 ( 
.A1(n_7683),
.A2(n_1429),
.B1(n_1376),
.B2(n_2116),
.Y(n_7686)
);

AOI22xp5_ASAP7_75t_L g7687 ( 
.A1(n_7685),
.A2(n_2099),
.B1(n_2115),
.B2(n_2110),
.Y(n_7687)
);

OAI21xp5_ASAP7_75t_L g7688 ( 
.A1(n_7687),
.A2(n_7686),
.B(n_657),
.Y(n_7688)
);

AOI21xp5_ASAP7_75t_L g7689 ( 
.A1(n_7688),
.A2(n_2107),
.B(n_2116),
.Y(n_7689)
);

INVx1_ASAP7_75t_L g7690 ( 
.A(n_7689),
.Y(n_7690)
);

OA21x2_ASAP7_75t_L g7691 ( 
.A1(n_7690),
.A2(n_658),
.B(n_660),
.Y(n_7691)
);

OAI21xp33_ASAP7_75t_L g7692 ( 
.A1(n_7690),
.A2(n_2095),
.B(n_2099),
.Y(n_7692)
);

OAI221xp5_ASAP7_75t_R g7693 ( 
.A1(n_7692),
.A2(n_2107),
.B1(n_2099),
.B2(n_2106),
.C(n_2095),
.Y(n_7693)
);

AOI221xp5_ASAP7_75t_L g7694 ( 
.A1(n_7691),
.A2(n_2095),
.B1(n_2106),
.B2(n_2110),
.C(n_2115),
.Y(n_7694)
);

AOI22xp33_ASAP7_75t_L g7695 ( 
.A1(n_7694),
.A2(n_2095),
.B1(n_2106),
.B2(n_2110),
.Y(n_7695)
);

AOI211xp5_ASAP7_75t_L g7696 ( 
.A1(n_7695),
.A2(n_7693),
.B(n_2110),
.C(n_2115),
.Y(n_7696)
);


endmodule