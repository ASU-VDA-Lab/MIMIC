module fake_jpeg_342_n_357 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_357);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_357;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_15),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_64),
.Y(n_118)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_62),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_65),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_76),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_87),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_83),
.Y(n_120)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_81),
.Y(n_170)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_20),
.B(n_2),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_21),
.B(n_2),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_98),
.Y(n_141)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_97),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_36),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_37),
.Y(n_98)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_38),
.B1(n_31),
.B2(n_58),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_100),
.B(n_104),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_40),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_21),
.B(n_3),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_27),
.B(n_54),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_107),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_27),
.B(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_112),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_46),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_110),
.Y(n_174)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_46),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_58),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_29),
.B(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_115),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_29),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g176 ( 
.A1(n_114),
.A2(n_19),
.B(n_106),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_52),
.C(n_38),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_117),
.B(n_123),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_69),
.A2(n_57),
.B1(n_58),
.B2(n_55),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_136),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_62),
.A2(n_85),
.B1(n_97),
.B2(n_81),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_78),
.A2(n_57),
.B1(n_55),
.B2(n_54),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_79),
.A2(n_115),
.B1(n_88),
.B2(n_100),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_94),
.A2(n_33),
.B1(n_53),
.B2(n_30),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_138),
.A2(n_140),
.B1(n_151),
.B2(n_164),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_33),
.B1(n_53),
.B2(n_30),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_82),
.A2(n_39),
.B1(n_51),
.B2(n_50),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_144),
.A2(n_119),
.B(n_149),
.C(n_166),
.Y(n_186)
);

AND2x4_ASAP7_75t_L g148 ( 
.A(n_70),
.B(n_51),
.Y(n_148)
);

OR2x4_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_176),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_96),
.A2(n_56),
.B1(n_50),
.B2(n_49),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_56),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_129),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_76),
.A2(n_49),
.B1(n_47),
.B2(n_45),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_155),
.B1(n_162),
.B2(n_178),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_91),
.A2(n_110),
.B1(n_112),
.B2(n_74),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_60),
.A2(n_47),
.B1(n_45),
.B2(n_41),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_104),
.A2(n_41),
.B1(n_5),
.B2(n_6),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_99),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_169),
.A2(n_75),
.B1(n_171),
.B2(n_175),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_59),
.A2(n_10),
.B1(n_16),
.B2(n_17),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_171),
.A2(n_175),
.B1(n_148),
.B2(n_117),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_68),
.A2(n_10),
.B1(n_16),
.B2(n_17),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_148),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_71),
.A2(n_72),
.B1(n_104),
.B2(n_107),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_107),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_194),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_184),
.A2(n_190),
.B1(n_221),
.B2(n_201),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_L g246 ( 
.A1(n_186),
.A2(n_187),
.B(n_189),
.Y(n_246)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_125),
.A2(n_178),
.B1(n_166),
.B2(n_138),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_195),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_132),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_148),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_202),
.Y(n_241)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_203),
.B(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_154),
.A2(n_142),
.B1(n_132),
.B2(n_161),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_210),
.B1(n_217),
.B2(n_218),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_118),
.B(n_134),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_215),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_161),
.A2(n_170),
.B1(n_172),
.B2(n_147),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_145),
.A2(n_174),
.B1(n_116),
.B2(n_163),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_216),
.B1(n_183),
.B2(n_193),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_130),
.B(n_133),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_212),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_144),
.A2(n_168),
.B(n_167),
.C(n_158),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_173),
.Y(n_224)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

INVx13_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_135),
.B(n_143),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_144),
.B1(n_157),
.B2(n_150),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_170),
.A2(n_172),
.B1(n_143),
.B2(n_159),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_159),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_213),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_122),
.B(n_160),
.Y(n_221)
);

AOI22x1_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_122),
.B1(n_158),
.B2(n_173),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_227),
.B1(n_250),
.B2(n_195),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_121),
.B1(n_139),
.B2(n_200),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_202),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_182),
.A2(n_121),
.B1(n_139),
.B2(n_198),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_200),
.A2(n_194),
.B1(n_197),
.B2(n_211),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_231),
.A2(n_248),
.B1(n_234),
.B2(n_246),
.Y(n_260)
);

AOI211xp5_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_206),
.B(n_231),
.C(n_230),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_237),
.A2(n_244),
.B1(n_236),
.B2(n_235),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_199),
.A2(n_186),
.B1(n_219),
.B2(n_190),
.Y(n_248)
);

AO22x1_ASAP7_75t_L g249 ( 
.A1(n_199),
.A2(n_193),
.B1(n_191),
.B2(n_196),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_249),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g251 ( 
.A(n_181),
.B(n_220),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_224),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_279)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_255),
.A2(n_273),
.B1(n_252),
.B2(n_223),
.Y(n_278)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_214),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_259),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_188),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_260),
.A2(n_261),
.B(n_269),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_180),
.B1(n_179),
.B2(n_217),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_240),
.B(n_230),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_265),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_240),
.Y(n_266)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_237),
.A2(n_249),
.B1(n_222),
.B2(n_233),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_222),
.B1(n_226),
.B2(n_232),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_226),
.A2(n_229),
.B1(n_245),
.B2(n_251),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_226),
.A2(n_245),
.B1(n_242),
.B2(n_249),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_228),
.A2(n_239),
.B1(n_241),
.B2(n_247),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_275),
.A2(n_243),
.B1(n_255),
.B2(n_253),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_236),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_277),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_223),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_278),
.B(n_268),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_289),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_243),
.B1(n_272),
.B2(n_271),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_283),
.A2(n_266),
.B1(n_262),
.B2(n_277),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_269),
.A2(n_260),
.B1(n_263),
.B2(n_257),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_267),
.A2(n_254),
.B(n_256),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_290),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_267),
.A2(n_264),
.B(n_258),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_293),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_273),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_274),
.Y(n_306)
);

AOI221xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_284),
.B1(n_289),
.B2(n_291),
.C(n_290),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_296),
.A2(n_306),
.B1(n_278),
.B2(n_287),
.Y(n_318)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_292),
.Y(n_298)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_302),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_284),
.B1(n_287),
.B2(n_291),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_276),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_293),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_307),
.Y(n_312)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_288),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_308),
.B1(n_283),
.B2(n_279),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_300),
.A2(n_279),
.B1(n_283),
.B2(n_290),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_313),
.A2(n_310),
.B1(n_299),
.B2(n_308),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_286),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_316),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_322),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_297),
.B(n_281),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_304),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_288),
.C(n_285),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_323),
.A2(n_329),
.B1(n_320),
.B2(n_315),
.Y(n_338)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_325),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_298),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_327),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_311),
.A2(n_310),
.B1(n_308),
.B2(n_301),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_302),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_314),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_324),
.B(n_306),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_334),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_322),
.C(n_313),
.Y(n_334)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_336),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_SL g337 ( 
.A(n_331),
.B(n_312),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_337),
.B(n_338),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_334),
.B(n_329),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_323),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_332),
.A2(n_324),
.B(n_328),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_342),
.A2(n_343),
.B(n_325),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_327),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_340),
.A2(n_335),
.B(n_327),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_345),
.A2(n_314),
.B(n_315),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_347),
.C(n_348),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_328),
.C(n_330),
.Y(n_348)
);

AO221x1_ASAP7_75t_L g350 ( 
.A1(n_347),
.A2(n_343),
.B1(n_339),
.B2(n_278),
.C(n_326),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_351),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_349),
.B(n_282),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_352),
.B(n_282),
.Y(n_354)
);

AOI321xp33_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_353),
.A3(n_320),
.B1(n_285),
.B2(n_309),
.C(n_307),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_305),
.C(n_280),
.Y(n_356)
);

BUFx24_ASAP7_75t_SL g357 ( 
.A(n_356),
.Y(n_357)
);


endmodule