module fake_jpeg_10651_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_17),
.B1(n_24),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_17),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_17),
.B1(n_24),
.B2(n_30),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_17),
.B1(n_24),
.B2(n_27),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_67),
.A2(n_35),
.B1(n_28),
.B2(n_16),
.Y(n_118)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_69),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_71),
.Y(n_104)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_73),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_76),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_80),
.Y(n_115)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_86),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_45),
.B1(n_39),
.B2(n_40),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_25),
.B1(n_23),
.B2(n_44),
.Y(n_103)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_96),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_90),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_43),
.B1(n_24),
.B2(n_39),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_91),
.B1(n_68),
.B2(n_70),
.Y(n_106)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_43),
.B1(n_40),
.B2(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_40),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_35),
.B1(n_65),
.B2(n_46),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_115),
.B1(n_104),
.B2(n_117),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_29),
.B1(n_20),
.B2(n_22),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_110),
.B1(n_30),
.B2(n_29),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_35),
.B1(n_46),
.B2(n_53),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_118),
.B1(n_119),
.B2(n_25),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_93),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_111),
.B(n_117),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_35),
.B(n_46),
.C(n_27),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_34),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_19),
.B1(n_29),
.B2(n_30),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_44),
.B(n_21),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_25),
.B(n_19),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_75),
.A2(n_71),
.B1(n_85),
.B2(n_89),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_125),
.B(n_21),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_44),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_78),
.Y(n_157)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_81),
.A3(n_89),
.B1(n_44),
.B2(n_74),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_128),
.A2(n_130),
.B(n_136),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_129),
.B(n_139),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_98),
.C(n_95),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_132),
.C(n_135),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_121),
.B(n_90),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_147),
.B1(n_156),
.B2(n_22),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_12),
.C(n_15),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_134),
.B(n_140),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_44),
.C(n_42),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_44),
.C(n_42),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_145),
.C(n_151),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_96),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_12),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_94),
.B1(n_97),
.B2(n_73),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_152),
.B1(n_153),
.B2(n_104),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_37),
.Y(n_144)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_108),
.C(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_37),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_149),
.Y(n_181)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_150),
.A2(n_157),
.B(n_105),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_42),
.C(n_37),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_102),
.A2(n_36),
.B1(n_42),
.B2(n_37),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_130),
.A3(n_155),
.B1(n_139),
.B2(n_142),
.Y(n_161)
);

AO21x2_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_55),
.B(n_34),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_112),
.B1(n_101),
.B2(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_103),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_159),
.A2(n_161),
.B1(n_167),
.B2(n_175),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_99),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_160),
.B(n_188),
.C(n_190),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_169),
.B1(n_184),
.B2(n_101),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_166),
.B(n_168),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_102),
.B1(n_103),
.B2(n_125),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_107),
.B1(n_125),
.B2(n_106),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_170),
.A2(n_179),
.B1(n_187),
.B2(n_33),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_172),
.B(n_176),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_155),
.A2(n_105),
.B1(n_114),
.B2(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_182),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_129),
.B1(n_133),
.B2(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_183),
.A2(n_192),
.B(n_113),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_100),
.B1(n_112),
.B2(n_127),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_172),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_128),
.A2(n_119),
.B1(n_114),
.B2(n_124),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_36),
.C(n_113),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_101),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_189),
.B(n_176),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_136),
.B(n_36),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_143),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_199),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_198),
.C(n_200),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_36),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_175),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_18),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_201),
.B(n_208),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_203),
.A2(n_212),
.B1(n_170),
.B2(n_165),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_113),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_206),
.A2(n_180),
.B1(n_193),
.B2(n_33),
.Y(n_237)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_216),
.C(n_32),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_16),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_192),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_211),
.B(n_214),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_163),
.A2(n_26),
.B1(n_33),
.B2(n_32),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_16),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_18),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_162),
.B(n_18),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_21),
.B1(n_55),
.B2(n_2),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_26),
.B(n_1),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_7),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_171),
.A2(n_21),
.B(n_1),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_223),
.B1(n_21),
.B2(n_8),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_171),
.A2(n_162),
.B(n_186),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_190),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_228),
.C(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_223),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_231),
.A2(n_238),
.B1(n_218),
.B2(n_204),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_161),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_167),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_241),
.C(n_247),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_242),
.B1(n_246),
.B2(n_218),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_208),
.A2(n_33),
.B1(n_32),
.B2(n_16),
.Y(n_238)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_8),
.C(n_15),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_245),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_55),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_0),
.C(n_2),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_8),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_194),
.C(n_215),
.Y(n_267)
);

AO22x1_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_199),
.B1(n_217),
.B2(n_214),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_251),
.A2(n_271),
.B(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_270),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_220),
.B(n_201),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_255),
.B(n_269),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_197),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_263),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_207),
.B1(n_217),
.B2(n_196),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_221),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_202),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_265),
.C(n_232),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_268),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_248),
.Y(n_282)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_227),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_272),
.B(n_256),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_195),
.B(n_234),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_276),
.B1(n_247),
.B2(n_256),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_240),
.B(n_230),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_257),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_257),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_241),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_278),
.C(n_280),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_11),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_213),
.B1(n_210),
.B2(n_242),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_285),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_261),
.Y(n_286)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_303),
.C(n_283),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_267),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_298),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_262),
.Y(n_294)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_258),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_299),
.B1(n_286),
.B2(n_281),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_273),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_13),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_9),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_302),
.Y(n_310)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_314),
.C(n_315),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_308),
.B(n_311),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_288),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_298),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_280),
.C(n_272),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_275),
.C(n_282),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_305),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_318),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_304),
.A2(n_292),
.B1(n_293),
.B2(n_297),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_9),
.C(n_3),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_323),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_0),
.B(n_4),
.Y(n_322)
);

A2O1A1O1Ixp25_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_308),
.B(n_310),
.C(n_5),
.D(n_6),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_4),
.C(n_5),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_309),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_319),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_5),
.Y(n_332)
);

NOR2x1_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_317),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_331),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_333),
.B(n_330),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_312),
.C(n_326),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_328),
.C(n_332),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_325),
.B(n_6),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_6),
.Y(n_339)
);


endmodule