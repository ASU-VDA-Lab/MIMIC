module fake_jpeg_14356_n_561 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_561);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_561;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVxp33_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_53),
.B(n_57),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_55),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_56),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_17),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g122 ( 
.A(n_58),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_80),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_16),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_79),
.Y(n_109)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_67),
.Y(n_121)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_16),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_35),
.A2(n_0),
.B(n_1),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_51),
.C(n_36),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_90),
.Y(n_126)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_3),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_22),
.B(n_2),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_95),
.Y(n_129)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_93),
.Y(n_130)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_22),
.B(n_2),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_96),
.Y(n_156)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_21),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_105),
.Y(n_134)
);

INVx2_ASAP7_75t_R g100 ( 
.A(n_44),
.Y(n_100)
);

OR2x4_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_44),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_21),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_21),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_32),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_110),
.B(n_38),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_45),
.B1(n_49),
.B2(n_47),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_111),
.A2(n_61),
.B1(n_60),
.B2(n_98),
.Y(n_181)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_67),
.Y(n_112)
);

INVx5_ASAP7_75t_SL g175 ( 
.A(n_112),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_19),
.C(n_42),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_117),
.B(n_94),
.C(n_84),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_125),
.B(n_40),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_135),
.B(n_97),
.Y(n_207)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_88),
.A2(n_82),
.B1(n_66),
.B2(n_65),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_139),
.A2(n_144),
.B1(n_39),
.B2(n_34),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_77),
.A2(n_39),
.B1(n_50),
.B2(n_34),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_51),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_72),
.B(n_23),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_164),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_87),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_56),
.Y(n_162)
);

CKINVDCx9p33_ASAP7_75t_R g184 ( 
.A(n_162),
.Y(n_184)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_58),
.Y(n_164)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_58),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_170),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_61),
.B(n_40),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_109),
.A2(n_111),
.B1(n_91),
.B2(n_81),
.Y(n_173)
);

AOI22x1_ASAP7_75t_L g240 ( 
.A1(n_173),
.A2(n_177),
.B1(n_157),
.B2(n_119),
.Y(n_240)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g282 ( 
.A(n_174),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g259 ( 
.A(n_176),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_75),
.B1(n_101),
.B2(n_71),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

OR2x4_ASAP7_75t_L g180 ( 
.A(n_115),
.B(n_102),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_180),
.A2(n_201),
.B(n_207),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_181),
.Y(n_268)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_145),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_186),
.B(n_205),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_118),
.A2(n_42),
.B1(n_23),
.B2(n_33),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_189),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_128),
.A2(n_89),
.B1(n_55),
.B2(n_59),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_190),
.A2(n_198),
.B1(n_217),
.B2(n_159),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_126),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_192),
.B(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

CKINVDCx9p33_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_197),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_146),
.A2(n_63),
.B1(n_54),
.B2(n_36),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_203),
.Y(n_283)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_206),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_129),
.B(n_96),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_208),
.B(n_210),
.Y(n_269)
);

CKINVDCx9p33_ASAP7_75t_R g209 ( 
.A(n_130),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_209),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_114),
.B(n_96),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_211),
.Y(n_278)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_212),
.Y(n_280)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_215),
.Y(n_272)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_221),
.Y(n_256)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_132),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_151),
.A2(n_78),
.B1(n_34),
.B2(n_50),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_218),
.A2(n_220),
.B1(n_226),
.B2(n_230),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_133),
.A2(n_33),
.B1(n_20),
.B2(n_49),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_108),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_119),
.B(n_20),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_150),
.Y(n_253)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_122),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_223),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_228),
.Y(n_260)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_107),
.A2(n_49),
.B1(n_47),
.B2(n_45),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_147),
.A2(n_38),
.B(n_47),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_107),
.B(n_74),
.Y(n_263)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_116),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_121),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_231),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_116),
.A2(n_46),
.B1(n_50),
.B2(n_86),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_157),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_87),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_161),
.C(n_156),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_257),
.C(n_279),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_124),
.B(n_73),
.C(n_160),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_235),
.B(n_254),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_187),
.B(n_143),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_238),
.B(n_270),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_240),
.A2(n_274),
.B1(n_276),
.B2(n_184),
.Y(n_301)
);

NAND2xp33_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_124),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g302 ( 
.A1(n_243),
.A2(n_262),
.B(n_184),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_253),
.B(n_284),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_201),
.B(n_160),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_201),
.B(n_156),
.C(n_136),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_173),
.A2(n_199),
.B1(n_177),
.B2(n_222),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_267),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_193),
.B(n_150),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_209),
.Y(n_286)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_172),
.A2(n_155),
.B(n_143),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_195),
.B(n_155),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_175),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_191),
.B(n_155),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_273),
.B(n_277),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_217),
.A2(n_136),
.B1(n_142),
.B2(n_137),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_180),
.B(n_46),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_194),
.B(n_73),
.C(n_137),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_142),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_287),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_182),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_176),
.C(n_175),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_290),
.B(n_279),
.C(n_250),
.Y(n_346)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_185),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_292),
.B(n_305),
.Y(n_334)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_293),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_179),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_294),
.B(n_308),
.Y(n_348)
);

BUFx12_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_295),
.Y(n_350)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_298),
.Y(n_339)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_299),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_268),
.A2(n_176),
.B1(n_197),
.B2(n_229),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_300),
.A2(n_282),
.B(n_174),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_301),
.A2(n_326),
.B1(n_258),
.B2(n_281),
.Y(n_341)
);

AO21x1_ASAP7_75t_L g365 ( 
.A1(n_302),
.A2(n_313),
.B(n_272),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_303),
.Y(n_359)
);

AND2x6_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_176),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_304),
.B(n_306),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_247),
.Y(n_305)
);

AND2x6_ASAP7_75t_L g306 ( 
.A(n_235),
.B(n_196),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_241),
.Y(n_307)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_307),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_212),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_242),
.Y(n_310)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_310),
.Y(n_369)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_311),
.Y(n_370)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_243),
.B(n_223),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_312),
.B(n_328),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_263),
.B(n_257),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_236),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_314),
.B(n_317),
.Y(n_337)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_255),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_240),
.A2(n_159),
.B1(n_113),
.B2(n_231),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_316),
.A2(n_325),
.B1(n_245),
.B2(n_271),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_275),
.B(n_185),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_269),
.B(n_213),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_318),
.B(n_322),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_239),
.B(n_183),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_321),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_233),
.B(n_183),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_238),
.B(n_203),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_259),
.Y(n_323)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_261),
.B(n_211),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_324),
.B(n_327),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_240),
.A2(n_113),
.B1(n_224),
.B2(n_178),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_276),
.A2(n_46),
.B1(n_202),
.B2(n_215),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_242),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_271),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_261),
.B(n_188),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_329),
.Y(n_345)
);

INVx13_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_330),
.Y(n_362)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_332),
.Y(n_358)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g340 ( 
.A1(n_301),
.A2(n_245),
.B1(n_258),
.B2(n_274),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_367),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_341),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_342),
.A2(n_352),
.B1(n_366),
.B2(n_372),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_285),
.A2(n_268),
.B(n_277),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_343),
.A2(n_296),
.B(n_303),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_346),
.B(n_225),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_264),
.B(n_248),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_351),
.A2(n_303),
.B(n_300),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_325),
.A2(n_244),
.B1(n_248),
.B2(n_272),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_289),
.B(n_256),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_361),
.C(n_373),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_308),
.A2(n_260),
.B1(n_244),
.B2(n_251),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_364),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_295),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_360),
.B(n_282),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_289),
.B(n_266),
.C(n_272),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_294),
.B(n_266),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_SL g389 ( 
.A1(n_365),
.A2(n_286),
.B(n_290),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_316),
.A2(n_278),
.B1(n_251),
.B2(n_252),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_313),
.A2(n_278),
.B1(n_252),
.B2(n_283),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_321),
.B(n_285),
.C(n_320),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_295),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_188),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_358),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_386),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_377),
.A2(n_343),
.B(n_346),
.Y(n_422)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_378),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_371),
.Y(n_379)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_379),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_320),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_381),
.B(n_388),
.C(n_396),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_382),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_304),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_383),
.A2(n_389),
.B(n_399),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_287),
.Y(n_384)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_372),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_285),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_336),
.B(n_288),
.Y(n_390)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_390),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_336),
.B(n_291),
.Y(n_392)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_392),
.Y(n_443)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_393),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_349),
.B(n_299),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_402),
.Y(n_424)
);

OAI22x1_ASAP7_75t_SL g395 ( 
.A1(n_342),
.A2(n_306),
.B1(n_312),
.B2(n_326),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_395),
.A2(n_400),
.B1(n_407),
.B2(n_357),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_319),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_334),
.B(n_309),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_397),
.B(n_403),
.Y(n_442)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_347),
.Y(n_398)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_398),
.Y(n_415)
);

OAI21xp33_ASAP7_75t_SL g400 ( 
.A1(n_359),
.A2(n_307),
.B(n_297),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_356),
.A2(n_332),
.B1(n_331),
.B2(n_311),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_283),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_352),
.A2(n_314),
.B1(n_315),
.B2(n_323),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_406),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_255),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_405),
.B(n_362),
.Y(n_437)
);

AND2x6_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_330),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_349),
.A2(n_298),
.B1(n_234),
.B2(n_204),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_348),
.B(n_234),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_353),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_337),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_411),
.A2(n_375),
.B1(n_399),
.B2(n_377),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_378),
.A2(n_348),
.B1(n_366),
.B2(n_340),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_412),
.A2(n_434),
.B1(n_438),
.B2(n_413),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g419 ( 
.A1(n_380),
.A2(n_340),
.B(n_367),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_419),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_345),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_420),
.B(n_429),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_351),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_428),
.Y(n_452)
);

NOR3xp33_ASAP7_75t_L g467 ( 
.A(n_422),
.B(n_440),
.C(n_171),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_394),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_396),
.B(n_350),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_431),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_374),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_432),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_433),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_409),
.A2(n_340),
.B1(n_347),
.B2(n_353),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_362),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_441),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_405),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_409),
.A2(n_370),
.B1(n_338),
.B2(n_369),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g440 ( 
.A(n_401),
.B(n_338),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_368),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_445),
.A2(n_429),
.B1(n_413),
.B2(n_443),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_426),
.A2(n_380),
.B1(n_391),
.B2(n_406),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_446),
.A2(n_468),
.B1(n_450),
.B2(n_465),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_447),
.A2(n_450),
.B1(n_455),
.B2(n_457),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_442),
.B(n_368),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_448),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_412),
.A2(n_395),
.B1(n_380),
.B2(n_375),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_423),
.A2(n_383),
.B(n_405),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_451),
.A2(n_467),
.B(n_469),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_421),
.B(n_381),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_453),
.B(n_430),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_434),
.A2(n_384),
.B1(n_408),
.B2(n_398),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_427),
.Y(n_456)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_456),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_419),
.A2(n_393),
.B1(n_385),
.B2(n_401),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_459),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_370),
.Y(n_460)
);

MAJx2_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_439),
.C(n_424),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_418),
.B(n_369),
.C(n_339),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_466),
.C(n_437),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_422),
.B(n_339),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_424),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_419),
.A2(n_344),
.B1(n_335),
.B2(n_246),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_465),
.A2(n_468),
.B1(n_470),
.B2(n_411),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_428),
.B(n_344),
.C(n_216),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_426),
.A2(n_335),
.B1(n_246),
.B2(n_171),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_423),
.A2(n_3),
.B(n_4),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_433),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_417),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_488),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_473),
.A2(n_484),
.B1(n_7),
.B2(n_8),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_444),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_475),
.A2(n_481),
.B1(n_483),
.B2(n_485),
.Y(n_511)
);

BUFx24_ASAP7_75t_SL g477 ( 
.A(n_451),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_477),
.B(n_489),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_478),
.A2(n_447),
.B1(n_469),
.B2(n_425),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_479),
.B(n_487),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_482),
.C(n_490),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_471),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_446),
.A2(n_439),
.B1(n_443),
.B2(n_416),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_452),
.B(n_430),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_457),
.B(n_437),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_455),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_416),
.C(n_425),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_452),
.Y(n_502)
);

AND2x2_ASAP7_75t_SL g493 ( 
.A(n_463),
.B(n_415),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_7),
.B(n_8),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_478),
.A2(n_449),
.B(n_459),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_495),
.A2(n_506),
.B(n_507),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_476),
.A2(n_449),
.B(n_462),
.C(n_459),
.Y(n_497)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_497),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_498),
.A2(n_500),
.B1(n_511),
.B2(n_486),
.Y(n_514)
);

AOI221xp5_ASAP7_75t_L g499 ( 
.A1(n_491),
.A2(n_458),
.B1(n_464),
.B2(n_438),
.C(n_436),
.Y(n_499)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_499),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_486),
.A2(n_466),
.B1(n_436),
.B2(n_415),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_508),
.Y(n_515)
);

OAI321xp33_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_414),
.A3(n_453),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_503)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_503),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_414),
.C(n_4),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_SL g526 ( 
.A(n_504),
.B(n_510),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_3),
.Y(n_505)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_505),
.Y(n_527)
);

A2O1A1O1Ixp25_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_3),
.B(n_4),
.C(n_6),
.D(n_7),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_487),
.B(n_8),
.C(n_9),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_472),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_520),
.Y(n_533)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_514),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_474),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_517),
.B(n_519),
.Y(n_539)
);

BUFx24_ASAP7_75t_SL g519 ( 
.A(n_497),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_496),
.B(n_488),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_493),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_493),
.Y(n_532)
);

NOR2x1_ASAP7_75t_SL g522 ( 
.A(n_501),
.B(n_479),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_522),
.A2(n_504),
.B1(n_510),
.B2(n_502),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_500),
.C(n_509),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_523),
.B(n_528),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_507),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_518),
.A2(n_495),
.B1(n_508),
.B2(n_498),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_530),
.B(n_534),
.Y(n_544)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_527),
.Y(n_531)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_531),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_532),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_506),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_536),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_523),
.B(n_482),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_537),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_14),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_538),
.A2(n_540),
.B1(n_525),
.B2(n_515),
.Y(n_547)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_516),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_520),
.C(n_513),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_543),
.B(n_547),
.Y(n_551)
);

NAND4xp25_ASAP7_75t_L g548 ( 
.A(n_542),
.B(n_536),
.C(n_529),
.D(n_525),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_R g554 ( 
.A(n_548),
.B(n_543),
.Y(n_554)
);

AOI322xp5_ASAP7_75t_L g549 ( 
.A1(n_541),
.A2(n_539),
.A3(n_530),
.B1(n_533),
.B2(n_515),
.C1(n_532),
.C2(n_521),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_549),
.B(n_550),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_544),
.A2(n_533),
.B(n_10),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_551),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_553),
.B(n_554),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_552),
.B(n_544),
.C(n_545),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_556),
.A2(n_546),
.B(n_11),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_557),
.Y(n_558)
);

BUFx24_ASAP7_75t_SL g559 ( 
.A(n_558),
.Y(n_559)
);

OAI222xp33_ASAP7_75t_L g560 ( 
.A1(n_559),
.A2(n_555),
.B1(n_11),
.B2(n_12),
.C1(n_14),
.C2(n_9),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_560),
.A2(n_12),
.B(n_556),
.Y(n_561)
);


endmodule