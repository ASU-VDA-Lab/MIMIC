module fake_netlist_1_1793_n_1478 (n_107, n_156, n_154, n_239, n_7, n_309, n_356, n_327, n_25, n_204, n_169, n_180, n_99, n_43, n_73, n_199, n_279, n_357, n_74, n_308, n_44, n_189, n_226, n_352, n_66, n_316, n_285, n_47, n_281, n_11, n_295, n_139, n_342, n_151, n_71, n_288, n_176, n_359, n_195, n_300, n_223, n_19, n_261, n_220, n_353, n_104, n_303, n_159, n_91, n_301, n_340, n_148, n_149, n_246, n_191, n_143, n_63, n_54, n_125, n_145, n_166, n_181, n_123, n_219, n_343, n_135, n_315, n_53, n_213, n_196, n_293, n_127, n_312, n_23, n_110, n_182, n_269, n_186, n_137, n_334, n_164, n_120, n_155, n_162, n_114, n_50, n_3, n_331, n_330, n_231, n_9, n_178, n_229, n_97, n_133, n_324, n_192, n_329, n_6, n_8, n_187, n_188, n_304, n_18, n_314, n_307, n_215, n_172, n_109, n_332, n_198, n_351, n_1, n_16, n_95, n_40, n_210, n_228, n_278, n_115, n_270, n_179, n_289, n_354, n_152, n_70, n_17, n_322, n_317, n_221, n_328, n_266, n_80, n_326, n_275, n_274, n_150, n_235, n_38, n_272, n_100, n_299, n_280, n_141, n_160, n_263, n_193, n_232, n_344, n_147, n_185, n_267, n_171, n_140, n_111, n_212, n_30, n_13, n_254, n_64, n_69, n_248, n_83, n_200, n_262, n_119, n_339, n_347, n_124, n_79, n_129, n_157, n_103, n_52, n_253, n_273, n_325, n_163, n_348, n_96, n_72, n_77, n_90, n_214, n_167, n_33, n_76, n_61, n_216, n_153, n_355, n_121, n_286, n_247, n_161, n_224, n_165, n_65, n_5, n_211, n_85, n_320, n_264, n_102, n_283, n_290, n_217, n_201, n_277, n_259, n_244, n_276, n_297, n_225, n_350, n_208, n_252, n_168, n_271, n_94, n_194, n_282, n_58, n_113, n_242, n_284, n_321, n_302, n_116, n_292, n_118, n_233, n_257, n_26, n_203, n_243, n_318, n_346, n_98, n_345, n_230, n_146, n_337, n_32, n_93, n_41, n_10, n_75, n_82, n_183, n_132, n_170, n_205, n_158, n_126, n_249, n_360, n_106, n_296, n_42, n_21, n_89, n_130, n_310, n_341, n_14, n_236, n_136, n_260, n_222, n_34, n_142, n_227, n_250, n_268, n_190, n_62, n_4, n_59, n_323, n_240, n_88, n_46, n_174, n_108, n_335, n_37, n_122, n_87, n_349, n_207, n_197, n_81, n_298, n_112, n_78, n_68, n_105, n_251, n_36, n_237, n_15, n_256, n_117, n_238, n_294, n_2, n_338, n_209, n_241, n_20, n_84, n_12, n_56, n_67, n_22, n_311, n_202, n_319, n_39, n_101, n_291, n_245, n_24, n_35, n_134, n_48, n_255, n_55, n_336, n_29, n_218, n_173, n_60, n_138, n_305, n_92, n_313, n_333, n_358, n_175, n_128, n_306, n_0, n_258, n_234, n_184, n_265, n_57, n_51, n_287, n_144, n_45, n_131, n_86, n_27, n_177, n_28, n_49, n_206, n_31, n_1478, n_912);
input n_107;
input n_156;
input n_154;
input n_239;
input n_7;
input n_309;
input n_356;
input n_327;
input n_25;
input n_204;
input n_169;
input n_180;
input n_99;
input n_43;
input n_73;
input n_199;
input n_279;
input n_357;
input n_74;
input n_308;
input n_44;
input n_189;
input n_226;
input n_352;
input n_66;
input n_316;
input n_285;
input n_47;
input n_281;
input n_11;
input n_295;
input n_139;
input n_342;
input n_151;
input n_71;
input n_288;
input n_176;
input n_359;
input n_195;
input n_300;
input n_223;
input n_19;
input n_261;
input n_220;
input n_353;
input n_104;
input n_303;
input n_159;
input n_91;
input n_301;
input n_340;
input n_148;
input n_149;
input n_246;
input n_191;
input n_143;
input n_63;
input n_54;
input n_125;
input n_145;
input n_166;
input n_181;
input n_123;
input n_219;
input n_343;
input n_135;
input n_315;
input n_53;
input n_213;
input n_196;
input n_293;
input n_127;
input n_312;
input n_23;
input n_110;
input n_182;
input n_269;
input n_186;
input n_137;
input n_334;
input n_164;
input n_120;
input n_155;
input n_162;
input n_114;
input n_50;
input n_3;
input n_331;
input n_330;
input n_231;
input n_9;
input n_178;
input n_229;
input n_97;
input n_133;
input n_324;
input n_192;
input n_329;
input n_6;
input n_8;
input n_187;
input n_188;
input n_304;
input n_18;
input n_314;
input n_307;
input n_215;
input n_172;
input n_109;
input n_332;
input n_198;
input n_351;
input n_1;
input n_16;
input n_95;
input n_40;
input n_210;
input n_228;
input n_278;
input n_115;
input n_270;
input n_179;
input n_289;
input n_354;
input n_152;
input n_70;
input n_17;
input n_322;
input n_317;
input n_221;
input n_328;
input n_266;
input n_80;
input n_326;
input n_275;
input n_274;
input n_150;
input n_235;
input n_38;
input n_272;
input n_100;
input n_299;
input n_280;
input n_141;
input n_160;
input n_263;
input n_193;
input n_232;
input n_344;
input n_147;
input n_185;
input n_267;
input n_171;
input n_140;
input n_111;
input n_212;
input n_30;
input n_13;
input n_254;
input n_64;
input n_69;
input n_248;
input n_83;
input n_200;
input n_262;
input n_119;
input n_339;
input n_347;
input n_124;
input n_79;
input n_129;
input n_157;
input n_103;
input n_52;
input n_253;
input n_273;
input n_325;
input n_163;
input n_348;
input n_96;
input n_72;
input n_77;
input n_90;
input n_214;
input n_167;
input n_33;
input n_76;
input n_61;
input n_216;
input n_153;
input n_355;
input n_121;
input n_286;
input n_247;
input n_161;
input n_224;
input n_165;
input n_65;
input n_5;
input n_211;
input n_85;
input n_320;
input n_264;
input n_102;
input n_283;
input n_290;
input n_217;
input n_201;
input n_277;
input n_259;
input n_244;
input n_276;
input n_297;
input n_225;
input n_350;
input n_208;
input n_252;
input n_168;
input n_271;
input n_94;
input n_194;
input n_282;
input n_58;
input n_113;
input n_242;
input n_284;
input n_321;
input n_302;
input n_116;
input n_292;
input n_118;
input n_233;
input n_257;
input n_26;
input n_203;
input n_243;
input n_318;
input n_346;
input n_98;
input n_345;
input n_230;
input n_146;
input n_337;
input n_32;
input n_93;
input n_41;
input n_10;
input n_75;
input n_82;
input n_183;
input n_132;
input n_170;
input n_205;
input n_158;
input n_126;
input n_249;
input n_360;
input n_106;
input n_296;
input n_42;
input n_21;
input n_89;
input n_130;
input n_310;
input n_341;
input n_14;
input n_236;
input n_136;
input n_260;
input n_222;
input n_34;
input n_142;
input n_227;
input n_250;
input n_268;
input n_190;
input n_62;
input n_4;
input n_59;
input n_323;
input n_240;
input n_88;
input n_46;
input n_174;
input n_108;
input n_335;
input n_37;
input n_122;
input n_87;
input n_349;
input n_207;
input n_197;
input n_81;
input n_298;
input n_112;
input n_78;
input n_68;
input n_105;
input n_251;
input n_36;
input n_237;
input n_15;
input n_256;
input n_117;
input n_238;
input n_294;
input n_2;
input n_338;
input n_209;
input n_241;
input n_20;
input n_84;
input n_12;
input n_56;
input n_67;
input n_22;
input n_311;
input n_202;
input n_319;
input n_39;
input n_101;
input n_291;
input n_245;
input n_24;
input n_35;
input n_134;
input n_48;
input n_255;
input n_55;
input n_336;
input n_29;
input n_218;
input n_173;
input n_60;
input n_138;
input n_305;
input n_92;
input n_313;
input n_333;
input n_358;
input n_175;
input n_128;
input n_306;
input n_0;
input n_258;
input n_234;
input n_184;
input n_265;
input n_57;
input n_51;
input n_287;
input n_144;
input n_45;
input n_131;
input n_86;
input n_27;
input n_177;
input n_28;
input n_49;
input n_206;
input n_31;
output n_1478;
output n_912;
wire n_890;
wire n_107;
wire n_759;
wire n_987;
wire n_658;
wire n_1202;
wire n_309;
wire n_1401;
wire n_356;
wire n_327;
wire n_1267;
wire n_1084;
wire n_1041;
wire n_169;
wire n_384;
wire n_959;
wire n_1152;
wire n_279;
wire n_1129;
wire n_1149;
wire n_357;
wire n_1207;
wire n_886;
wire n_595;
wire n_875;
wire n_952;
wire n_1451;
wire n_47;
wire n_766;
wire n_744;
wire n_1448;
wire n_399;
wire n_1452;
wire n_942;
wire n_295;
wire n_1474;
wire n_139;
wire n_151;
wire n_900;
wire n_869;
wire n_935;
wire n_359;
wire n_300;
wire n_487;
wire n_405;
wire n_482;
wire n_1050;
wire n_707;
wire n_1450;
wire n_220;
wire n_1467;
wire n_1471;
wire n_159;
wire n_301;
wire n_340;
wire n_963;
wire n_1278;
wire n_246;
wire n_676;
wire n_143;
wire n_446;
wire n_402;
wire n_54;
wire n_876;
wire n_1324;
wire n_1198;
wire n_145;
wire n_1412;
wire n_166;
wire n_1059;
wire n_621;
wire n_1445;
wire n_981;
wire n_213;
wire n_196;
wire n_1167;
wire n_1089;
wire n_1286;
wire n_1045;
wire n_424;
wire n_110;
wire n_1019;
wire n_1374;
wire n_1468;
wire n_1024;
wire n_660;
wire n_433;
wire n_392;
wire n_155;
wire n_1171;
wire n_331;
wire n_814;
wire n_678;
wire n_991;
wire n_1091;
wire n_133;
wire n_1244;
wire n_1367;
wire n_548;
wire n_443;
wire n_304;
wire n_682;
wire n_1402;
wire n_441;
wire n_868;
wire n_920;
wire n_517;
wire n_386;
wire n_1209;
wire n_653;
wire n_351;
wire n_1;
wire n_1218;
wire n_829;
wire n_984;
wire n_366;
wire n_837;
wire n_549;
wire n_720;
wire n_1092;
wire n_17;
wire n_221;
wire n_711;
wire n_773;
wire n_266;
wire n_1311;
wire n_793;
wire n_679;
wire n_684;
wire n_879;
wire n_544;
wire n_275;
wire n_691;
wire n_1122;
wire n_274;
wire n_1407;
wire n_1110;
wire n_1464;
wire n_38;
wire n_965;
wire n_100;
wire n_1277;
wire n_844;
wire n_695;
wire n_344;
wire n_878;
wire n_367;
wire n_795;
wire n_687;
wire n_212;
wire n_1203;
wire n_728;
wire n_254;
wire n_704;
wire n_435;
wire n_841;
wire n_69;
wire n_1021;
wire n_1454;
wire n_1186;
wire n_1300;
wire n_1012;
wire n_124;
wire n_1463;
wire n_1175;
wire n_1127;
wire n_1423;
wire n_1386;
wire n_904;
wire n_1016;
wire n_103;
wire n_253;
wire n_677;
wire n_692;
wire n_951;
wire n_163;
wire n_1421;
wire n_1433;
wire n_77;
wire n_214;
wire n_167;
wire n_1134;
wire n_76;
wire n_1384;
wire n_1320;
wire n_470;
wire n_61;
wire n_216;
wire n_153;
wire n_355;
wire n_1066;
wire n_286;
wire n_408;
wire n_1003;
wire n_247;
wire n_1090;
wire n_165;
wire n_413;
wire n_1126;
wire n_1405;
wire n_290;
wire n_1031;
wire n_792;
wire n_277;
wire n_885;
wire n_631;
wire n_1410;
wire n_854;
wire n_523;
wire n_985;
wire n_901;
wire n_419;
wire n_1183;
wire n_519;
wire n_271;
wire n_1132;
wire n_785;
wire n_1137;
wire n_94;
wire n_1085;
wire n_997;
wire n_858;
wire n_1191;
wire n_58;
wire n_242;
wire n_284;
wire n_321;
wire n_811;
wire n_734;
wire n_233;
wire n_698;
wire n_257;
wire n_26;
wire n_1173;
wire n_477;
wire n_318;
wire n_1379;
wire n_98;
wire n_714;
wire n_32;
wire n_531;
wire n_406;
wire n_372;
wire n_820;
wire n_923;
wire n_702;
wire n_1301;
wire n_647;
wire n_445;
wire n_1303;
wire n_732;
wire n_926;
wire n_845;
wire n_10;
wire n_1036;
wire n_761;
wire n_1075;
wire n_510;
wire n_360;
wire n_1040;
wire n_1067;
wire n_296;
wire n_975;
wire n_89;
wire n_130;
wire n_639;
wire n_1345;
wire n_1008;
wire n_34;
wire n_395;
wire n_1392;
wire n_250;
wire n_1120;
wire n_565;
wire n_323;
wire n_1101;
wire n_1369;
wire n_1416;
wire n_1275;
wire n_240;
wire n_768;
wire n_568;
wire n_1287;
wire n_46;
wire n_174;
wire n_108;
wire n_335;
wire n_37;
wire n_515;
wire n_802;
wire n_672;
wire n_466;
wire n_87;
wire n_1027;
wire n_572;
wire n_81;
wire n_1292;
wire n_1473;
wire n_36;
wire n_917;
wire n_680;
wire n_767;
wire n_237;
wire n_1034;
wire n_633;
wire n_803;
wire n_398;
wire n_796;
wire n_1263;
wire n_1424;
wire n_662;
wire n_391;
wire n_241;
wire n_874;
wire n_449;
wire n_1070;
wire n_56;
wire n_455;
wire n_67;
wire n_401;
wire n_1159;
wire n_1434;
wire n_877;
wire n_725;
wire n_930;
wire n_1318;
wire n_1396;
wire n_1063;
wire n_291;
wire n_1233;
wire n_664;
wire n_35;
wire n_1196;
wire n_659;
wire n_968;
wire n_1093;
wire n_336;
wire n_1241;
wire n_556;
wire n_1376;
wire n_648;
wire n_60;
wire n_936;
wire n_1289;
wire n_924;
wire n_305;
wire n_1158;
wire n_358;
wire n_627;
wire n_750;
wire n_1459;
wire n_589;
wire n_128;
wire n_697;
wire n_642;
wire n_234;
wire n_848;
wire n_1005;
wire n_1153;
wire n_1361;
wire n_514;
wire n_625;
wire n_403;
wire n_995;
wire n_738;
wire n_511;
wire n_1319;
wire n_49;
wire n_1417;
wire n_646;
wire n_156;
wire n_154;
wire n_1099;
wire n_994;
wire n_1257;
wire n_204;
wire n_439;
wire n_180;
wire n_73;
wire n_1172;
wire n_74;
wire n_308;
wire n_518;
wire n_681;
wire n_189;
wire n_447;
wire n_903;
wire n_1368;
wire n_66;
wire n_379;
wire n_626;
wire n_1347;
wire n_1337;
wire n_475;
wire n_281;
wire n_1296;
wire n_516;
wire n_1282;
wire n_1389;
wire n_342;
wire n_557;
wire n_438;
wire n_1447;
wire n_461;
wire n_1382;
wire n_830;
wire n_562;
wire n_967;
wire n_526;
wire n_261;
wire n_104;
wire n_709;
wire n_1200;
wire n_821;
wire n_468;
wire n_91;
wire n_148;
wire n_378;
wire n_752;
wire n_823;
wire n_191;
wire n_63;
wire n_387;
wire n_1350;
wire n_961;
wire n_492;
wire n_1100;
wire n_1128;
wire n_219;
wire n_343;
wire n_555;
wire n_1259;
wire n_880;
wire n_312;
wire n_742;
wire n_23;
wire n_1048;
wire n_269;
wire n_751;
wire n_186;
wire n_164;
wire n_114;
wire n_1229;
wire n_50;
wire n_1322;
wire n_574;
wire n_478;
wire n_1225;
wire n_1141;
wire n_998;
wire n_1461;
wire n_824;
wire n_601;
wire n_736;
wire n_215;
wire n_172;
wire n_979;
wire n_332;
wire n_670;
wire n_1112;
wire n_755;
wire n_1193;
wire n_765;
wire n_1449;
wire n_179;
wire n_289;
wire n_721;
wire n_485;
wire n_354;
wire n_980;
wire n_70;
wire n_1399;
wire n_458;
wire n_322;
wire n_1123;
wire n_317;
wire n_800;
wire n_973;
wire n_1466;
wire n_1470;
wire n_522;
wire n_1055;
wire n_326;
wire n_532;
wire n_1206;
wire n_635;
wire n_1107;
wire n_1342;
wire n_1023;
wire n_299;
wire n_1477;
wire n_1072;
wire n_509;
wire n_1043;
wire n_263;
wire n_1230;
wire n_193;
wire n_267;
wire n_638;
wire n_873;
wire n_585;
wire n_450;
wire n_140;
wire n_779;
wire n_13;
wire n_64;
wire n_970;
wire n_921;
wire n_1373;
wire n_927;
wire n_339;
wire n_696;
wire n_748;
wire n_774;
wire n_1080;
wire n_1280;
wire n_1385;
wire n_743;
wire n_944;
wire n_96;
wire n_669;
wire n_770;
wire n_364;
wire n_33;
wire n_464;
wire n_1279;
wire n_1119;
wire n_590;
wire n_121;
wire n_161;
wire n_224;
wire n_537;
wire n_1117;
wire n_843;
wire n_85;
wire n_264;
wire n_733;
wire n_846;
wire n_791;
wire n_1334;
wire n_1157;
wire n_932;
wire n_244;
wire n_1061;
wire n_297;
wire n_350;
wire n_616;
wire n_208;
wire n_528;
wire n_168;
wire n_1271;
wire n_1011;
wire n_1087;
wire n_758;
wire n_775;
wire n_113;
wire n_498;
wire n_538;
wire n_1214;
wire n_302;
wire n_292;
wire n_547;
wire n_741;
wire n_705;
wire n_828;
wire n_1456;
wire n_988;
wire n_996;
wire n_1360;
wire n_1327;
wire n_1283;
wire n_1164;
wire n_146;
wire n_641;
wire n_93;
wire n_1294;
wire n_1472;
wire n_1332;
wire n_41;
wire n_826;
wire n_1009;
wire n_1079;
wire n_898;
wire n_417;
wire n_1215;
wire n_1192;
wire n_1248;
wire n_818;
wire n_1297;
wire n_75;
wire n_82;
wire n_183;
wire n_550;
wire n_582;
wire n_784;
wire n_170;
wire n_915;
wire n_1427;
wire n_363;
wire n_1078;
wire n_724;
wire n_1419;
wire n_21;
wire n_1148;
wire n_1380;
wire n_939;
wire n_640;
wire n_1228;
wire n_976;
wire n_1430;
wire n_938;
wire n_657;
wire n_964;
wire n_385;
wire n_227;
wire n_454;
wire n_551;
wire n_268;
wire n_190;
wire n_62;
wire n_4;
wire n_956;
wire n_781;
wire n_1071;
wire n_376;
wire n_694;
wire n_88;
wire n_807;
wire n_613;
wire n_207;
wire n_1258;
wire n_1190;
wire n_298;
wire n_630;
wire n_1395;
wire n_1290;
wire n_983;
wire n_1052;
wire n_78;
wire n_68;
wire n_919;
wire n_598;
wire n_810;
wire n_251;
wire n_916;
wire n_465;
wire n_1333;
wire n_881;
wire n_520;
wire n_668;
wire n_338;
wire n_907;
wire n_20;
wire n_782;
wire n_832;
wire n_790;
wire n_504;
wire n_456;
wire n_319;
wire n_1328;
wire n_1227;
wire n_933;
wire n_719;
wire n_788;
wire n_655;
wire n_1208;
wire n_1103;
wire n_472;
wire n_1142;
wire n_1010;
wire n_457;
wire n_1346;
wire n_255;
wire n_1170;
wire n_513;
wire n_29;
wire n_893;
wire n_382;
wire n_894;
wire n_536;
wire n_474;
wire n_1387;
wire n_745;
wire n_706;
wire n_1370;
wire n_1165;
wire n_1210;
wire n_958;
wire n_0;
wire n_619;
wire n_258;
wire n_974;
wire n_1155;
wire n_607;
wire n_184;
wire n_1251;
wire n_1453;
wire n_144;
wire n_1130;
wire n_420;
wire n_1341;
wire n_86;
wire n_28;
wire n_206;
wire n_1362;
wire n_349;
wire n_673;
wire n_1124;
wire n_1364;
wire n_25;
wire n_592;
wire n_1238;
wire n_545;
wire n_99;
wire n_43;
wire n_199;
wire n_1184;
wire n_1340;
wire n_831;
wire n_1295;
wire n_729;
wire n_394;
wire n_44;
wire n_352;
wire n_689;
wire n_1268;
wire n_1306;
wire n_316;
wire n_586;
wire n_1388;
wire n_1252;
wire n_1131;
wire n_1426;
wire n_645;
wire n_497;
wire n_11;
wire n_1314;
wire n_1088;
wire n_1242;
wire n_1197;
wire n_805;
wire n_1315;
wire n_373;
wire n_753;
wire n_71;
wire n_288;
wire n_176;
wire n_931;
wire n_195;
wire n_1400;
wire n_723;
wire n_833;
wire n_1281;
wire n_409;
wire n_838;
wire n_534;
wire n_423;
wire n_483;
wire n_353;
wire n_303;
wire n_1187;
wire n_566;
wire n_149;
wire n_567;
wire n_1435;
wire n_780;
wire n_1224;
wire n_864;
wire n_125;
wire n_596;
wire n_1046;
wire n_1111;
wire n_1243;
wire n_494;
wire n_1115;
wire n_135;
wire n_481;
wire n_1147;
wire n_127;
wire n_182;
wire n_529;
wire n_656;
wire n_1246;
wire n_1397;
wire n_1226;
wire n_137;
wire n_1274;
wire n_651;
wire n_882;
wire n_999;
wire n_636;
wire n_614;
wire n_737;
wire n_1391;
wire n_428;
wire n_178;
wire n_1276;
wire n_708;
wire n_229;
wire n_442;
wire n_1176;
wire n_1348;
wire n_699;
wire n_857;
wire n_1273;
wire n_1199;
wire n_8;
wire n_1185;
wire n_578;
wire n_928;
wire n_187;
wire n_188;
wire n_18;
wire n_628;
wire n_425;
wire n_905;
wire n_109;
wire n_198;
wire n_1310;
wire n_426;
wire n_716;
wire n_892;
wire n_115;
wire n_476;
wire n_989;
wire n_599;
wire n_1232;
wire n_715;
wire n_849;
wire n_1077;
wire n_404;
wire n_1288;
wire n_362;
wire n_688;
wire n_1428;
wire n_152;
wire n_1475;
wire n_1102;
wire n_1177;
wire n_506;
wire n_328;
wire n_1305;
wire n_1411;
wire n_388;
wire n_1260;
wire n_763;
wire n_632;
wire n_906;
wire n_615;
wire n_1145;
wire n_701;
wire n_1335;
wire n_888;
wire n_661;
wire n_909;
wire n_493;
wire n_972;
wire n_690;
wire n_272;
wire n_1442;
wire n_561;
wire n_1413;
wire n_1057;
wire n_581;
wire n_280;
wire n_1068;
wire n_1352;
wire n_377;
wire n_1044;
wire n_1013;
wire n_1143;
wire n_185;
wire n_955;
wire n_1007;
wire n_950;
wire n_171;
wire n_899;
wire n_111;
wire n_978;
wire n_30;
wire n_634;
wire n_1444;
wire n_559;
wire n_407;
wire n_527;
wire n_200;
wire n_986;
wire n_262;
wire n_1349;
wire n_503;
wire n_969;
wire n_1138;
wire n_856;
wire n_1081;
wire n_347;
wire n_79;
wire n_1265;
wire n_1284;
wire n_521;
wire n_157;
wire n_808;
wire n_1113;
wire n_1038;
wire n_434;
wire n_624;
wire n_1240;
wire n_273;
wire n_571;
wire n_325;
wire n_524;
wire n_1118;
wire n_1420;
wire n_530;
wire n_348;
wire n_762;
wire n_685;
wire n_90;
wire n_72;
wire n_594;
wire n_1114;
wire n_1030;
wire n_1253;
wire n_861;
wire n_809;
wire n_908;
wire n_1239;
wire n_1022;
wire n_463;
wire n_1125;
wire n_484;
wire n_431;
wire n_860;
wire n_710;
wire n_560;
wire n_525;
wire n_1174;
wire n_393;
wire n_211;
wire n_283;
wire n_1406;
wire n_217;
wire n_1264;
wire n_259;
wire n_1178;
wire n_666;
wire n_276;
wire n_225;
wire n_815;
wire n_922;
wire n_839;
wire n_1403;
wire n_1109;
wire n_739;
wire n_1221;
wire n_1356;
wire n_501;
wire n_1443;
wire n_1414;
wire n_1330;
wire n_593;
wire n_597;
wire n_1097;
wire n_1234;
wire n_1151;
wire n_203;
wire n_460;
wire n_1458;
wire n_1235;
wire n_637;
wire n_957;
wire n_872;
wire n_539;
wire n_713;
wire n_467;
wire n_760;
wire n_665;
wire n_1436;
wire n_390;
wire n_1001;
wire n_1161;
wire n_1321;
wire n_778;
wire n_1393;
wire n_925;
wire n_158;
wire n_249;
wire n_749;
wire n_1069;
wire n_1098;
wire n_106;
wire n_605;
wire n_835;
wire n_437;
wire n_940;
wire n_1150;
wire n_700;
wire n_1033;
wire n_1381;
wire n_1236;
wire n_822;
wire n_381;
wire n_142;
wire n_754;
wire n_453;
wire n_59;
wire n_1121;
wire n_914;
wire n_945;
wire n_852;
wire n_1336;
wire n_122;
wire n_374;
wire n_1042;
wire n_197;
wire n_541;
wire n_1285;
wire n_112;
wire n_735;
wire n_552;
wire n_1323;
wire n_962;
wire n_1422;
wire n_416;
wire n_1299;
wire n_1205;
wire n_414;
wire n_469;
wire n_1313;
wire n_1331;
wire n_429;
wire n_1270;
wire n_804;
wire n_1460;
wire n_117;
wire n_577;
wire n_238;
wire n_294;
wire n_2;
wire n_1256;
wire n_618;
wire n_412;
wire n_22;
wire n_683;
wire n_479;
wire n_1266;
wire n_584;
wire n_311;
wire n_813;
wire n_819;
wire n_1096;
wire n_39;
wire n_953;
wire n_489;
wire n_245;
wire n_764;
wire n_486;
wire n_794;
wire n_1261;
wire n_1343;
wire n_1394;
wire n_1017;
wire n_1195;
wire n_1291;
wire n_543;
wire n_218;
wire n_173;
wire n_488;
wire n_1105;
wire n_799;
wire n_937;
wire n_462;
wire n_495;
wire n_430;
wire n_418;
wire n_175;
wire n_897;
wire n_512;
wire n_1188;
wire n_265;
wire n_57;
wire n_51;
wire n_1465;
wire n_1231;
wire n_131;
wire n_27;
wire n_1180;
wire n_1365;
wire n_448;
wire n_415;
wire n_31;
wire n_1309;
wire n_1432;
wire n_239;
wire n_7;
wire n_895;
wire n_1029;
wire n_1014;
wire n_929;
wire n_769;
wire n_370;
wire n_1015;
wire n_604;
wire n_440;
wire n_1375;
wire n_786;
wire n_1249;
wire n_1359;
wire n_1425;
wire n_226;
wire n_535;
wire n_1116;
wire n_285;
wire n_564;
wire n_1047;
wire n_471;
wire n_1049;
wire n_949;
wire n_1035;
wire n_1104;
wire n_371;
wire n_579;
wire n_608;
wire n_368;
wire n_1020;
wire n_859;
wire n_1438;
wire n_223;
wire n_1440;
wire n_19;
wire n_1372;
wire n_971;
wire n_569;
wire n_410;
wire n_502;
wire n_1262;
wire n_1312;
wire n_1462;
wire n_1136;
wire n_1298;
wire n_629;
wire n_1189;
wire n_558;
wire n_181;
wire n_123;
wire n_553;
wire n_1398;
wire n_817;
wire n_776;
wire n_397;
wire n_315;
wire n_53;
wire n_1476;
wire n_1201;
wire n_1058;
wire n_836;
wire n_293;
wire n_1439;
wire n_1028;
wire n_990;
wire n_663;
wire n_1338;
wire n_887;
wire n_507;
wire n_334;
wire n_1095;
wire n_1062;
wire n_993;
wire n_806;
wire n_120;
wire n_1053;
wire n_650;
wire n_1378;
wire n_162;
wire n_977;
wire n_772;
wire n_816;
wire n_789;
wire n_1255;
wire n_3;
wire n_884;
wire n_330;
wire n_231;
wire n_1307;
wire n_9;
wire n_1211;
wire n_1404;
wire n_1083;
wire n_652;
wire n_97;
wire n_982;
wire n_324;
wire n_422;
wire n_192;
wire n_329;
wire n_1409;
wire n_6;
wire n_1383;
wire n_1293;
wire n_1160;
wire n_883;
wire n_801;
wire n_912;
wire n_314;
wire n_307;
wire n_934;
wire n_16;
wire n_95;
wire n_40;
wire n_210;
wire n_1371;
wire n_228;
wire n_863;
wire n_671;
wire n_1144;
wire n_278;
wire n_270;
wire n_1135;
wire n_1415;
wire n_617;
wire n_396;
wire n_1139;
wire n_851;
wire n_588;
wire n_375;
wire n_1162;
wire n_855;
wire n_911;
wire n_491;
wire n_1216;
wire n_1329;
wire n_80;
wire n_1237;
wire n_546;
wire n_756;
wire n_1437;
wire n_992;
wire n_576;
wire n_1366;
wire n_1351;
wire n_622;
wire n_910;
wire n_150;
wire n_235;
wire n_533;
wire n_686;
wire n_1269;
wire n_141;
wire n_160;
wire n_1182;
wire n_499;
wire n_1377;
wire n_757;
wire n_1429;
wire n_1060;
wire n_232;
wire n_812;
wire n_783;
wire n_147;
wire n_1065;
wire n_644;
wire n_1326;
wire n_746;
wire n_1064;
wire n_1358;
wire n_1441;
wire n_583;
wire n_1408;
wire n_248;
wire n_866;
wire n_1457;
wire n_83;
wire n_1106;
wire n_603;
wire n_1032;
wire n_119;
wire n_667;
wire n_1076;
wire n_1018;
wire n_129;
wire n_611;
wire n_421;
wire n_52;
wire n_1179;
wire n_850;
wire n_1308;
wire n_1074;
wire n_787;
wire n_1390;
wire n_1272;
wire n_1108;
wire n_609;
wire n_946;
wire n_1082;
wire n_65;
wire n_5;
wire n_496;
wire n_1181;
wire n_1316;
wire n_320;
wire n_102;
wire n_201;
wire n_1363;
wire n_612;
wire n_771;
wire n_827;
wire n_1037;
wire n_747;
wire n_252;
wire n_966;
wire n_693;
wire n_896;
wire n_1212;
wire n_1056;
wire n_194;
wire n_825;
wire n_282;
wire n_1223;
wire n_703;
wire n_1254;
wire n_116;
wire n_1213;
wire n_1247;
wire n_118;
wire n_587;
wire n_554;
wire n_722;
wire n_1245;
wire n_1357;
wire n_243;
wire n_346;
wire n_1154;
wire n_345;
wire n_230;
wire n_452;
wire n_1455;
wire n_337;
wire n_726;
wire n_847;
wire n_842;
wire n_918;
wire n_623;
wire n_451;
wire n_500;
wire n_948;
wire n_1026;
wire n_575;
wire n_600;
wire n_731;
wire n_1006;
wire n_132;
wire n_643;
wire n_1418;
wire n_205;
wire n_126;
wire n_473;
wire n_389;
wire n_834;
wire n_427;
wire n_1194;
wire n_42;
wire n_1086;
wire n_871;
wire n_620;
wire n_480;
wire n_1073;
wire n_1039;
wire n_341;
wire n_310;
wire n_14;
wire n_236;
wire n_727;
wire n_136;
wire n_260;
wire n_891;
wire n_1317;
wire n_1002;
wire n_1004;
wire n_580;
wire n_610;
wire n_222;
wire n_1302;
wire n_853;
wire n_1325;
wire n_798;
wire n_943;
wire n_606;
wire n_1353;
wire n_712;
wire n_777;
wire n_954;
wire n_902;
wire n_459;
wire n_1446;
wire n_717;
wire n_865;
wire n_380;
wire n_867;
wire n_649;
wire n_602;
wire n_1355;
wire n_444;
wire n_105;
wire n_1220;
wire n_889;
wire n_870;
wire n_432;
wire n_913;
wire n_730;
wire n_369;
wire n_1146;
wire n_361;
wire n_1354;
wire n_1163;
wire n_654;
wire n_15;
wire n_960;
wire n_256;
wire n_365;
wire n_1469;
wire n_1222;
wire n_591;
wire n_1025;
wire n_209;
wire n_84;
wire n_12;
wire n_1133;
wire n_1250;
wire n_1169;
wire n_383;
wire n_202;
wire n_542;
wire n_862;
wire n_101;
wire n_1168;
wire n_941;
wire n_1304;
wire n_508;
wire n_24;
wire n_1204;
wire n_490;
wire n_540;
wire n_947;
wire n_840;
wire n_400;
wire n_1094;
wire n_134;
wire n_48;
wire n_563;
wire n_1339;
wire n_55;
wire n_718;
wire n_1140;
wire n_1156;
wire n_138;
wire n_573;
wire n_505;
wire n_740;
wire n_313;
wire n_92;
wire n_333;
wire n_306;
wire n_1344;
wire n_675;
wire n_1431;
wire n_1219;
wire n_1000;
wire n_674;
wire n_570;
wire n_411;
wire n_287;
wire n_45;
wire n_1217;
wire n_177;
wire n_1054;
wire n_1166;
wire n_436;
wire n_1051;
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_269), .Y(n_361) );
BUFx10_ASAP7_75t_L g362 ( .A(n_351), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_317), .Y(n_363) );
INVx2_ASAP7_75t_SL g364 ( .A(n_339), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_137), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_32), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_262), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_279), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_204), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_22), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_203), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_358), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_206), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_3), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_34), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_85), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_135), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_169), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_16), .Y(n_379) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_343), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_113), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_266), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_243), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_10), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_175), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_94), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_222), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_104), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_312), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_106), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_12), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_21), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_54), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_102), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_199), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_354), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_313), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_261), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_333), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_360), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_256), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_88), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_85), .Y(n_403) );
INVx4_ASAP7_75t_R g404 ( .A(n_284), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_291), .Y(n_405) );
INVxp33_ASAP7_75t_SL g406 ( .A(n_37), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_210), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_249), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_124), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_48), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_278), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_240), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_157), .Y(n_413) );
INVxp33_ASAP7_75t_L g414 ( .A(n_346), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_109), .Y(n_415) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_232), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_42), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_77), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_246), .Y(n_419) );
BUFx3_ASAP7_75t_L g420 ( .A(n_331), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_200), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_11), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_344), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_301), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_160), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_178), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_213), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_188), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_28), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_171), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_117), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_233), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_318), .Y(n_433) );
INVxp33_ASAP7_75t_L g434 ( .A(n_139), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_181), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_242), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_123), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_326), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_248), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_134), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_226), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_270), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_359), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_253), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_352), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_66), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_202), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_221), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_286), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_143), .Y(n_450) );
BUFx10_ASAP7_75t_L g451 ( .A(n_309), .Y(n_451) );
INVxp33_ASAP7_75t_L g452 ( .A(n_36), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_349), .Y(n_453) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_23), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_35), .Y(n_455) );
BUFx5_ASAP7_75t_L g456 ( .A(n_111), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_276), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_5), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_115), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_258), .Y(n_460) );
BUFx3_ASAP7_75t_L g461 ( .A(n_329), .Y(n_461) );
INVxp33_ASAP7_75t_SL g462 ( .A(n_274), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_308), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_225), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_19), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_158), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_357), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_214), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_25), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_350), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_79), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_337), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_145), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_323), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_234), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_155), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_142), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_23), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_90), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_310), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_32), .Y(n_481) );
INVxp33_ASAP7_75t_SL g482 ( .A(n_194), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_186), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_110), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_47), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_132), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_25), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_97), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_150), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_219), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_119), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_59), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_68), .B(n_12), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_275), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_320), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_104), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_292), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_324), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_67), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_207), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_151), .Y(n_501) );
INVxp33_ASAP7_75t_SL g502 ( .A(n_102), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_106), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_16), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_78), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_296), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_133), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_96), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_91), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_154), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_280), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_68), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_250), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_138), .Y(n_514) );
INVxp33_ASAP7_75t_L g515 ( .A(n_103), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_172), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_267), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_216), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_128), .Y(n_519) );
NOR2xp67_ASAP7_75t_L g520 ( .A(n_183), .B(n_170), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_11), .Y(n_521) );
BUFx3_ASAP7_75t_L g522 ( .A(n_231), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_263), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_341), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_76), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_227), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_27), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_152), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_305), .Y(n_529) );
BUFx3_ASAP7_75t_L g530 ( .A(n_153), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_126), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_332), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_265), .Y(n_533) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_247), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_239), .B(n_140), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_1), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_277), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_8), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_65), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_141), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_81), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_345), .B(n_281), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_114), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_507), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_376), .B(n_0), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_507), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_527), .B(n_449), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_499), .B(n_0), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_475), .Y(n_549) );
BUFx3_ASAP7_75t_L g550 ( .A(n_420), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_365), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_365), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_365), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_431), .B(n_1), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_456), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_365), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_380), .Y(n_557) );
INVx3_ASAP7_75t_L g558 ( .A(n_362), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_456), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_456), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_456), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_380), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_411), .B(n_2), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_406), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_380), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_380), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_456), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_456), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_468), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_378), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_375), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_468), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_375), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_459), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_361), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_378), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_383), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_362), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_468), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_459), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_499), .Y(n_581) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_468), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_363), .Y(n_583) );
AND2x6_ASAP7_75t_L g584 ( .A(n_420), .B(n_120), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_583), .B(n_364), .Y(n_585) );
AO22x1_ASAP7_75t_L g586 ( .A1(n_584), .A2(n_414), .B1(n_434), .B2(n_462), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_548), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_555), .Y(n_588) );
INVx3_ASAP7_75t_L g589 ( .A(n_548), .Y(n_589) );
INVx5_ASAP7_75t_L g590 ( .A(n_584), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_558), .B(n_414), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_583), .B(n_474), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_558), .B(n_452), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_558), .B(n_537), .Y(n_594) );
BUFx3_ASAP7_75t_L g595 ( .A(n_550), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_558), .B(n_366), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_555), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_559), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_547), .B(n_454), .Y(n_599) );
NAND2xp33_ASAP7_75t_L g600 ( .A(n_584), .B(n_368), .Y(n_600) );
OAI22xp33_ASAP7_75t_L g601 ( .A1(n_564), .A2(n_479), .B1(n_515), .B2(n_452), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_559), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_578), .B(n_581), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_578), .B(n_374), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_552), .Y(n_605) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_548), .B(n_542), .Y(n_606) );
INVx2_ASAP7_75t_SL g607 ( .A(n_550), .Y(n_607) );
BUFx3_ASAP7_75t_L g608 ( .A(n_550), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_560), .Y(n_609) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_552), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_578), .B(n_515), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_548), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_578), .B(n_362), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_584), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_552), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_549), .B(n_451), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_552), .Y(n_617) );
INVx4_ASAP7_75t_L g618 ( .A(n_584), .Y(n_618) );
BUFx3_ASAP7_75t_L g619 ( .A(n_584), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_552), .Y(n_620) );
BUFx3_ASAP7_75t_L g621 ( .A(n_584), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_560), .Y(n_622) );
INVx4_ASAP7_75t_SL g623 ( .A(n_584), .Y(n_623) );
INVx3_ASAP7_75t_L g624 ( .A(n_544), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_544), .B(n_434), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_561), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_544), .B(n_451), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_570), .A2(n_381), .B1(n_384), .B2(n_379), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_546), .B(n_451), .Y(n_629) );
AND3x4_ASAP7_75t_L g630 ( .A(n_570), .B(n_520), .C(n_502), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_624), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_624), .Y(n_632) );
BUFx3_ASAP7_75t_L g633 ( .A(n_595), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_593), .Y(n_634) );
BUFx3_ASAP7_75t_L g635 ( .A(n_595), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_624), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_591), .B(n_563), .Y(n_637) );
NOR2xp33_ASAP7_75t_R g638 ( .A(n_600), .B(n_575), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_612), .A2(n_502), .B1(n_406), .B2(n_581), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_624), .Y(n_640) );
NAND2x1p5_ASAP7_75t_L g641 ( .A(n_627), .B(n_493), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_612), .A2(n_545), .B1(n_567), .B2(n_561), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_630), .A2(n_568), .B1(n_567), .B2(n_482), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_593), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_627), .B(n_554), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_611), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_630), .A2(n_400), .B1(n_408), .B2(n_361), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_611), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_629), .B(n_546), .Y(n_649) );
BUFx3_ASAP7_75t_L g650 ( .A(n_595), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_629), .B(n_546), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_629), .B(n_462), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_618), .B(n_568), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_625), .B(n_571), .Y(n_654) );
AOI21xp33_ASAP7_75t_L g655 ( .A1(n_599), .A2(n_611), .B(n_594), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_596), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_596), .B(n_571), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_594), .B(n_514), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_596), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_613), .B(n_573), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_596), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_587), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g663 ( .A(n_630), .B(n_408), .C(n_400), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_606), .A2(n_494), .B1(n_501), .B2(n_426), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_618), .B(n_367), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_592), .B(n_573), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_587), .Y(n_667) );
INVx3_ASAP7_75t_L g668 ( .A(n_587), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_587), .A2(n_388), .B1(n_390), .B2(n_386), .Y(n_669) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_619), .Y(n_670) );
NOR2xp33_ASAP7_75t_SL g671 ( .A(n_618), .B(n_426), .Y(n_671) );
INVx3_ASAP7_75t_L g672 ( .A(n_589), .Y(n_672) );
BUFx2_ASAP7_75t_L g673 ( .A(n_599), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_604), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_592), .B(n_418), .Y(n_675) );
INVx4_ASAP7_75t_L g676 ( .A(n_623), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_599), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_588), .A2(n_371), .B(n_369), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_606), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_606), .A2(n_501), .B1(n_516), .B2(n_494), .Y(n_680) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_619), .Y(n_681) );
AND2x4_ASAP7_75t_L g682 ( .A(n_604), .B(n_574), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_604), .Y(n_683) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_619), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_604), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_589), .Y(n_686) );
BUFx10_ASAP7_75t_L g687 ( .A(n_604), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_589), .A2(n_422), .B1(n_429), .B2(n_391), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_588), .A2(n_373), .B(n_372), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_616), .B(n_603), .Y(n_690) );
BUFx3_ASAP7_75t_L g691 ( .A(n_608), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_606), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_603), .B(n_574), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_589), .B(n_580), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g695 ( .A(n_586), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_601), .B(n_418), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_618), .B(n_377), .Y(n_697) );
NOR2xp67_ASAP7_75t_L g698 ( .A(n_585), .B(n_576), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_590), .B(n_387), .Y(n_699) );
NAND2xp33_ASAP7_75t_L g700 ( .A(n_590), .B(n_382), .Y(n_700) );
AO22x1_ASAP7_75t_L g701 ( .A1(n_586), .A2(n_543), .B1(n_541), .B2(n_417), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_585), .B(n_580), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_597), .A2(n_397), .B(n_396), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_597), .Y(n_704) );
NOR2x2_ASAP7_75t_L g705 ( .A(n_628), .B(n_370), .Y(n_705) );
INVx2_ASAP7_75t_SL g706 ( .A(n_590), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_608), .B(n_389), .Y(n_707) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_628), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_623), .B(n_543), .Y(n_709) );
CKINVDCx5p33_ASAP7_75t_R g710 ( .A(n_621), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_608), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_598), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_598), .B(n_413), .Y(n_713) );
OAI21x1_ASAP7_75t_L g714 ( .A1(n_704), .A2(n_609), .B(n_602), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_664), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_712), .A2(n_609), .B(n_622), .C(n_602), .Y(n_716) );
AND2x4_ASAP7_75t_L g717 ( .A(n_634), .B(n_623), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_656), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_668), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_675), .B(n_626), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_673), .B(n_402), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_668), .Y(n_722) );
AO32x2_ASAP7_75t_L g723 ( .A1(n_679), .A2(n_607), .A3(n_614), .B1(n_577), .B2(n_576), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_668), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_659), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_672), .Y(n_726) );
INVxp67_ASAP7_75t_L g727 ( .A(n_680), .Y(n_727) );
BUFx4f_ASAP7_75t_L g728 ( .A(n_641), .Y(n_728) );
BUFx2_ASAP7_75t_L g729 ( .A(n_692), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_653), .A2(n_614), .B(n_621), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_708), .A2(n_528), .B1(n_626), .B2(n_622), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_661), .Y(n_732) );
BUFx3_ASAP7_75t_L g733 ( .A(n_641), .Y(n_733) );
INVx5_ASAP7_75t_L g734 ( .A(n_687), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_644), .B(n_623), .Y(n_735) );
O2A1O1Ixp33_ASAP7_75t_L g736 ( .A1(n_655), .A2(n_410), .B(n_455), .C(n_446), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_674), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_672), .Y(n_738) );
OR2x6_ASAP7_75t_L g739 ( .A(n_679), .B(n_458), .Y(n_739) );
BUFx2_ASAP7_75t_L g740 ( .A(n_705), .Y(n_740) );
INVx2_ASAP7_75t_SL g741 ( .A(n_675), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_645), .B(n_607), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_646), .B(n_623), .Y(n_743) );
O2A1O1Ixp5_ASAP7_75t_SL g744 ( .A1(n_678), .A2(n_399), .B(n_401), .C(n_398), .Y(n_744) );
INVx4_ASAP7_75t_L g745 ( .A(n_687), .Y(n_745) );
AND2x4_ASAP7_75t_L g746 ( .A(n_648), .B(n_623), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_672), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_687), .Y(n_748) );
BUFx4f_ASAP7_75t_SL g749 ( .A(n_696), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_L g750 ( .A1(n_696), .A2(n_469), .B(n_478), .C(n_465), .Y(n_750) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_670), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_SL g752 ( .A1(n_690), .A2(n_577), .B(n_535), .C(n_553), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_683), .Y(n_753) );
BUFx8_ASAP7_75t_SL g754 ( .A(n_677), .Y(n_754) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_670), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_662), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_665), .A2(n_590), .B(n_534), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_708), .A2(n_392), .B1(n_393), .B2(n_370), .Y(n_758) );
BUFx2_ASAP7_75t_L g759 ( .A(n_705), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_662), .Y(n_760) );
AND2x4_ASAP7_75t_L g761 ( .A(n_657), .B(n_484), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_685), .Y(n_762) );
A2O1A1Ixp33_ASAP7_75t_L g763 ( .A1(n_637), .A2(n_487), .B(n_488), .C(n_485), .Y(n_763) );
O2A1O1Ixp33_ASAP7_75t_L g764 ( .A1(n_649), .A2(n_492), .B(n_496), .C(n_491), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_694), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_638), .Y(n_766) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_670), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_665), .A2(n_590), .B(n_416), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_694), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_667), .Y(n_770) );
BUFx3_ASAP7_75t_L g771 ( .A(n_657), .Y(n_771) );
BUFx4f_ASAP7_75t_L g772 ( .A(n_657), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_647), .Y(n_773) );
BUFx4f_ASAP7_75t_L g774 ( .A(n_682), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_667), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_643), .A2(n_393), .B1(n_394), .B2(n_392), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_697), .A2(n_590), .B(n_407), .Y(n_777) );
BUFx6f_ASAP7_75t_L g778 ( .A(n_670), .Y(n_778) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_701), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_697), .A2(n_590), .B(n_409), .Y(n_780) );
AOI21x1_ASAP7_75t_L g781 ( .A1(n_699), .A2(n_615), .B(n_605), .Y(n_781) );
INVx1_ASAP7_75t_SL g782 ( .A(n_709), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_694), .Y(n_783) );
BUFx2_ASAP7_75t_L g784 ( .A(n_709), .Y(n_784) );
NAND2xp5_ASAP7_75t_SL g785 ( .A(n_671), .B(n_590), .Y(n_785) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_681), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_652), .B(n_403), .Y(n_787) );
CKINVDCx11_ASAP7_75t_R g788 ( .A(n_682), .Y(n_788) );
INVx3_ASAP7_75t_L g789 ( .A(n_682), .Y(n_789) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_698), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_663), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_666), .B(n_471), .Y(n_792) );
BUFx3_ASAP7_75t_L g793 ( .A(n_631), .Y(n_793) );
NOR2xp33_ASAP7_75t_SL g794 ( .A(n_676), .B(n_481), .Y(n_794) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_681), .Y(n_795) );
OR2x6_ASAP7_75t_L g796 ( .A(n_651), .B(n_504), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_695), .A2(n_503), .B1(n_521), .B2(n_512), .Y(n_797) );
INVx1_ASAP7_75t_SL g798 ( .A(n_633), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_686), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_686), .Y(n_800) );
CKINVDCx8_ASAP7_75t_R g801 ( .A(n_660), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_658), .A2(n_639), .B1(n_642), .B2(n_669), .Y(n_802) );
OAI22xp5_ASAP7_75t_SL g803 ( .A1(n_688), .A2(n_508), .B1(n_509), .B2(n_505), .Y(n_803) );
OAI21xp33_ASAP7_75t_L g804 ( .A1(n_654), .A2(n_536), .B(n_525), .Y(n_804) );
INVx4_ASAP7_75t_L g805 ( .A(n_676), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_711), .Y(n_806) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_681), .Y(n_807) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_681), .Y(n_808) );
HB1xp67_ASAP7_75t_SL g809 ( .A(n_676), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_711), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_693), .A2(n_539), .B1(n_538), .B2(n_419), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_633), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g813 ( .A1(n_702), .A2(n_415), .B1(n_448), .B2(n_436), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_631), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_635), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_689), .A2(n_415), .B1(n_421), .B2(n_405), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_703), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g818 ( .A1(n_713), .A2(n_425), .B(n_424), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_635), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_632), .B(n_427), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_632), .B(n_428), .Y(n_821) );
NAND2x1p5_ASAP7_75t_L g822 ( .A(n_650), .B(n_415), .Y(n_822) );
BUFx8_ASAP7_75t_SL g823 ( .A(n_636), .Y(n_823) );
NAND2xp5_ASAP7_75t_SL g824 ( .A(n_710), .B(n_460), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_650), .Y(n_825) );
OAI21x1_ASAP7_75t_SL g826 ( .A1(n_707), .A2(n_385), .B(n_383), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_636), .B(n_415), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_640), .B(n_430), .Y(n_828) );
NAND2xp33_ASAP7_75t_L g829 ( .A(n_710), .B(n_467), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_691), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_691), .A2(n_435), .B1(n_437), .B2(n_432), .Y(n_831) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_684), .Y(n_832) );
O2A1O1Ixp5_ASAP7_75t_SL g833 ( .A1(n_699), .A2(n_438), .B(n_440), .C(n_439), .Y(n_833) );
BUFx2_ASAP7_75t_L g834 ( .A(n_684), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_684), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_684), .Y(n_836) );
INVx2_ASAP7_75t_SL g837 ( .A(n_706), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_706), .B(n_441), .Y(n_838) );
NAND2xp5_ASAP7_75t_SL g839 ( .A(n_700), .B(n_480), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_700), .Y(n_840) );
BUFx6f_ASAP7_75t_L g841 ( .A(n_679), .Y(n_841) );
INVx3_ASAP7_75t_L g842 ( .A(n_687), .Y(n_842) );
INVx3_ASAP7_75t_L g843 ( .A(n_687), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_675), .B(n_442), .Y(n_844) );
OAI21x1_ASAP7_75t_L g845 ( .A1(n_714), .A2(n_395), .B(n_385), .Y(n_845) );
AOI21x1_ASAP7_75t_L g846 ( .A1(n_826), .A2(n_412), .B(n_395), .Y(n_846) );
OAI22xp33_ASAP7_75t_L g847 ( .A1(n_794), .A2(n_464), .B1(n_518), .B2(n_461), .Y(n_847) );
OAI21x1_ASAP7_75t_L g848 ( .A1(n_781), .A2(n_423), .B(n_412), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_741), .A2(n_444), .B1(n_445), .B2(n_443), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_756), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_760), .Y(n_851) );
OAI21x1_ASAP7_75t_L g852 ( .A1(n_822), .A2(n_433), .B(n_423), .Y(n_852) );
INVx3_ASAP7_75t_SL g853 ( .A(n_739), .Y(n_853) );
OAI21xp5_ASAP7_75t_L g854 ( .A1(n_744), .A2(n_450), .B(n_447), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_770), .Y(n_855) );
BUFx12f_ASAP7_75t_L g856 ( .A(n_788), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_761), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_720), .B(n_453), .Y(n_858) );
BUFx6f_ASAP7_75t_L g859 ( .A(n_841), .Y(n_859) );
OAI21x1_ASAP7_75t_L g860 ( .A1(n_822), .A2(n_526), .B(n_433), .Y(n_860) );
A2O1A1Ixp33_ASAP7_75t_SL g861 ( .A1(n_736), .A2(n_535), .B(n_553), .C(n_551), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_792), .B(n_728), .Y(n_862) );
CKINVDCx12_ASAP7_75t_R g863 ( .A(n_739), .Y(n_863) );
OR2x2_ASAP7_75t_L g864 ( .A(n_758), .B(n_4), .Y(n_864) );
BUFx3_ASAP7_75t_L g865 ( .A(n_734), .Y(n_865) );
A2O1A1Ixp33_ASAP7_75t_L g866 ( .A1(n_720), .A2(n_526), .B(n_463), .C(n_466), .Y(n_866) );
INVx2_ASAP7_75t_SL g867 ( .A(n_728), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_733), .B(n_5), .Y(n_868) );
AO21x1_ASAP7_75t_L g869 ( .A1(n_840), .A2(n_470), .B(n_457), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_754), .Y(n_870) );
NOR2x1_ASAP7_75t_SL g871 ( .A(n_739), .B(n_461), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_775), .Y(n_872) );
AND2x2_ASAP7_75t_SL g873 ( .A(n_794), .B(n_472), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_823), .Y(n_874) );
OR2x2_ASAP7_75t_L g875 ( .A(n_758), .B(n_6), .Y(n_875) );
BUFx3_ASAP7_75t_L g876 ( .A(n_734), .Y(n_876) );
OAI21x1_ASAP7_75t_L g877 ( .A1(n_833), .A2(n_476), .B(n_473), .Y(n_877) );
OAI21x1_ASAP7_75t_L g878 ( .A1(n_820), .A2(n_483), .B(n_477), .Y(n_878) );
AND2x4_ASAP7_75t_L g879 ( .A(n_734), .B(n_486), .Y(n_879) );
OAI21x1_ASAP7_75t_L g880 ( .A1(n_820), .A2(n_490), .B(n_489), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_796), .Y(n_881) );
OAI21x1_ASAP7_75t_L g882 ( .A1(n_821), .A2(n_497), .B(n_495), .Y(n_882) );
A2O1A1Ixp33_ASAP7_75t_L g883 ( .A1(n_764), .A2(n_498), .B(n_506), .C(n_500), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_817), .B(n_510), .Y(n_884) );
AO21x2_ASAP7_75t_L g885 ( .A1(n_752), .A2(n_513), .B(n_511), .Y(n_885) );
OA21x2_ASAP7_75t_L g886 ( .A1(n_821), .A2(n_519), .B(n_517), .Y(n_886) );
AND2x4_ASAP7_75t_L g887 ( .A(n_745), .B(n_524), .Y(n_887) );
OAI21xp5_ASAP7_75t_L g888 ( .A1(n_716), .A2(n_531), .B(n_529), .Y(n_888) );
INVx2_ASAP7_75t_L g889 ( .A(n_800), .Y(n_889) );
OAI21x1_ASAP7_75t_L g890 ( .A1(n_828), .A2(n_540), .B(n_532), .Y(n_890) );
AND2x4_ASAP7_75t_L g891 ( .A(n_745), .B(n_464), .Y(n_891) );
AOI22x1_ASAP7_75t_L g892 ( .A1(n_818), .A2(n_553), .B1(n_556), .B2(n_551), .Y(n_892) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_729), .Y(n_893) );
A2O1A1Ixp33_ASAP7_75t_L g894 ( .A1(n_804), .A2(n_518), .B(n_530), .C(n_522), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_731), .A2(n_533), .B1(n_523), .B2(n_530), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_802), .B(n_727), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_718), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_844), .B(n_6), .Y(n_898) );
INVx6_ASAP7_75t_L g899 ( .A(n_841), .Y(n_899) );
OR2x2_ASAP7_75t_L g900 ( .A(n_721), .B(n_7), .Y(n_900) );
AOI21xp5_ASAP7_75t_L g901 ( .A1(n_838), .A2(n_615), .B(n_605), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_725), .Y(n_902) );
AO21x2_ASAP7_75t_L g903 ( .A1(n_838), .A2(n_556), .B(n_551), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_844), .B(n_9), .Y(n_904) );
OAI21x1_ASAP7_75t_L g905 ( .A1(n_743), .A2(n_617), .B(n_562), .Y(n_905) );
NOR2x1_ASAP7_75t_SL g906 ( .A(n_841), .B(n_522), .Y(n_906) );
OA21x2_ASAP7_75t_L g907 ( .A1(n_816), .A2(n_617), .B(n_562), .Y(n_907) );
OAI21x1_ASAP7_75t_L g908 ( .A1(n_836), .A2(n_617), .B(n_562), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_789), .B(n_9), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_782), .A2(n_557), .B1(n_566), .B2(n_565), .Y(n_910) );
NAND2x1p5_ASAP7_75t_L g911 ( .A(n_772), .B(n_557), .Y(n_911) );
UNKNOWN g912 ( );
INVx2_ASAP7_75t_L g913 ( .A(n_799), .Y(n_913) );
O2A1O1Ixp33_ASAP7_75t_L g914 ( .A1(n_763), .A2(n_565), .B(n_569), .C(n_566), .Y(n_914) );
OAI21x1_ASAP7_75t_L g915 ( .A1(n_806), .A2(n_566), .B(n_565), .Y(n_915) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_715), .A2(n_569), .B1(n_579), .B2(n_572), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_784), .A2(n_572), .B1(n_579), .B2(n_569), .Y(n_917) );
OAI21x1_ASAP7_75t_L g918 ( .A1(n_810), .A2(n_579), .B(n_572), .Y(n_918) );
AO31x2_ASAP7_75t_L g919 ( .A1(n_831), .A2(n_552), .A3(n_582), .B(n_404), .Y(n_919) );
BUFx3_ASAP7_75t_L g920 ( .A(n_772), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_732), .Y(n_921) );
OA21x2_ASAP7_75t_L g922 ( .A1(n_827), .A2(n_582), .B(n_610), .Y(n_922) );
AO21x1_ASAP7_75t_L g923 ( .A1(n_831), .A2(n_582), .B(n_121), .Y(n_923) );
BUFx3_ASAP7_75t_L g924 ( .A(n_774), .Y(n_924) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_787), .B(n_13), .Y(n_925) );
OA21x2_ASAP7_75t_L g926 ( .A1(n_814), .A2(n_582), .B(n_610), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_751), .Y(n_927) );
OAI21x1_ASAP7_75t_L g928 ( .A1(n_730), .A2(n_582), .B(n_122), .Y(n_928) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_766), .Y(n_929) );
OAI221xp5_ASAP7_75t_L g930 ( .A1(n_776), .A2(n_13), .B1(n_14), .B2(n_15), .C(n_17), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_740), .B(n_14), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_782), .A2(n_18), .B1(n_15), .B2(n_17), .Y(n_932) );
BUFx2_ASAP7_75t_L g933 ( .A(n_749), .Y(n_933) );
O2A1O1Ixp33_ASAP7_75t_SL g934 ( .A1(n_785), .A2(n_127), .B(n_129), .C(n_125), .Y(n_934) );
OA21x2_ASAP7_75t_L g935 ( .A1(n_742), .A2(n_620), .B(n_610), .Y(n_935) );
INVxp67_ASAP7_75t_L g936 ( .A(n_742), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_759), .A2(n_620), .B1(n_610), .B2(n_22), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_751), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_748), .A2(n_24), .B1(n_19), .B2(n_20), .Y(n_939) );
OAI21x1_ASAP7_75t_L g940 ( .A1(n_777), .A2(n_131), .B(n_130), .Y(n_940) );
O2A1O1Ixp33_ASAP7_75t_SL g941 ( .A1(n_779), .A2(n_144), .B(n_146), .C(n_136), .Y(n_941) );
OA21x2_ASAP7_75t_L g942 ( .A1(n_780), .A2(n_620), .B(n_610), .Y(n_942) );
NAND2x1p5_ASAP7_75t_L g943 ( .A(n_748), .B(n_24), .Y(n_943) );
CKINVDCx11_ASAP7_75t_R g944 ( .A(n_801), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_791), .A2(n_620), .B1(n_610), .B2(n_28), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_789), .B(n_26), .Y(n_946) );
BUFx3_ASAP7_75t_L g947 ( .A(n_835), .Y(n_947) );
BUFx6f_ASAP7_75t_L g948 ( .A(n_751), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_737), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g950 ( .A1(n_771), .A2(n_29), .B1(n_26), .B2(n_27), .Y(n_950) );
BUFx2_ASAP7_75t_L g951 ( .A(n_803), .Y(n_951) );
AO31x2_ASAP7_75t_L g952 ( .A1(n_811), .A2(n_31), .A3(n_29), .B(n_30), .Y(n_952) );
OAI21x1_ASAP7_75t_L g953 ( .A1(n_812), .A2(n_148), .B(n_147), .Y(n_953) );
AO21x2_ASAP7_75t_L g954 ( .A1(n_753), .A2(n_620), .B(n_610), .Y(n_954) );
INVx2_ASAP7_75t_L g955 ( .A(n_755), .Y(n_955) );
BUFx3_ASAP7_75t_L g956 ( .A(n_834), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g957 ( .A1(n_773), .A2(n_620), .B1(n_33), .B2(n_30), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_755), .Y(n_958) );
NOR2xp33_ASAP7_75t_SL g959 ( .A(n_805), .B(n_31), .Y(n_959) );
OAI21x1_ASAP7_75t_L g960 ( .A1(n_815), .A2(n_156), .B(n_149), .Y(n_960) );
INVx5_ASAP7_75t_L g961 ( .A(n_842), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_755), .Y(n_962) );
OAI21x1_ASAP7_75t_L g963 ( .A1(n_819), .A2(n_161), .B(n_159), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g964 ( .A1(n_750), .A2(n_33), .B1(n_34), .B2(n_35), .C(n_36), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_767), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_809), .A2(n_39), .B1(n_37), .B2(n_38), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_762), .A2(n_40), .B1(n_38), .B2(n_39), .Y(n_967) );
OAI21xp5_ASAP7_75t_L g968 ( .A1(n_757), .A2(n_163), .B(n_162), .Y(n_968) );
OAI21x1_ASAP7_75t_L g969 ( .A1(n_825), .A2(n_165), .B(n_164), .Y(n_969) );
OAI21x1_ASAP7_75t_L g970 ( .A1(n_830), .A2(n_167), .B(n_166), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g971 ( .A1(n_803), .A2(n_42), .B1(n_40), .B2(n_41), .Y(n_971) );
INVx2_ASAP7_75t_L g972 ( .A(n_767), .Y(n_972) );
NAND2x1p5_ASAP7_75t_L g973 ( .A(n_842), .B(n_41), .Y(n_973) );
OAI22xp33_ASAP7_75t_L g974 ( .A1(n_811), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_974) );
BUFx12f_ASAP7_75t_L g975 ( .A(n_805), .Y(n_975) );
INVx3_ASAP7_75t_L g976 ( .A(n_843), .Y(n_976) );
INVx4_ASAP7_75t_L g977 ( .A(n_843), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_767), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_765), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_769), .B(n_46), .Y(n_980) );
BUFx6f_ASAP7_75t_L g981 ( .A(n_778), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_783), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_790), .B(n_46), .Y(n_983) );
OAI21x1_ASAP7_75t_L g984 ( .A1(n_768), .A2(n_173), .B(n_168), .Y(n_984) );
AO31x2_ASAP7_75t_L g985 ( .A1(n_719), .A2(n_47), .A3(n_48), .B(n_49), .Y(n_985) );
AND2x4_ASAP7_75t_L g986 ( .A(n_717), .B(n_49), .Y(n_986) );
OAI21x1_ASAP7_75t_L g987 ( .A1(n_722), .A2(n_176), .B(n_174), .Y(n_987) );
INVx3_ASAP7_75t_L g988 ( .A(n_717), .Y(n_988) );
BUFx2_ASAP7_75t_L g989 ( .A(n_793), .Y(n_989) );
O2A1O1Ixp33_ASAP7_75t_L g990 ( .A1(n_813), .A2(n_50), .B(n_51), .C(n_52), .Y(n_990) );
OAI21x1_ASAP7_75t_L g991 ( .A1(n_724), .A2(n_179), .B(n_177), .Y(n_991) );
OAI21xp5_ASAP7_75t_L g992 ( .A1(n_726), .A2(n_182), .B(n_180), .Y(n_992) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_798), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_798), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_994) );
OAI21x1_ASAP7_75t_L g995 ( .A1(n_738), .A2(n_185), .B(n_184), .Y(n_995) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_912), .A2(n_824), .B1(n_829), .B2(n_747), .C(n_839), .Y(n_996) );
OAI21xp5_ASAP7_75t_L g997 ( .A1(n_896), .A2(n_832), .B(n_746), .Y(n_997) );
AOI21xp5_ASAP7_75t_L g998 ( .A1(n_901), .A2(n_786), .B(n_778), .Y(n_998) );
AOI21xp33_ASAP7_75t_L g999 ( .A1(n_861), .A2(n_837), .B(n_746), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_913), .Y(n_1000) );
OAI22xp33_ASAP7_75t_SL g1001 ( .A1(n_943), .A2(n_723), .B1(n_735), .B2(n_55), .Y(n_1001) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_936), .B(n_735), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g1003 ( .A1(n_951), .A2(n_808), .B1(n_807), .B2(n_795), .C(n_786), .Y(n_1003) );
A2O1A1Ixp33_ASAP7_75t_L g1004 ( .A1(n_936), .A2(n_808), .B(n_807), .C(n_795), .Y(n_1004) );
AOI221xp5_ASAP7_75t_L g1005 ( .A1(n_925), .A2(n_808), .B1(n_807), .B2(n_795), .C(n_786), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g1006 ( .A1(n_873), .A2(n_778), .B1(n_723), .B2(n_55), .Y(n_1006) );
NAND2xp33_ASAP7_75t_R g1007 ( .A(n_933), .B(n_53), .Y(n_1007) );
A2O1A1Ixp33_ASAP7_75t_L g1008 ( .A1(n_925), .A2(n_723), .B(n_54), .C(n_56), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_873), .A2(n_53), .B1(n_56), .B2(n_57), .Y(n_1009) );
AOI21xp5_ASAP7_75t_L g1010 ( .A1(n_901), .A2(n_189), .B(n_187), .Y(n_1010) );
INVx1_ASAP7_75t_SL g1011 ( .A(n_853), .Y(n_1011) );
NAND3xp33_ASAP7_75t_L g1012 ( .A(n_945), .B(n_58), .C(n_60), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_862), .B(n_60), .Y(n_1013) );
OA21x2_ASAP7_75t_L g1014 ( .A1(n_845), .A2(n_191), .B(n_190), .Y(n_1014) );
INVx1_ASAP7_75t_SL g1015 ( .A(n_893), .Y(n_1015) );
BUFx4f_ASAP7_75t_SL g1016 ( .A(n_856), .Y(n_1016) );
INVx2_ASAP7_75t_L g1017 ( .A(n_913), .Y(n_1017) );
AOI221xp5_ASAP7_75t_L g1018 ( .A1(n_930), .A2(n_974), .B1(n_884), .B2(n_866), .C(n_881), .Y(n_1018) );
AOI22xp33_ASAP7_75t_SL g1019 ( .A1(n_959), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_850), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_897), .Y(n_1021) );
O2A1O1Ixp33_ASAP7_75t_L g1022 ( .A1(n_883), .A2(n_61), .B(n_62), .C(n_63), .Y(n_1022) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_864), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_902), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_921), .B(n_67), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_949), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_850), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1028 ( .A(n_867), .B(n_920), .Y(n_1028) );
OAI21xp5_ASAP7_75t_L g1029 ( .A1(n_866), .A2(n_69), .B(n_70), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_847), .A2(n_71), .B1(n_72), .B2(n_73), .Y(n_1030) );
OAI22xp33_ASAP7_75t_L g1031 ( .A1(n_875), .A2(n_74), .B1(n_75), .B2(n_76), .Y(n_1031) );
A2O1A1Ixp33_ASAP7_75t_L g1032 ( .A1(n_990), .A2(n_75), .B(n_77), .C(n_78), .Y(n_1032) );
AOI21xp33_ASAP7_75t_L g1033 ( .A1(n_861), .A2(n_79), .B(n_80), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_863), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_1034) );
AO21x2_ASAP7_75t_L g1035 ( .A1(n_854), .A2(n_193), .B(n_192), .Y(n_1035) );
OAI22xp33_ASAP7_75t_L g1036 ( .A1(n_900), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_849), .A2(n_83), .B1(n_86), .B2(n_87), .Y(n_1037) );
AOI21x1_ASAP7_75t_L g1038 ( .A1(n_846), .A2(n_196), .B(n_195), .Y(n_1038) );
AOI21xp5_ASAP7_75t_L g1039 ( .A1(n_848), .A2(n_198), .B(n_197), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_986), .A2(n_89), .B1(n_91), .B2(n_92), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_868), .B(n_92), .Y(n_1041) );
INVx2_ASAP7_75t_L g1042 ( .A(n_851), .Y(n_1042) );
INVx1_ASAP7_75t_SL g1043 ( .A(n_989), .Y(n_1043) );
AOI22xp5_ASAP7_75t_L g1044 ( .A1(n_974), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_1044) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_871), .A2(n_93), .B1(n_95), .B2(n_96), .Y(n_1045) );
BUFx12f_ASAP7_75t_L g1046 ( .A(n_856), .Y(n_1046) );
NAND3xp33_ASAP7_75t_L g1047 ( .A(n_945), .B(n_98), .C(n_99), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_986), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_1048) );
OAI21xp5_ASAP7_75t_L g1049 ( .A1(n_898), .A2(n_100), .B(n_101), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_851), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_973), .Y(n_1051) );
AND2x4_ASAP7_75t_L g1052 ( .A(n_924), .B(n_101), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_947), .B(n_105), .Y(n_1053) );
AOI211xp5_ASAP7_75t_L g1054 ( .A1(n_966), .A2(n_107), .B(n_108), .C(n_109), .Y(n_1054) );
INVx2_ASAP7_75t_L g1055 ( .A(n_855), .Y(n_1055) );
NAND2xp5_ASAP7_75t_SL g1056 ( .A(n_961), .B(n_112), .Y(n_1056) );
AOI22xp5_ASAP7_75t_L g1057 ( .A1(n_964), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_1057) );
AND2x4_ASAP7_75t_L g1058 ( .A(n_865), .B(n_116), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_857), .B(n_117), .Y(n_1059) );
AO31x2_ASAP7_75t_L g1060 ( .A1(n_923), .A2(n_118), .A3(n_119), .B(n_201), .Y(n_1060) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_943), .A2(n_118), .B1(n_205), .B2(n_208), .Y(n_1061) );
BUFx5_ASAP7_75t_L g1062 ( .A(n_865), .Y(n_1062) );
OAI21x1_ASAP7_75t_L g1063 ( .A1(n_905), .A2(n_209), .B(n_211), .Y(n_1063) );
AND2x4_ASAP7_75t_L g1064 ( .A(n_876), .B(n_212), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g1065 ( .A1(n_904), .A2(n_215), .B1(n_217), .B2(n_218), .C(n_220), .Y(n_1065) );
INVx2_ASAP7_75t_L g1066 ( .A(n_855), .Y(n_1066) );
INVx11_ASAP7_75t_L g1067 ( .A(n_975), .Y(n_1067) );
AO21x2_ASAP7_75t_L g1068 ( .A1(n_894), .A2(n_223), .B(n_224), .Y(n_1068) );
INVx2_ASAP7_75t_L g1069 ( .A(n_872), .Y(n_1069) );
OR2x2_ASAP7_75t_L g1070 ( .A(n_947), .B(n_228), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_931), .A2(n_229), .B1(n_230), .B2(n_235), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_879), .A2(n_236), .B1(n_237), .B2(n_238), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_973), .Y(n_1073) );
HB1xp67_ASAP7_75t_L g1074 ( .A(n_993), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_872), .Y(n_1075) );
OAI211xp5_ASAP7_75t_L g1076 ( .A1(n_971), .A2(n_241), .B(n_244), .C(n_245), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_979), .Y(n_1077) );
AND2x6_ASAP7_75t_L g1078 ( .A(n_876), .B(n_251), .Y(n_1078) );
OAI21xp33_ASAP7_75t_L g1079 ( .A1(n_894), .A2(n_252), .B(n_254), .Y(n_1079) );
BUFx12f_ASAP7_75t_L g1080 ( .A(n_944), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_982), .B(n_356), .Y(n_1081) );
AOI221xp5_ASAP7_75t_L g1082 ( .A1(n_858), .A2(n_255), .B1(n_257), .B2(n_259), .C(n_260), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_980), .Y(n_1083) );
INVx2_ASAP7_75t_L g1084 ( .A(n_889), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_889), .Y(n_1085) );
AOI21x1_ASAP7_75t_L g1086 ( .A1(n_935), .A2(n_264), .B(n_268), .Y(n_1086) );
OAI211xp5_ASAP7_75t_L g1087 ( .A1(n_990), .A2(n_271), .B(n_272), .C(n_273), .Y(n_1087) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_874), .Y(n_1088) );
OAI211xp5_ASAP7_75t_L g1089 ( .A1(n_967), .A2(n_282), .B(n_283), .C(n_285), .Y(n_1089) );
BUFx5_ASAP7_75t_L g1090 ( .A(n_956), .Y(n_1090) );
OAI21x1_ASAP7_75t_L g1091 ( .A1(n_928), .A2(n_287), .B(n_288), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_887), .B(n_289), .Y(n_1092) );
OAI221xp5_ASAP7_75t_L g1093 ( .A1(n_937), .A2(n_290), .B1(n_293), .B2(n_294), .C(n_295), .Y(n_1093) );
AO221x1_ASAP7_75t_L g1094 ( .A1(n_932), .A2(n_297), .B1(n_298), .B2(n_299), .C(n_300), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_988), .B(n_302), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_952), .Y(n_1096) );
BUFx4f_ASAP7_75t_SL g1097 ( .A(n_870), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_957), .A2(n_303), .B1(n_304), .B2(n_306), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_879), .B(n_307), .Y(n_1099) );
OR2x2_ASAP7_75t_L g1100 ( .A(n_895), .B(n_311), .Y(n_1100) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_870), .Y(n_1101) );
INVx4_ASAP7_75t_L g1102 ( .A(n_961), .Y(n_1102) );
NAND3xp33_ASAP7_75t_L g1103 ( .A(n_937), .B(n_314), .C(n_315), .Y(n_1103) );
AND2x4_ASAP7_75t_SL g1104 ( .A(n_977), .B(n_316), .Y(n_1104) );
OAI22xp33_ASAP7_75t_L g1105 ( .A1(n_950), .A2(n_319), .B1(n_321), .B2(n_322), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_891), .B(n_325), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_967), .A2(n_327), .B1(n_328), .B2(n_330), .Y(n_1107) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_891), .B(n_334), .Y(n_1108) );
INVx2_ASAP7_75t_L g1109 ( .A(n_935), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_935), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_952), .Y(n_1111) );
OR2x2_ASAP7_75t_L g1112 ( .A(n_956), .B(n_335), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_952), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_952), .Y(n_1114) );
BUFx8_ASAP7_75t_SL g1115 ( .A(n_929), .Y(n_1115) );
NAND2xp5_ASAP7_75t_SL g1116 ( .A(n_961), .B(n_336), .Y(n_1116) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_993), .A2(n_338), .B1(n_340), .B2(n_342), .Y(n_1117) );
BUFx12f_ASAP7_75t_L g1118 ( .A(n_944), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_869), .A2(n_347), .B1(n_348), .B2(n_353), .Y(n_1119) );
INVx2_ASAP7_75t_SL g1120 ( .A(n_961), .Y(n_1120) );
OA21x2_ASAP7_75t_L g1121 ( .A1(n_877), .A2(n_355), .B(n_963), .Y(n_1121) );
AOI22x1_ASAP7_75t_L g1122 ( .A1(n_968), .A2(n_977), .B1(n_911), .B2(n_888), .Y(n_1122) );
OAI21xp33_ASAP7_75t_L g1123 ( .A1(n_917), .A2(n_909), .B(n_946), .Y(n_1123) );
A2O1A1Ixp33_ASAP7_75t_L g1124 ( .A1(n_914), .A2(n_880), .B(n_882), .C(n_890), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_983), .A2(n_885), .B1(n_939), .B2(n_916), .Y(n_1125) );
AOI21xp5_ASAP7_75t_L g1126 ( .A1(n_954), .A2(n_942), .B(n_885), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_886), .B(n_985), .Y(n_1127) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_976), .B(n_859), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1129 ( .A(n_886), .B(n_911), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_886), .B(n_976), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_985), .B(n_994), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_916), .A2(n_917), .B1(n_892), .B2(n_878), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_899), .A2(n_910), .B1(n_903), .B2(n_907), .Y(n_1133) );
OR2x2_ASAP7_75t_L g1134 ( .A(n_919), .B(n_985), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_919), .B(n_906), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_899), .A2(n_903), .B1(n_907), .B2(n_859), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1109), .Y(n_1137) );
INVx3_ASAP7_75t_L g1138 ( .A(n_1102), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1021), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1110), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1024), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1142 ( .A(n_1015), .B(n_919), .Y(n_1142) );
AND2x4_ASAP7_75t_L g1143 ( .A(n_1051), .B(n_859), .Y(n_1143) );
OAI22xp33_ASAP7_75t_L g1144 ( .A1(n_1034), .A2(n_899), .B1(n_992), .B2(n_859), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1000), .B(n_972), .Y(n_1145) );
AND2x4_ASAP7_75t_L g1146 ( .A(n_1073), .B(n_962), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1026), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1017), .B(n_972), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1020), .B(n_927), .Y(n_1149) );
NOR2xp33_ASAP7_75t_SL g1150 ( .A(n_1097), .B(n_981), .Y(n_1150) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1027), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1077), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1042), .B(n_927), .Y(n_1153) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1050), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1074), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1055), .B(n_962), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1066), .B(n_938), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1025), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1069), .B(n_938), .Y(n_1159) );
AND2x4_ASAP7_75t_L g1160 ( .A(n_1102), .B(n_978), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1075), .B(n_965), .Y(n_1161) );
NAND2x1_ASAP7_75t_L g1162 ( .A(n_1078), .B(n_948), .Y(n_1162) );
OR2x2_ASAP7_75t_L g1163 ( .A(n_1015), .B(n_1096), .Y(n_1163) );
INVx4_ASAP7_75t_L g1164 ( .A(n_1078), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1018), .B(n_1013), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1084), .B(n_965), .Y(n_1166) );
INVx4_ASAP7_75t_L g1167 ( .A(n_1078), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1111), .B(n_958), .Y(n_1168) );
INVx1_ASAP7_75t_SL g1169 ( .A(n_1011), .Y(n_1169) );
AND2x4_ASAP7_75t_L g1170 ( .A(n_1128), .B(n_955), .Y(n_1170) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1085), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1172 ( .A(n_1043), .B(n_955), .Y(n_1172) );
AND2x4_ASAP7_75t_SL g1173 ( .A(n_1002), .B(n_948), .Y(n_1173) );
INVx2_ASAP7_75t_L g1174 ( .A(n_1086), .Y(n_1174) );
NAND2xp33_ASAP7_75t_R g1175 ( .A(n_1101), .B(n_926), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1113), .B(n_978), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1044), .B(n_926), .Y(n_1177) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1129), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1044), .B(n_926), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1029), .B(n_922), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_1012), .A2(n_852), .B1(n_860), .B2(n_922), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1127), .B(n_922), .Y(n_1182) );
OR2x6_ASAP7_75t_L g1183 ( .A(n_1064), .B(n_981), .Y(n_1183) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1014), .Y(n_1184) );
BUFx2_ASAP7_75t_L g1185 ( .A(n_1062), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1083), .B(n_981), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_1114), .B(n_981), .Y(n_1187) );
AOI22xp5_ASAP7_75t_SL g1188 ( .A1(n_1088), .A2(n_948), .B1(n_941), .B2(n_942), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1058), .B(n_954), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1049), .B(n_984), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1053), .Y(n_1191) );
CKINVDCx11_ASAP7_75t_R g1192 ( .A(n_1046), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1002), .B(n_995), .Y(n_1193) );
CKINVDCx5p33_ASAP7_75t_R g1194 ( .A(n_1067), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1052), .Y(n_1195) );
BUFx6f_ASAP7_75t_L g1196 ( .A(n_1120), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1011), .B(n_940), .Y(n_1197) );
NOR2xp33_ASAP7_75t_L g1198 ( .A(n_1028), .B(n_934), .Y(n_1198) );
INVx2_ASAP7_75t_SL g1199 ( .A(n_1062), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1090), .B(n_991), .Y(n_1200) );
INVx2_ASAP7_75t_SL g1201 ( .A(n_1062), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1090), .B(n_987), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1090), .B(n_970), .Y(n_1203) );
BUFx3_ASAP7_75t_L g1204 ( .A(n_1062), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1041), .B(n_942), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1090), .B(n_969), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1059), .Y(n_1207) );
BUFx2_ASAP7_75t_L g1208 ( .A(n_1090), .Y(n_1208) );
NOR2x1_ASAP7_75t_SL g1209 ( .A(n_1108), .B(n_934), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1023), .B(n_941), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1064), .B(n_953), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1099), .B(n_960), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1131), .B(n_918), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1070), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1034), .B(n_915), .Y(n_1215) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_1031), .A2(n_908), .B1(n_1057), .B2(n_1047), .Y(n_1216) );
INVx3_ASAP7_75t_L g1217 ( .A(n_1078), .Y(n_1217) );
INVx1_ASAP7_75t_SL g1218 ( .A(n_1016), .Y(n_1218) );
AND2x4_ASAP7_75t_L g1219 ( .A(n_997), .B(n_1130), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1054), .B(n_1092), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1037), .Y(n_1221) );
INVx2_ASAP7_75t_L g1222 ( .A(n_1134), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1036), .Y(n_1223) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1091), .Y(n_1224) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1063), .Y(n_1225) );
INVx2_ASAP7_75t_SL g1226 ( .A(n_1104), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1054), .B(n_1006), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1006), .B(n_1032), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1229 ( .A(n_1112), .B(n_1135), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1106), .B(n_1040), .Y(n_1230) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1121), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1048), .B(n_1009), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1028), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1121), .Y(n_1234) );
INVx2_ASAP7_75t_SL g1235 ( .A(n_1056), .Y(n_1235) );
OAI21xp5_ASAP7_75t_L g1236 ( .A1(n_1008), .A2(n_1047), .B(n_1012), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1030), .Y(n_1237) );
INVx5_ASAP7_75t_L g1238 ( .A(n_1080), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1057), .B(n_1060), .Y(n_1239) );
NAND2x1p5_ASAP7_75t_L g1240 ( .A(n_1100), .B(n_1116), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1022), .Y(n_1241) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1060), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1125), .B(n_1126), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1081), .Y(n_1244) );
NOR2xp33_ASAP7_75t_SL g1245 ( .A(n_1118), .B(n_1115), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1019), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1060), .B(n_1045), .Y(n_1247) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1038), .Y(n_1248) );
AND2x4_ASAP7_75t_L g1249 ( .A(n_1004), .B(n_1095), .Y(n_1249) );
BUFx2_ASAP7_75t_L g1250 ( .A(n_1005), .Y(n_1250) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1068), .Y(n_1251) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1068), .Y(n_1252) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1137), .Y(n_1253) );
BUFx2_ASAP7_75t_L g1254 ( .A(n_1164), .Y(n_1254) );
INVx3_ASAP7_75t_L g1255 ( .A(n_1164), .Y(n_1255) );
INVx1_ASAP7_75t_SL g1256 ( .A(n_1194), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1178), .B(n_1136), .Y(n_1257) );
OAI31xp33_ASAP7_75t_L g1258 ( .A1(n_1227), .A2(n_1001), .A3(n_1087), .B(n_1093), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1137), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1140), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1178), .B(n_1133), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1182), .B(n_1035), .Y(n_1262) );
BUFx3_ASAP7_75t_L g1263 ( .A(n_1196), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1140), .Y(n_1264) );
INVx2_ASAP7_75t_L g1265 ( .A(n_1182), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1222), .B(n_1033), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1222), .Y(n_1267) );
OR2x2_ASAP7_75t_L g1268 ( .A(n_1163), .B(n_1003), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_1220), .A2(n_1094), .B1(n_1103), .B2(n_1001), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1189), .B(n_1124), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1271 ( .A(n_1163), .B(n_1103), .Y(n_1271) );
OAI33xp33_ASAP7_75t_L g1272 ( .A1(n_1155), .A2(n_1105), .A3(n_1117), .B1(n_1098), .B2(n_1007), .B3(n_1079), .Y(n_1272) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1229), .B(n_1107), .Y(n_1273) );
AND2x4_ASAP7_75t_L g1274 ( .A(n_1164), .B(n_1167), .Y(n_1274) );
NOR3xp33_ASAP7_75t_L g1275 ( .A(n_1246), .B(n_1076), .C(n_1061), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1168), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1189), .B(n_1107), .Y(n_1277) );
INVx2_ASAP7_75t_L g1278 ( .A(n_1176), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1213), .B(n_1079), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_1220), .A2(n_996), .B1(n_1122), .B2(n_1123), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1176), .Y(n_1281) );
INVx2_ASAP7_75t_L g1282 ( .A(n_1151), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1213), .B(n_1119), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1187), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1239), .B(n_999), .Y(n_1285) );
INVx3_ASAP7_75t_L g1286 ( .A(n_1167), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1239), .B(n_1132), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1219), .B(n_1072), .Y(n_1288) );
BUFx2_ASAP7_75t_L g1289 ( .A(n_1208), .Y(n_1289) );
OAI21xp33_ASAP7_75t_L g1290 ( .A1(n_1227), .A2(n_1247), .B(n_1236), .Y(n_1290) );
AOI211xp5_ASAP7_75t_SL g1291 ( .A1(n_1217), .A2(n_1089), .B(n_1082), .C(n_1065), .Y(n_1291) );
INVx2_ASAP7_75t_L g1292 ( .A(n_1151), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1187), .Y(n_1293) );
INVx2_ASAP7_75t_L g1294 ( .A(n_1154), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1219), .B(n_1071), .Y(n_1295) );
HB1xp67_ASAP7_75t_L g1296 ( .A(n_1172), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1229), .B(n_998), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1142), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1142), .Y(n_1299) );
AOI221xp5_ASAP7_75t_L g1300 ( .A1(n_1223), .A2(n_1010), .B1(n_1039), .B2(n_1158), .C(n_1165), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1205), .B(n_1243), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1219), .B(n_1154), .Y(n_1302) );
OAI33xp33_ASAP7_75t_L g1303 ( .A1(n_1139), .A2(n_1141), .A3(n_1152), .B1(n_1147), .B2(n_1191), .B3(n_1214), .Y(n_1303) );
INVxp67_ASAP7_75t_L g1304 ( .A(n_1169), .Y(n_1304) );
OAI21xp5_ASAP7_75t_L g1305 ( .A1(n_1216), .A2(n_1241), .B(n_1210), .Y(n_1305) );
INVx2_ASAP7_75t_L g1306 ( .A(n_1171), .Y(n_1306) );
AND2x4_ASAP7_75t_L g1307 ( .A(n_1217), .B(n_1200), .Y(n_1307) );
BUFx2_ASAP7_75t_L g1308 ( .A(n_1208), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1145), .B(n_1148), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1145), .B(n_1148), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1149), .B(n_1153), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1242), .Y(n_1312) );
HB1xp67_ASAP7_75t_L g1313 ( .A(n_1186), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1149), .B(n_1153), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1156), .B(n_1157), .Y(n_1315) );
HB1xp67_ASAP7_75t_L g1316 ( .A(n_1186), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1243), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1159), .B(n_1161), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_1232), .A2(n_1230), .B1(n_1228), .B2(n_1221), .Y(n_1319) );
INVxp67_ASAP7_75t_SL g1320 ( .A(n_1175), .Y(n_1320) );
OAI21xp5_ASAP7_75t_SL g1321 ( .A1(n_1226), .A2(n_1144), .B(n_1240), .Y(n_1321) );
NAND3xp33_ASAP7_75t_SL g1322 ( .A(n_1245), .B(n_1218), .C(n_1150), .Y(n_1322) );
OAI21xp5_ASAP7_75t_L g1323 ( .A1(n_1215), .A2(n_1247), .B(n_1237), .Y(n_1323) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1231), .Y(n_1324) );
OR2x2_ASAP7_75t_L g1325 ( .A(n_1195), .B(n_1138), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1159), .B(n_1161), .Y(n_1326) );
INVx2_ASAP7_75t_L g1327 ( .A(n_1231), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1166), .B(n_1179), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1166), .B(n_1179), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_1207), .B(n_1233), .Y(n_1330) );
INVx2_ASAP7_75t_SL g1331 ( .A(n_1138), .Y(n_1331) );
INVxp67_ASAP7_75t_L g1332 ( .A(n_1138), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1259), .Y(n_1333) );
INVx2_ASAP7_75t_L g1334 ( .A(n_1324), .Y(n_1334) );
INVx2_ASAP7_75t_L g1335 ( .A(n_1324), .Y(n_1335) );
AND2x4_ASAP7_75t_L g1336 ( .A(n_1307), .B(n_1202), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1265), .B(n_1177), .Y(n_1337) );
AOI22xp5_ASAP7_75t_L g1338 ( .A1(n_1319), .A2(n_1244), .B1(n_1250), .B2(n_1235), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1260), .Y(n_1339) );
INVx2_ASAP7_75t_L g1340 ( .A(n_1327), .Y(n_1340) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1260), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1309), .B(n_1146), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1328), .B(n_1180), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1328), .B(n_1193), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1329), .B(n_1193), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1310), .B(n_1146), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1329), .B(n_1211), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1270), .B(n_1211), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1310), .B(n_1185), .Y(n_1349) );
INVx2_ASAP7_75t_L g1350 ( .A(n_1253), .Y(n_1350) );
BUFx2_ASAP7_75t_L g1351 ( .A(n_1254), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1264), .Y(n_1352) );
AOI32xp33_ASAP7_75t_L g1353 ( .A1(n_1254), .A2(n_1190), .A3(n_1215), .B1(n_1198), .B2(n_1235), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1270), .B(n_1212), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1311), .B(n_1201), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1287), .B(n_1212), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1311), .B(n_1199), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1314), .B(n_1199), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1267), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1287), .B(n_1190), .Y(n_1360) );
INVx2_ASAP7_75t_L g1361 ( .A(n_1282), .Y(n_1361) );
INVx2_ASAP7_75t_L g1362 ( .A(n_1282), .Y(n_1362) );
OR2x2_ASAP7_75t_L g1363 ( .A(n_1301), .B(n_1197), .Y(n_1363) );
INVx2_ASAP7_75t_L g1364 ( .A(n_1292), .Y(n_1364) );
OAI21x1_ASAP7_75t_L g1365 ( .A1(n_1305), .A2(n_1234), .B(n_1174), .Y(n_1365) );
NAND3xp33_ASAP7_75t_L g1366 ( .A(n_1275), .B(n_1188), .C(n_1238), .Y(n_1366) );
OR2x2_ASAP7_75t_L g1367 ( .A(n_1317), .B(n_1183), .Y(n_1367) );
OR2x2_ASAP7_75t_L g1368 ( .A(n_1317), .B(n_1183), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1285), .B(n_1202), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1302), .B(n_1252), .Y(n_1370) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1298), .B(n_1183), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1323), .B(n_1251), .Y(n_1372) );
INVx2_ASAP7_75t_L g1373 ( .A(n_1292), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1261), .B(n_1203), .Y(n_1374) );
NAND4xp25_ASAP7_75t_SL g1375 ( .A(n_1256), .B(n_1192), .C(n_1238), .D(n_1181), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1261), .B(n_1203), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1298), .B(n_1206), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1378 ( .A(n_1299), .B(n_1183), .Y(n_1378) );
OR2x2_ASAP7_75t_L g1379 ( .A(n_1299), .B(n_1240), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1312), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1315), .B(n_1206), .Y(n_1381) );
AND2x4_ASAP7_75t_L g1382 ( .A(n_1307), .B(n_1204), .Y(n_1382) );
AOI211x1_ASAP7_75t_SL g1383 ( .A1(n_1322), .A2(n_1174), .B(n_1248), .C(n_1184), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1294), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1318), .B(n_1204), .Y(n_1385) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_1284), .B(n_1162), .Y(n_1386) );
INVx2_ASAP7_75t_L g1387 ( .A(n_1294), .Y(n_1387) );
INVx2_ASAP7_75t_L g1388 ( .A(n_1306), .Y(n_1388) );
NAND2x1p5_ASAP7_75t_L g1389 ( .A(n_1255), .B(n_1160), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1318), .B(n_1143), .Y(n_1390) );
OR2x2_ASAP7_75t_L g1391 ( .A(n_1349), .B(n_1296), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1385), .B(n_1313), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1360), .B(n_1290), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1385), .B(n_1316), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1347), .B(n_1326), .Y(n_1395) );
NOR2xp33_ASAP7_75t_SL g1396 ( .A(n_1366), .B(n_1321), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1360), .B(n_1290), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1347), .B(n_1326), .Y(n_1398) );
AND2x4_ASAP7_75t_L g1399 ( .A(n_1351), .B(n_1274), .Y(n_1399) );
AND2x4_ASAP7_75t_L g1400 ( .A(n_1351), .B(n_1274), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1356), .B(n_1284), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1359), .B(n_1276), .Y(n_1402) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1333), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1344), .B(n_1304), .Y(n_1404) );
INVxp67_ASAP7_75t_L g1405 ( .A(n_1355), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1344), .B(n_1289), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1345), .B(n_1289), .Y(n_1407) );
AOI21xp5_ASAP7_75t_L g1408 ( .A1(n_1375), .A2(n_1321), .B(n_1258), .Y(n_1408) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1333), .Y(n_1409) );
OR2x2_ASAP7_75t_L g1410 ( .A(n_1381), .B(n_1278), .Y(n_1410) );
OAI21xp33_ASAP7_75t_L g1411 ( .A1(n_1353), .A2(n_1280), .B(n_1269), .Y(n_1411) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1354), .B(n_1281), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1343), .B(n_1308), .Y(n_1413) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1339), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1341), .Y(n_1415) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_1357), .B(n_1293), .Y(n_1416) );
NAND2xp5_ASAP7_75t_L g1417 ( .A(n_1354), .B(n_1281), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1352), .Y(n_1418) );
AND2x4_ASAP7_75t_L g1419 ( .A(n_1382), .B(n_1274), .Y(n_1419) );
OR2x2_ASAP7_75t_L g1420 ( .A(n_1358), .B(n_1293), .Y(n_1420) );
NAND2x1_ASAP7_75t_L g1421 ( .A(n_1382), .B(n_1274), .Y(n_1421) );
OR2x2_ASAP7_75t_L g1422 ( .A(n_1343), .B(n_1297), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1348), .B(n_1307), .Y(n_1423) );
OAI221xp5_ASAP7_75t_L g1424 ( .A1(n_1411), .A2(n_1338), .B1(n_1353), .B2(n_1258), .C(n_1320), .Y(n_1424) );
O2A1O1Ixp33_ASAP7_75t_L g1425 ( .A1(n_1408), .A2(n_1330), .B(n_1303), .C(n_1272), .Y(n_1425) );
INVx2_ASAP7_75t_L g1426 ( .A(n_1392), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1427 ( .A(n_1393), .B(n_1348), .Y(n_1427) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1416), .Y(n_1428) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1420), .Y(n_1429) );
INVxp67_ASAP7_75t_L g1430 ( .A(n_1391), .Y(n_1430) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1403), .Y(n_1431) );
OAI221xp5_ASAP7_75t_L g1432 ( .A1(n_1396), .A2(n_1300), .B1(n_1389), .B2(n_1255), .C(n_1286), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1393), .B(n_1369), .Y(n_1433) );
OAI21xp5_ASAP7_75t_L g1434 ( .A1(n_1421), .A2(n_1332), .B(n_1331), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1409), .Y(n_1435) );
OAI22xp5_ASAP7_75t_L g1436 ( .A1(n_1405), .A2(n_1346), .B1(n_1342), .B2(n_1390), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1397), .B(n_1374), .Y(n_1437) );
OAI22xp33_ASAP7_75t_L g1438 ( .A1(n_1422), .A2(n_1331), .B1(n_1273), .B2(n_1379), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1395), .B(n_1374), .Y(n_1439) );
OAI22xp5_ASAP7_75t_L g1440 ( .A1(n_1399), .A2(n_1336), .B1(n_1382), .B2(n_1268), .Y(n_1440) );
OR2x2_ASAP7_75t_L g1441 ( .A(n_1410), .B(n_1363), .Y(n_1441) );
OAI31xp33_ASAP7_75t_L g1442 ( .A1(n_1400), .A2(n_1291), .A3(n_1288), .B(n_1295), .Y(n_1442) );
AOI22xp5_ASAP7_75t_L g1443 ( .A1(n_1424), .A2(n_1404), .B1(n_1417), .B2(n_1412), .Y(n_1443) );
AOI21xp33_ASAP7_75t_L g1444 ( .A1(n_1425), .A2(n_1325), .B(n_1402), .Y(n_1444) );
AOI22xp5_ASAP7_75t_L g1445 ( .A1(n_1424), .A2(n_1417), .B1(n_1412), .B2(n_1406), .Y(n_1445) );
AND4x1_ASAP7_75t_L g1446 ( .A(n_1442), .B(n_1383), .C(n_1398), .D(n_1413), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1426), .B(n_1423), .Y(n_1447) );
AO22x1_ASAP7_75t_L g1448 ( .A1(n_1434), .A2(n_1419), .B1(n_1394), .B2(n_1407), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1431), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1428), .B(n_1401), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1451 ( .A(n_1429), .B(n_1376), .Y(n_1451) );
INVx2_ASAP7_75t_L g1452 ( .A(n_1435), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1433), .B(n_1376), .Y(n_1453) );
AOI222xp33_ASAP7_75t_L g1454 ( .A1(n_1430), .A2(n_1372), .B1(n_1415), .B2(n_1414), .C1(n_1418), .C2(n_1337), .Y(n_1454) );
AOI22xp5_ASAP7_75t_L g1455 ( .A1(n_1443), .A2(n_1440), .B1(n_1436), .B2(n_1432), .Y(n_1455) );
AOI221xp5_ASAP7_75t_L g1456 ( .A1(n_1444), .A2(n_1438), .B1(n_1427), .B2(n_1437), .C(n_1439), .Y(n_1456) );
NOR2xp67_ASAP7_75t_L g1457 ( .A(n_1445), .B(n_1441), .Y(n_1457) );
AOI31xp33_ASAP7_75t_L g1458 ( .A1(n_1454), .A2(n_1386), .A3(n_1271), .B(n_1368), .Y(n_1458) );
OAI21xp5_ASAP7_75t_L g1459 ( .A1(n_1446), .A2(n_1271), .B(n_1367), .Y(n_1459) );
OAI22xp33_ASAP7_75t_L g1460 ( .A1(n_1448), .A2(n_1371), .B1(n_1378), .B2(n_1263), .Y(n_1460) );
AOI221xp5_ASAP7_75t_L g1461 ( .A1(n_1458), .A2(n_1449), .B1(n_1450), .B2(n_1452), .C(n_1451), .Y(n_1461) );
AOI221xp5_ASAP7_75t_L g1462 ( .A1(n_1456), .A2(n_1453), .B1(n_1447), .B2(n_1337), .C(n_1377), .Y(n_1462) );
OA21x2_ASAP7_75t_L g1463 ( .A1(n_1459), .A2(n_1365), .B(n_1335), .Y(n_1463) );
AOI211xp5_ASAP7_75t_SL g1464 ( .A1(n_1460), .A2(n_1283), .B(n_1266), .C(n_1277), .Y(n_1464) );
NOR3xp33_ASAP7_75t_L g1465 ( .A(n_1455), .B(n_1143), .C(n_1266), .Y(n_1465) );
O2A1O1Ixp33_ASAP7_75t_L g1466 ( .A1(n_1457), .A2(n_1249), .B(n_1263), .C(n_1380), .Y(n_1466) );
AND2x4_ASAP7_75t_L g1467 ( .A(n_1465), .B(n_1370), .Y(n_1467) );
NAND4xp75_ASAP7_75t_L g1468 ( .A(n_1461), .B(n_1279), .C(n_1262), .D(n_1257), .Y(n_1468) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1462), .Y(n_1469) );
NOR4xp25_ASAP7_75t_L g1470 ( .A(n_1469), .B(n_1466), .C(n_1463), .D(n_1464), .Y(n_1470) );
NOR3xp33_ASAP7_75t_SL g1471 ( .A(n_1468), .B(n_1384), .C(n_1209), .Y(n_1471) );
INVx2_ASAP7_75t_L g1472 ( .A(n_1467), .Y(n_1472) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1472), .Y(n_1473) );
AOI22xp5_ASAP7_75t_L g1474 ( .A1(n_1473), .A2(n_1470), .B1(n_1471), .B2(n_1173), .Y(n_1474) );
OAI22xp5_ASAP7_75t_SL g1475 ( .A1(n_1474), .A2(n_1224), .B1(n_1225), .B2(n_1170), .Y(n_1475) );
AOI222xp33_ASAP7_75t_SL g1476 ( .A1(n_1475), .A2(n_1340), .B1(n_1334), .B2(n_1388), .C1(n_1361), .C2(n_1387), .Y(n_1476) );
AO221x2_ASAP7_75t_L g1477 ( .A1(n_1476), .A2(n_1362), .B1(n_1387), .B2(n_1373), .C(n_1364), .Y(n_1477) );
AOI22xp5_ASAP7_75t_L g1478 ( .A1(n_1477), .A2(n_1350), .B1(n_1364), .B2(n_1388), .Y(n_1478) );
endmodule