module fake_jpeg_13073_n_312 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_51),
.Y(n_139)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_53),
.Y(n_132)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_61),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_1),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_66),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_17),
.B(n_2),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_73),
.B(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_22),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_74),
.B(n_84),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_75),
.A2(n_4),
.B1(n_8),
.B2(n_11),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_25),
.B(n_13),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_88),
.Y(n_106)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_77),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_78),
.B(n_85),
.Y(n_130)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_86),
.Y(n_143)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_35),
.B(n_3),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_38),
.B(n_4),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_93),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_67),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_40),
.B1(n_18),
.B2(n_29),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_98),
.A2(n_120),
.B1(n_146),
.B2(n_147),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_48),
.A2(n_39),
.B1(n_33),
.B2(n_32),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_107),
.A2(n_121),
.B1(n_128),
.B2(n_105),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_59),
.A2(n_78),
.B1(n_87),
.B2(n_85),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_124),
.B1(n_103),
.B2(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_32),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_25),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_66),
.A2(n_29),
.B1(n_33),
.B2(n_9),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_50),
.A2(n_29),
.B1(n_8),
.B2(n_11),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_60),
.B(n_12),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_123),
.B(n_138),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_53),
.A2(n_13),
.B1(n_58),
.B2(n_75),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_117),
.B(n_143),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_84),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_76),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_96),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_55),
.A2(n_34),
.B1(n_66),
.B2(n_51),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_55),
.A2(n_34),
.B1(n_66),
.B2(n_51),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_149),
.A2(n_161),
.B1(n_180),
.B2(n_183),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_151),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_108),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_160),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_127),
.C(n_102),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_115),
.B1(n_109),
.B2(n_107),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_164),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_106),
.Y(n_164)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_98),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_110),
.B(n_104),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_120),
.A2(n_147),
.B1(n_115),
.B2(n_121),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_179),
.B1(n_185),
.B2(n_158),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_134),
.B1(n_139),
.B2(n_110),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_109),
.B(n_101),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_161),
.Y(n_189)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_114),
.B(n_129),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_139),
.A2(n_119),
.B1(n_111),
.B2(n_131),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_181),
.Y(n_191)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_105),
.A2(n_124),
.B1(n_128),
.B2(n_75),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_112),
.B(n_130),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_162),
.B(n_148),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_95),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_202),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_193),
.A2(n_201),
.B1(n_152),
.B2(n_187),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_183),
.B1(n_185),
.B2(n_170),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_160),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_176),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_214),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_165),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_215),
.Y(n_216)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_213),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_219),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_210),
.A2(n_185),
.B1(n_154),
.B2(n_186),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_218),
.A2(n_193),
.B1(n_189),
.B2(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_225),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_190),
.B(n_169),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_153),
.C(n_175),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_237),
.Y(n_244)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

NOR2x1_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_205),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_233),
.B(n_238),
.Y(n_250)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_230),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_229),
.Y(n_242)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_236),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_182),
.C(n_177),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_156),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_194),
.B1(n_212),
.B2(n_190),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_239),
.B1(n_222),
.B2(n_224),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_249),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_234),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_211),
.B(n_191),
.Y(n_251)
);

AO221x1_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_238),
.B1(n_237),
.B2(n_218),
.C(n_219),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_225),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_231),
.A2(n_207),
.B(n_197),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_254),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_250),
.B1(n_245),
.B2(n_248),
.Y(n_275)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

OAI322xp33_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_251),
.A3(n_249),
.B1(n_253),
.B2(n_254),
.C1(n_244),
.C2(n_257),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_261),
.A2(n_263),
.B1(n_240),
.B2(n_247),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_220),
.C(n_227),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_242),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_238),
.C(n_207),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_270),
.C(n_248),
.Y(n_277)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_235),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_265),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_230),
.CI(n_226),
.CON(n_268),
.SN(n_268)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_247),
.CI(n_255),
.CON(n_279),
.SN(n_279)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_271),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_206),
.C(n_204),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_257),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_280),
.B1(n_282),
.B2(n_260),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_275),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_250),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_277),
.C(n_259),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_258),
.B1(n_261),
.B2(n_267),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_269),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_270),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_286),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_278),
.A2(n_258),
.B(n_267),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_279),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_263),
.B(n_266),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_274),
.B1(n_278),
.B2(n_279),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_271),
.C(n_255),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_291),
.C(n_283),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_243),
.C(n_268),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_296),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_287),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_291),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_294),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_298),
.B(n_301),
.Y(n_304)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_299),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_302),
.B(n_296),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_300),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_300),
.C(n_301),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_290),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_304),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_308),
.B(n_309),
.C(n_293),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_285),
.C(n_268),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_243),
.Y(n_312)
);


endmodule