module fake_jpeg_11212_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_19),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g62 ( 
.A(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_1),
.Y(n_60)
);

NAND4xp25_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_39),
.C(n_38),
.D(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_5),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_49),
.B1(n_48),
.B2(n_52),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_4),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_6),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_37),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_78),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_45),
.C(n_68),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_79),
.C(n_85),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_61),
.B1(n_49),
.B2(n_43),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_82),
.B1(n_12),
.B2(n_23),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_53),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_42),
.C(n_21),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_83),
.B(n_87),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_6),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_9),
.C(n_10),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_88),
.A2(n_66),
.B1(n_14),
.B2(n_15),
.Y(n_90)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_93),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_66),
.B1(n_18),
.B2(n_22),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_94),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_30),
.B(n_31),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_111),
.B(n_101),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_32),
.C(n_34),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.C(n_110),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_97),
.B(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_118),
.Y(n_121)
);

OA21x2_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_116),
.B(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_106),
.Y(n_124)
);


endmodule