module fake_jpeg_20487_n_71 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_70;
wire n_15;
wire n_66;

INVx2_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_19),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_17),
.B(n_0),
.Y(n_20)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_16),
.B(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_20),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_15),
.B1(n_9),
.B2(n_8),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_23),
.B1(n_9),
.B2(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_34),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_18),
.C(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_22),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_28),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_21),
.B1(n_19),
.B2(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_19),
.B1(n_13),
.B2(n_10),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_22),
.B1(n_1),
.B2(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_44),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_32),
.C(n_41),
.Y(n_51)
);

XOR2x1_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_52),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_54),
.C(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_40),
.Y(n_52)
);

AO22x1_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_39),
.B1(n_36),
.B2(n_10),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_49),
.B1(n_3),
.B2(n_0),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_12),
.B(n_3),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_12),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_49),
.C(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_49),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_62),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_6),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_65),
.B(n_69),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_62),
.Y(n_71)
);


endmodule