module fake_jpeg_15951_n_355 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_355);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_52),
.Y(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_20),
.B(n_21),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_67),
.A2(n_37),
.B(n_30),
.C(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_17),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_27),
.B1(n_21),
.B2(n_33),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_33),
.B1(n_27),
.B2(n_37),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_41),
.B1(n_37),
.B2(n_27),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_37),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_79),
.B(n_100),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_39),
.C(n_43),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_82),
.B(n_32),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_91),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_84),
.B(n_98),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_104),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_88),
.Y(n_118)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_37),
.B(n_28),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_94),
.B(n_95),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_30),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_51),
.B1(n_48),
.B2(n_44),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_105),
.B1(n_111),
.B2(n_115),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_25),
.B(n_28),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_64),
.B(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_59),
.B(n_25),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_77),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_40),
.B1(n_31),
.B2(n_26),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_59),
.A2(n_43),
.B1(n_23),
.B2(n_24),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_77),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_64),
.A2(n_17),
.B1(n_34),
.B2(n_19),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_19),
.B1(n_34),
.B2(n_31),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_80),
.B1(n_96),
.B2(n_105),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_23),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_134),
.Y(n_157)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_24),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_95),
.B(n_24),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_138),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_137),
.B(n_108),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_24),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_140),
.B(n_82),
.Y(n_154)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_79),
.A2(n_31),
.B1(n_26),
.B2(n_32),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_103),
.B1(n_110),
.B2(n_81),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_152),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_150),
.B(n_155),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_156),
.B1(n_162),
.B2(n_165),
.Y(n_180)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_128),
.C(n_32),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_139),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_100),
.B1(n_94),
.B2(n_92),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_163),
.B(n_170),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_119),
.A2(n_90),
.B1(n_100),
.B2(n_111),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_119),
.A2(n_106),
.B(n_109),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_146),
.B(n_123),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_93),
.B1(n_111),
.B2(n_114),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_85),
.B1(n_97),
.B2(n_99),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_168),
.B1(n_169),
.B2(n_142),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_85),
.B1(n_97),
.B2(n_111),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_89),
.B1(n_26),
.B2(n_31),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_174),
.B1(n_122),
.B2(n_118),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_126),
.A2(n_107),
.B1(n_116),
.B2(n_88),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_35),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_177),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_32),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_179),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_9),
.B(n_16),
.C(n_15),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_188),
.B1(n_207),
.B2(n_158),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_183),
.A2(n_185),
.B(n_189),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_146),
.B(n_134),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_135),
.B(n_127),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_179),
.A2(n_144),
.B1(n_145),
.B2(n_124),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_191),
.B(n_196),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_124),
.B(n_132),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_140),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_199),
.C(n_204),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_122),
.B1(n_132),
.B2(n_137),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_205),
.B1(n_160),
.B2(n_177),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_128),
.B(n_125),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_159),
.B(n_153),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_203),
.A2(n_210),
.B(n_163),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_121),
.C(n_118),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_161),
.A2(n_120),
.B1(n_32),
.B2(n_35),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_2),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_35),
.B1(n_9),
.B2(n_10),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_0),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_1),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_170),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_173),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_213),
.C(n_2),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_35),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_215),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_198),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_184),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_218),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_226),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_198),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_202),
.B1(n_201),
.B2(n_205),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_183),
.B(n_176),
.CI(n_152),
.CON(n_224),
.SN(n_224)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_185),
.B(n_11),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_149),
.B(n_35),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_210),
.B(n_206),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_199),
.B(n_11),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_149),
.Y(n_231)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

XOR2x2_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_16),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_191),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_212),
.B(n_15),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_242),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_14),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_195),
.C(n_213),
.Y(n_248)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_14),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_240),
.B(n_13),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_195),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_3),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_246),
.C(n_249),
.Y(n_276)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_180),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_12),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_204),
.C(n_211),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_210),
.B1(n_187),
.B2(n_191),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_250),
.A2(n_253),
.B1(n_260),
.B2(n_261),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_190),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_259),
.C(n_201),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_226),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_247),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_258),
.B(n_12),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_182),
.C(n_186),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_231),
.A2(n_188),
.B1(n_186),
.B2(n_182),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_187),
.B(n_202),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_238),
.B1(n_230),
.B2(n_242),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_254),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_270),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_256),
.A2(n_217),
.B(n_216),
.Y(n_269)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_227),
.B1(n_224),
.B2(n_234),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_271),
.A2(n_274),
.B1(n_286),
.B2(n_250),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_224),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_273),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_241),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_223),
.B1(n_221),
.B2(n_225),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_219),
.B(n_222),
.C(n_228),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_277),
.B(n_288),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_229),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.C(n_289),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_235),
.Y(n_279)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_244),
.A2(n_222),
.B(n_225),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_263),
.B1(n_262),
.B2(n_5),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_261),
.A2(n_237),
.B1(n_201),
.B2(n_12),
.Y(n_286)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_243),
.C(n_260),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_301),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_252),
.C(n_248),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_280),
.A2(n_253),
.B(n_251),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_286),
.B(n_277),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_270),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_303),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_247),
.C(n_267),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_278),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_319),
.C(n_321),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_275),
.B(n_272),
.Y(n_311)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_288),
.B1(n_284),
.B2(n_271),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_312),
.A2(n_317),
.B1(n_298),
.B2(n_304),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_293),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_316),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_296),
.B(n_306),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_281),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_300),
.A2(n_289),
.B1(n_4),
.B2(n_5),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_11),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_3),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_297),
.Y(n_322)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_322),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_302),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_321),
.C(n_308),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_326),
.A2(n_330),
.B1(n_317),
.B2(n_4),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_332),
.Y(n_335)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_309),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_331),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_315),
.A2(n_295),
.B(n_305),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_314),
.A2(n_303),
.B(n_301),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_339),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_333),
.B(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_338),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_310),
.C(n_313),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_316),
.C(n_290),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_290),
.C(n_318),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_340),
.B(n_341),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_328),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_344),
.B(n_335),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_337),
.A2(n_327),
.B(n_4),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_345),
.B(n_335),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_347),
.A2(n_348),
.B(n_349),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_342),
.B(n_3),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_350),
.A2(n_346),
.B(n_343),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_351),
.A2(n_5),
.B(n_6),
.Y(n_352)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_8),
.B(n_6),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_8),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_6),
.B(n_7),
.Y(n_355)
);


endmodule