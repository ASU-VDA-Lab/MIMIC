module fake_jpeg_18644_n_345 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_48),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_52),
.A2(n_38),
.B1(n_20),
.B2(n_31),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_38),
.B1(n_23),
.B2(n_25),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_64),
.B1(n_23),
.B2(n_21),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_31),
.B1(n_20),
.B2(n_22),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_70),
.Y(n_81)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_28),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_75),
.B(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_42),
.B1(n_49),
.B2(n_45),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_78),
.A2(n_60),
.B1(n_69),
.B2(n_55),
.Y(n_121)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_84),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_66),
.B1(n_56),
.B2(n_69),
.Y(n_115)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_34),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_86),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_103),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_96),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_28),
.B1(n_32),
.B2(n_63),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_56),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_32),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_50),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_126),
.C(n_130),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_110),
.B(n_111),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_76),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_121),
.B1(n_129),
.B2(n_106),
.Y(n_142)
);

NAND2x1_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_50),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_102),
.Y(n_143)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_25),
.B(n_30),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_95),
.A2(n_36),
.B(n_26),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_88),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_136),
.Y(n_141)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_81),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_118),
.C(n_128),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_139),
.B(n_144),
.Y(n_182)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_142),
.A2(n_54),
.B1(n_94),
.B2(n_93),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_119),
.B(n_130),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_26),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_152),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_78),
.B1(n_100),
.B2(n_96),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_146),
.A2(n_159),
.B1(n_127),
.B2(n_122),
.Y(n_179)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_84),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_77),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_109),
.B(n_26),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_153),
.A2(n_157),
.B1(n_136),
.B2(n_120),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_43),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_43),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_106),
.A2(n_67),
.B1(n_51),
.B2(n_45),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_162),
.A2(n_168),
.B(n_80),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_110),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_164),
.A2(n_26),
.B(n_35),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_121),
.B1(n_111),
.B2(n_107),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_177),
.B1(n_188),
.B2(n_116),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_125),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_187),
.Y(n_195)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_183),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_107),
.C(n_8),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_86),
.B(n_141),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_127),
.B1(n_120),
.B2(n_128),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_184),
.B1(n_73),
.B2(n_39),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_122),
.B1(n_94),
.B2(n_123),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_93),
.B1(n_116),
.B2(n_117),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_156),
.C(n_143),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_24),
.C(n_26),
.Y(n_207)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_143),
.A2(n_134),
.B1(n_90),
.B2(n_99),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_164),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_196),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_191),
.C(n_198),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_146),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_R g192 ( 
.A(n_162),
.B(n_161),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_192),
.B(n_163),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_193),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_133),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

AO22x2_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_159),
.B1(n_155),
.B2(n_160),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_138),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_197),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_153),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_157),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_207),
.C(n_209),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_206),
.B1(n_196),
.B2(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_138),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_213),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_117),
.B1(n_77),
.B2(n_51),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_210),
.B1(n_214),
.B2(n_211),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_138),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_211),
.B(n_192),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_39),
.C(n_24),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_36),
.B1(n_14),
.B2(n_17),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_215),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_36),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_36),
.B1(n_13),
.B2(n_17),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_29),
.B1(n_37),
.B2(n_33),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_218),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_37),
.B1(n_33),
.B2(n_27),
.Y(n_218)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_173),
.Y(n_226)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_244),
.B1(n_210),
.B2(n_217),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_208),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_235),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_187),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_239),
.B1(n_234),
.B2(n_238),
.Y(n_259)
);

OAI32xp33_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_163),
.A3(n_178),
.B1(n_171),
.B2(n_169),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_241),
.B(n_212),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_185),
.B1(n_12),
.B2(n_13),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_190),
.B(n_169),
.C(n_166),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_198),
.C(n_207),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_191),
.B1(n_199),
.B2(n_166),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_258),
.C(n_266),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_235),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_222),
.B(n_209),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_255),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_221),
.B1(n_233),
.B2(n_241),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_264),
.B1(n_231),
.B2(n_224),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_83),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_227),
.A2(n_35),
.B1(n_27),
.B2(n_11),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_263),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_240),
.C(n_244),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_262),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_238),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_219),
.B(n_237),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_37),
.C(n_33),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_83),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_27),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_267),
.A2(n_277),
.B1(n_37),
.B2(n_33),
.Y(n_300)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_219),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_245),
.Y(n_287)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_275),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_221),
.B1(n_233),
.B2(n_229),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_281),
.Y(n_286)
);

AOI21x1_ASAP7_75t_SL g280 ( 
.A1(n_248),
.A2(n_228),
.B(n_231),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_232),
.B(n_258),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_257),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_284),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_260),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_282),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_259),
.B(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_289),
.B(n_285),
.Y(n_309)
);

OA21x2_ASAP7_75t_SL g292 ( 
.A1(n_275),
.A2(n_247),
.B(n_230),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_292),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_296),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_9),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_300),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_35),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_271),
.B(n_293),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_267),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_278),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_304),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_281),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_291),
.C(n_290),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_273),
.C(n_282),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_300),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_268),
.B1(n_279),
.B2(n_269),
.Y(n_307)
);

OA22x2_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_308),
.B1(n_312),
.B2(n_298),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_276),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_289),
.A2(n_270),
.B1(n_273),
.B2(n_285),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_295),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_287),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_291),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_319),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_322),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_321),
.Y(n_332)
);

NAND4xp25_ASAP7_75t_SL g322 ( 
.A(n_311),
.B(n_301),
.C(n_288),
.D(n_4),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_7),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_324),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_7),
.Y(n_324)
);

NOR2x1_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_307),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_5),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_302),
.B1(n_306),
.B2(n_4),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_329),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_10),
.C(n_3),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_11),
.C(n_3),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_5),
.C(n_6),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_323),
.Y(n_333)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_333),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_334),
.A2(n_335),
.B(n_337),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_5),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_331),
.B(n_327),
.Y(n_341)
);

AOI322xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_331),
.A3(n_325),
.B1(n_338),
.B2(n_336),
.C1(n_14),
.C2(n_13),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_342),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_16),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_16),
.B(n_1),
.Y(n_345)
);


endmodule