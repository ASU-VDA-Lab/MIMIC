module fake_jpeg_20817_n_164 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp67_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_39),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_35),
.Y(n_62)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_42),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.C(n_1),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_1),
.C(n_2),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_43),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_54),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_22),
.B1(n_19),
.B2(n_28),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_59),
.B1(n_44),
.B2(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_22),
.B1(n_18),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_32),
.B1(n_42),
.B2(n_33),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_3),
.B(n_4),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_61),
.B(n_5),
.C(n_7),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_32),
.A2(n_18),
.B1(n_19),
.B2(n_25),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_3),
.B(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_27),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_41),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_75),
.B1(n_80),
.B2(n_85),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_36),
.A3(n_15),
.B1(n_30),
.B2(n_21),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_49),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_15),
.B(n_30),
.C(n_24),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_24),
.B(n_25),
.C(n_20),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_78),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_74),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_36),
.B1(n_31),
.B2(n_17),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_44),
.A2(n_31),
.B1(n_17),
.B2(n_5),
.Y(n_79)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_82),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_41),
.B1(n_31),
.B2(n_17),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_59),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_64),
.B(n_61),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_85),
.B1(n_86),
.B2(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_62),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_62),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_70),
.C(n_41),
.Y(n_111)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

XNOR2x1_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_87),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_112),
.B(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_80),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_115),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_97),
.C(n_103),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_71),
.C(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_73),
.C(n_62),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_117),
.B(n_97),
.Y(n_127)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_120),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_90),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_101),
.B1(n_102),
.B2(n_97),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_129),
.B1(n_132),
.B2(n_111),
.Y(n_136)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_113),
.C(n_112),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_118),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_101),
.B1(n_92),
.B2(n_90),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_109),
.B(n_116),
.C(n_110),
.D(n_114),
.Y(n_131)
);

INVxp67_ASAP7_75t_R g141 ( 
.A(n_131),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_107),
.B1(n_106),
.B2(n_119),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_129),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_138),
.C(n_142),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_115),
.C(n_98),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_105),
.B1(n_95),
.B2(n_78),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_130),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_127),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_118),
.C(n_95),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_146),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_138),
.Y(n_144)
);

AOI31xp33_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_128),
.A3(n_131),
.B(n_142),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_133),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_141),
.A3(n_123),
.B1(n_128),
.B2(n_131),
.C1(n_124),
.C2(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_145),
.A2(n_122),
.B1(n_135),
.B2(n_141),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_145),
.B(n_130),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_153),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_147),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_11),
.A3(n_14),
.B1(n_9),
.B2(n_10),
.C1(n_84),
.C2(n_74),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_153),
.A3(n_150),
.B1(n_83),
.B2(n_76),
.C1(n_62),
.C2(n_47),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_140),
.B(n_125),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_150),
.B(n_13),
.Y(n_160)
);

OAI311xp33_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_160),
.A3(n_156),
.B1(n_9),
.C1(n_7),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_5),
.C(n_7),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.Y(n_164)
);


endmodule