module fake_jpeg_22467_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_44),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_49),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_7),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_20),
.Y(n_69)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_57),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_34),
.B1(n_38),
.B2(n_27),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_63),
.B1(n_77),
.B2(n_82),
.Y(n_88)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_34),
.B1(n_38),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_34),
.B1(n_38),
.B2(n_25),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_26),
.Y(n_89)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_70),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_25),
.B1(n_28),
.B2(n_37),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_17),
.C(n_31),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_73),
.B(n_8),
.Y(n_119)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_28),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_37),
.B1(n_28),
.B2(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_37),
.B1(n_24),
.B2(n_22),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_18),
.B1(n_33),
.B2(n_19),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_30),
.B1(n_29),
.B2(n_35),
.Y(n_116)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_22),
.B1(n_24),
.B2(n_31),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_94),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_112),
.Y(n_128)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_103),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_97),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_36),
.B1(n_21),
.B2(n_26),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_93),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_21),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_21),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_29),
.B1(n_18),
.B2(n_33),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_107),
.B1(n_113),
.B2(n_116),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_30),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_109),
.Y(n_147)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_36),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_61),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_65),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_0),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_79),
.B(n_19),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_36),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_55),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_80),
.B(n_12),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_53),
.A2(n_8),
.B(n_14),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_7),
.B(n_13),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_54),
.B(n_0),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_8),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_55),
.A2(n_26),
.B1(n_20),
.B2(n_36),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_125),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_131),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_84),
.B(n_81),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_139),
.B(n_154),
.Y(n_162)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_132),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_57),
.B1(n_26),
.B2(n_20),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_117),
.B1(n_105),
.B2(n_93),
.Y(n_174)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_134),
.Y(n_169)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_65),
.C(n_20),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_155),
.C(n_107),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_141),
.B(n_112),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_95),
.A2(n_0),
.B(n_1),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_146),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_145),
.B1(n_153),
.B2(n_85),
.Y(n_172)
);

AO21x2_ASAP7_75t_L g145 ( 
.A1(n_93),
.A2(n_2),
.B(n_3),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_100),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_109),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_148),
.B(n_156),
.Y(n_158)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_102),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_86),
.A2(n_3),
.B(n_4),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_4),
.C(n_5),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_160),
.Y(n_207)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_176),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_94),
.C(n_111),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_173),
.C(n_183),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_165),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_99),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_123),
.B(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_99),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_178),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_185),
.B1(n_145),
.B2(n_150),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_96),
.C(n_110),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_174),
.A2(n_180),
.B1(n_188),
.B2(n_6),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_99),
.B(n_112),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_177),
.B(n_154),
.Y(n_195)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_120),
.B(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_120),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_93),
.B1(n_115),
.B2(n_108),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_115),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_182),
.A2(n_186),
.B1(n_191),
.B2(n_163),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_96),
.C(n_108),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_93),
.B1(n_121),
.B2(n_87),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_145),
.A2(n_87),
.B1(n_97),
.B2(n_91),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_147),
.B(n_113),
.Y(n_190)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_192),
.A2(n_174),
.B1(n_185),
.B2(n_189),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_126),
.B1(n_157),
.B2(n_137),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_214),
.B1(n_216),
.B2(n_218),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_196),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_141),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_155),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_209),
.C(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_205),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_153),
.B(n_141),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_219),
.B(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_138),
.B(n_130),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_211),
.B(n_217),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_181),
.C(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_212),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_162),
.A2(n_151),
.B(n_127),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_215),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_134),
.B1(n_133),
.B2(n_124),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_125),
.B1(n_6),
.B2(n_5),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_159),
.A2(n_188),
.B(n_166),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_172),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_218)
);

NAND2x1p5_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_180),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_219),
.B1(n_189),
.B2(n_200),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_158),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_193),
.B1(n_211),
.B2(n_218),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_228),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_199),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_227),
.C(n_209),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_171),
.C(n_160),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_198),
.B(n_190),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_231),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_235),
.B1(n_197),
.B2(n_203),
.Y(n_256)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_205),
.B(n_158),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_244),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_238),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_243),
.B(n_233),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_184),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_240),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_161),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_177),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_176),
.Y(n_246)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_247),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_192),
.B1(n_197),
.B2(n_208),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_248),
.A2(n_259),
.B1(n_264),
.B2(n_235),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_258),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_234),
.B1(n_247),
.B2(n_227),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_207),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_220),
.B1(n_194),
.B2(n_170),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_266),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_201),
.C(n_196),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_265),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_234),
.B1(n_243),
.B2(n_237),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_232),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_267),
.Y(n_273)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_271),
.Y(n_286)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_263),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_276),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_246),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_257),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_277),
.A2(n_278),
.B1(n_254),
.B2(n_226),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_230),
.B1(n_226),
.B2(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_281),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_250),
.A2(n_224),
.B1(n_244),
.B2(n_228),
.Y(n_282)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_245),
.Y(n_283)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_245),
.B(n_224),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_284),
.A2(n_266),
.B(n_229),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_256),
.A2(n_248),
.B1(n_264),
.B2(n_254),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_265),
.B(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_259),
.C(n_249),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_292),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_289),
.C(n_269),
.Y(n_300)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_255),
.C(n_262),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_280),
.C(n_258),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_300),
.A2(n_307),
.B(n_287),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_304),
.C(n_305),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_294),
.C(n_288),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_281),
.C(n_285),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_274),
.C(n_277),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_286),
.B(n_282),
.CI(n_278),
.CON(n_308),
.SN(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_270),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_312),
.Y(n_320)
);

XOR2x1_ASAP7_75t_SL g311 ( 
.A(n_308),
.B(n_292),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_295),
.B(n_286),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_270),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_313),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_297),
.B1(n_299),
.B2(n_295),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_299),
.B(n_309),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_316),
.A2(n_287),
.B(n_306),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_321),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_320),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

NAND4xp25_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_317),
.C(n_311),
.D(n_315),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_326),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_315),
.C(n_310),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_293),
.C(n_324),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_312),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_325),
.Y(n_331)
);


endmodule