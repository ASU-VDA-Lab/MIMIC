module fake_jpeg_163_n_240 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_240);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_240;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_41),
.Y(n_69)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_27),
.B(n_0),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_42),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_1),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_20),
.B(n_2),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_55),
.Y(n_73)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_3),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_3),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_61),
.Y(n_81)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_64),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_36),
.B1(n_35),
.B2(n_18),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_66),
.A2(n_78),
.B1(n_61),
.B2(n_53),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_36),
.B1(n_37),
.B2(n_31),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_75),
.B1(n_76),
.B2(n_42),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_28),
.B1(n_18),
.B2(n_38),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_79),
.B1(n_84),
.B2(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_7),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_31),
.B1(n_23),
.B2(n_28),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_17),
.B1(n_30),
.B2(n_25),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_34),
.B1(n_25),
.B2(n_21),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_34),
.B1(n_25),
.B2(n_17),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_34),
.B1(n_22),
.B2(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_39),
.B(n_4),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_86),
.B(n_88),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_41),
.B(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_49),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_56),
.B(n_4),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_59),
.B1(n_52),
.B2(n_62),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_22),
.B1(n_5),
.B2(n_7),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_62),
.B1(n_63),
.B2(n_12),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_58),
.B(n_4),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_114),
.B(n_119),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_58),
.C(n_59),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_5),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_112),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_83),
.B1(n_91),
.B2(n_81),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_94),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_70),
.A2(n_64),
.B(n_10),
.C(n_11),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_8),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_117),
.Y(n_152)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_82),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_62),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_87),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_10),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_126),
.B(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_53),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_124),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_70),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_82),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_116),
.CI(n_113),
.CON(n_134),
.SN(n_134)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_137),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_138),
.B1(n_145),
.B2(n_150),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_123),
.CI(n_108),
.CON(n_137),
.SN(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_120),
.B1(n_109),
.B2(n_92),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_78),
.B(n_94),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_146),
.B(n_98),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_96),
.B1(n_91),
.B2(n_83),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_88),
.B(n_69),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_68),
.B1(n_85),
.B2(n_69),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_149),
.A2(n_107),
.B1(n_127),
.B2(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_61),
.B1(n_68),
.B2(n_63),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_63),
.B1(n_85),
.B2(n_97),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_87),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_162),
.B1(n_170),
.B2(n_177),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_133),
.A2(n_118),
.B1(n_124),
.B2(n_130),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_178),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_112),
.C(n_86),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_146),
.C(n_148),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_174),
.B(n_145),
.Y(n_180)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_171),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_130),
.B1(n_124),
.B2(n_118),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_98),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_143),
.B(n_138),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_87),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_176),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_136),
.A2(n_98),
.B1(n_100),
.B2(n_111),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_12),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_179),
.B(n_135),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_147),
.C(n_137),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_161),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_172),
.C(n_169),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_152),
.A3(n_132),
.B1(n_134),
.B2(n_137),
.C1(n_178),
.C2(n_167),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_192),
.C(n_171),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_155),
.B(n_134),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_177),
.B(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_158),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_135),
.A3(n_142),
.B1(n_151),
.B2(n_149),
.C1(n_14),
.C2(n_100),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_150),
.B1(n_151),
.B2(n_156),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_194),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_142),
.B1(n_100),
.B2(n_77),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_179),
.B(n_161),
.C(n_176),
.D(n_164),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_199),
.B(n_183),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_184),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_191),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_203),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_206),
.C(n_181),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_207),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_166),
.C(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_208),
.A2(n_209),
.B1(n_195),
.B2(n_182),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_77),
.B1(n_188),
.B2(n_189),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_213),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_217),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_184),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_185),
.C(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_218),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_197),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_183),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_204),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_200),
.B(n_193),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_214),
.B(n_206),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_225),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_204),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_199),
.B(n_212),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_229),
.B(n_200),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_221),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_228),
.B(n_196),
.Y(n_234)
);

OAI221xp5_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_220),
.B1(n_213),
.B2(n_225),
.C(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_219),
.C(n_181),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_233),
.B(n_234),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_235),
.C(n_196),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_238),
.C(n_190),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_235),
.B(n_190),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_77),
.Y(n_240)
);


endmodule