module fake_jpeg_30154_n_494 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_494);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_494;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_48),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_55),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_14),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_63),
.Y(n_115)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_34),
.B(n_13),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_69),
.Y(n_99)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_34),
.B(n_13),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g143 ( 
.A(n_73),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_74),
.B(n_80),
.Y(n_141)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_40),
.B(n_46),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_89),
.Y(n_138)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_90),
.Y(n_144)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_13),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_92),
.Y(n_96)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

BUFx4f_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_26),
.B1(n_23),
.B2(n_43),
.Y(n_103)
);

INVx2_ASAP7_75t_R g94 ( 
.A(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_38),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_100),
.B(n_48),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_47),
.A2(n_20),
.B1(n_35),
.B2(n_29),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_101),
.A2(n_28),
.B1(n_36),
.B2(n_42),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_44),
.B1(n_43),
.B2(n_37),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_102),
.A2(n_105),
.B1(n_122),
.B2(n_31),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_49),
.A2(n_44),
.B1(n_43),
.B2(n_37),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_44),
.B1(n_43),
.B2(n_26),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_110),
.A2(n_127),
.B1(n_130),
.B2(n_41),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_19),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_113),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_18),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_19),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_118),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_18),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_50),
.A2(n_44),
.B1(n_22),
.B2(n_24),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_59),
.A2(n_26),
.B1(n_24),
.B2(n_36),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_73),
.A2(n_36),
.B1(n_28),
.B2(n_24),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_54),
.B(n_46),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_146),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_56),
.B(n_35),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_149),
.A2(n_152),
.B1(n_154),
.B2(n_121),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_144),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_150),
.B(n_160),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_147),
.A2(n_92),
.B1(n_77),
.B2(n_86),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_99),
.B(n_20),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_153),
.B(n_157),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_148),
.A2(n_76),
.B1(n_82),
.B2(n_58),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_115),
.B(n_29),
.Y(n_157)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_74),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_74),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_163),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_96),
.A2(n_79),
.B1(n_87),
.B2(n_85),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_165),
.A2(n_183),
.B1(n_131),
.B2(n_136),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_166),
.A2(n_133),
.B1(n_132),
.B2(n_98),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_96),
.B(n_125),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_171),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_41),
.B1(n_31),
.B2(n_16),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_93),
.C(n_64),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_169),
.B(n_174),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_97),
.B(n_28),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_97),
.B(n_38),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_180),
.Y(n_212)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_138),
.B(n_38),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_126),
.B(n_58),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_185),
.Y(n_221)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_124),
.A2(n_84),
.B1(n_83),
.B2(n_81),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_140),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_138),
.B(n_38),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_192),
.Y(n_234)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_188),
.Y(n_222)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_189),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_41),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_190),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_117),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_191),
.B(n_104),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_108),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_126),
.B(n_66),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_193),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_117),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_194),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_139),
.B(n_65),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_196),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_SL g200 ( 
.A1(n_167),
.A2(n_112),
.B(n_120),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_200),
.B(n_169),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_157),
.C(n_151),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_151),
.B(n_108),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_155),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_233),
.B1(n_235),
.B2(n_183),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_102),
.B(n_121),
.C(n_112),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_204),
.A2(n_123),
.B(n_106),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_211),
.A2(n_176),
.B1(n_185),
.B2(n_163),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_202),
.B1(n_158),
.B2(n_210),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_166),
.A2(n_98),
.B1(n_131),
.B2(n_136),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_171),
.B1(n_192),
.B2(n_173),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_195),
.A2(n_123),
.B(n_137),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_204),
.B(n_218),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_158),
.A2(n_132),
.B1(n_133),
.B2(n_142),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_238),
.A2(n_245),
.B1(n_258),
.B2(n_269),
.Y(n_287)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_228),
.C(n_210),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_248),
.C(n_199),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_241),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_174),
.B(n_190),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_242),
.A2(n_270),
.B(n_53),
.Y(n_293)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_190),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_243),
.B(n_252),
.Y(n_307)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_255),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_228),
.C(n_234),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_204),
.A2(n_165),
.B1(n_174),
.B2(n_180),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_249),
.A2(n_267),
.B1(n_231),
.B2(n_208),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_250),
.A2(n_256),
.B(n_268),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_251),
.B(n_253),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_155),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_186),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_254),
.B(n_261),
.CI(n_263),
.CON(n_282),
.SN(n_282)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_212),
.B(n_184),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_222),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_265),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_216),
.A2(n_156),
.B1(n_164),
.B2(n_142),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_198),
.B(n_150),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_262),
.Y(n_274)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_260),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_212),
.B(n_191),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_205),
.B(n_189),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_177),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_220),
.C(n_198),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_188),
.B1(n_106),
.B2(n_107),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_199),
.A2(n_227),
.B1(n_233),
.B2(n_221),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_227),
.A2(n_176),
.B1(n_187),
.B2(n_175),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_231),
.B1(n_214),
.B2(n_208),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_206),
.B(n_172),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_207),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_275),
.A2(n_293),
.B(n_296),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_221),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_279),
.C(n_283),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_288),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_213),
.C(n_215),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_159),
.B1(n_214),
.B2(n_178),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_284),
.A2(n_292),
.B1(n_297),
.B2(n_299),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_215),
.C(n_207),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_294),
.C(n_300),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_249),
.A2(n_159),
.B1(n_107),
.B2(n_214),
.Y(n_289)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_247),
.A2(n_225),
.B1(n_162),
.B2(n_170),
.Y(n_290)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_290),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_253),
.B(n_194),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_242),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_225),
.B1(n_219),
.B2(n_226),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_219),
.C(n_229),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_250),
.A2(n_229),
.B(n_217),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_256),
.A2(n_226),
.B1(n_179),
.B2(n_217),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_256),
.A2(n_182),
.B1(n_104),
.B2(n_224),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_31),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_16),
.B1(n_170),
.B2(n_162),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_267),
.B1(n_264),
.B2(n_266),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_250),
.C(n_293),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_243),
.B(n_272),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_310),
.A2(n_322),
.B(n_299),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_312),
.B(n_12),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_314),
.B(n_316),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_315),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_274),
.B(n_252),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_259),
.Y(n_317)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_298),
.A2(n_251),
.B(n_257),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_323),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_324),
.A2(n_290),
.B1(n_289),
.B2(n_275),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_307),
.B(n_237),
.Y(n_326)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_295),
.B(n_243),
.Y(n_327)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_328),
.Y(n_363)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_280),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_332),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_262),
.Y(n_331)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_244),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_277),
.B(n_255),
.C(n_237),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_339),
.C(n_286),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_285),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_334),
.Y(n_369)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_303),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_335),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_349)
);

INVx11_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_297),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_303),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_245),
.C(n_260),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_282),
.B(n_239),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_340),
.A2(n_341),
.B1(n_246),
.B2(n_265),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_282),
.B(n_236),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_283),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_343),
.B(n_347),
.Y(n_394)
);

OA22x2_ASAP7_75t_L g345 ( 
.A1(n_308),
.A2(n_287),
.B1(n_302),
.B2(n_305),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_351),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_321),
.A2(n_302),
.B1(n_278),
.B2(n_284),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_312),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_352),
.B(n_365),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_354),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_320),
.A2(n_302),
.B1(n_288),
.B2(n_287),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_291),
.C(n_307),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_356),
.C(n_358),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_294),
.C(n_282),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_357),
.A2(n_367),
.B(n_331),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_333),
.C(n_312),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_321),
.A2(n_292),
.B1(n_304),
.B2(n_301),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_360),
.A2(n_370),
.B1(n_324),
.B2(n_311),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_320),
.A2(n_258),
.B1(n_304),
.B2(n_300),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_362),
.B(n_373),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_309),
.B(n_246),
.C(n_241),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_315),
.C(n_329),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_313),
.A2(n_241),
.B(n_265),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_310),
.A2(n_170),
.B1(n_162),
.B2(n_16),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_371),
.B(n_327),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_311),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_SL g375 ( 
.A(n_361),
.B(n_313),
.C(n_322),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_375),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_364),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_376),
.B(n_377),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_342),
.B(n_317),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_348),
.B(n_314),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_385),
.Y(n_416)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_364),
.Y(n_381)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_309),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_393),
.Y(n_412)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_359),
.Y(n_383)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_383),
.Y(n_422)
);

FAx1_ASAP7_75t_SL g384 ( 
.A(n_355),
.B(n_341),
.CI(n_340),
.CON(n_384),
.SN(n_384)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_391),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_369),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_372),
.B(n_318),
.Y(n_387)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_387),
.Y(n_421)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_388),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_389),
.A2(n_395),
.B1(n_351),
.B2(n_362),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_350),
.B(n_326),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_390),
.B(n_369),
.Y(n_401)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_363),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_398),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_367),
.A2(n_316),
.B1(n_330),
.B2(n_334),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_399),
.C(n_358),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_361),
.A2(n_338),
.B(n_335),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_375),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_352),
.B(n_332),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_343),
.B(n_328),
.C(n_323),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_404),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_403),
.A2(n_374),
.B1(n_400),
.B2(n_389),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_379),
.A2(n_353),
.B1(n_354),
.B2(n_357),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_395),
.A2(n_356),
.B1(n_345),
.B2(n_366),
.Y(n_407)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_407),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_408),
.B(n_409),
.C(n_411),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_345),
.C(n_371),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_374),
.A2(n_349),
.B1(n_360),
.B2(n_345),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_410),
.A2(n_418),
.B1(n_417),
.B2(n_420),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_368),
.C(n_370),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_379),
.A2(n_373),
.B1(n_344),
.B2(n_315),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_418),
.Y(n_438)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_415),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_344),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_336),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_419),
.B(n_378),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_436),
.Y(n_441)
);

AO21x1_ASAP7_75t_L g425 ( 
.A1(n_415),
.A2(n_392),
.B(n_374),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_11),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_384),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_428),
.Y(n_442)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_427),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_403),
.A2(n_400),
.B1(n_382),
.B2(n_396),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_399),
.C(n_386),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_409),
.C(n_411),
.Y(n_443)
);

NOR2x1_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_384),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_439),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_433),
.A2(n_435),
.B1(n_412),
.B2(n_405),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_417),
.A2(n_406),
.B(n_402),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_434),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_406),
.A2(n_386),
.B1(n_336),
.B2(n_398),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_407),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_393),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_11),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_412),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_443),
.B(n_444),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_434),
.B(n_422),
.Y(n_444)
);

AOI21xp33_ASAP7_75t_L g445 ( 
.A1(n_437),
.A2(n_405),
.B(n_419),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_445),
.A2(n_455),
.B(n_425),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_448),
.B(n_450),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_12),
.Y(n_451)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_451),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_432),
.A2(n_11),
.B1(n_10),
.B2(n_2),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_453),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_10),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_454),
.B(n_456),
.C(n_440),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_423),
.B(n_0),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_0),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_461),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_443),
.B(n_432),
.C(n_430),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_2),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_442),
.A2(n_437),
.B(n_438),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_460),
.A2(n_468),
.B(n_469),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_446),
.A2(n_431),
.B1(n_433),
.B2(n_436),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_449),
.A2(n_435),
.B1(n_425),
.B2(n_427),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_466),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_465),
.B(n_441),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_439),
.C(n_428),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_454),
.A2(n_438),
.B(n_424),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_453),
.A2(n_456),
.B(n_441),
.Y(n_469)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_471),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_464),
.A2(n_450),
.B(n_1),
.Y(n_472)
);

AOI32xp33_ASAP7_75t_L g482 ( 
.A1(n_472),
.A2(n_477),
.A3(n_479),
.B1(n_462),
.B2(n_4),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_0),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_474),
.B(n_475),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_459),
.B(n_0),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_1),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_476),
.Y(n_483)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

NOR4xp25_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_462),
.C(n_457),
.D(n_458),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_480),
.B(n_482),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_478),
.B(n_3),
.C(n_5),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_485),
.A2(n_3),
.B(n_6),
.Y(n_489)
);

AOI321xp33_ASAP7_75t_L g487 ( 
.A1(n_484),
.A2(n_479),
.A3(n_473),
.B1(n_472),
.B2(n_7),
.C(n_3),
.Y(n_487)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_487),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_481),
.B(n_473),
.C(n_5),
.Y(n_488)
);

OAI321xp33_ASAP7_75t_L g490 ( 
.A1(n_488),
.A2(n_489),
.A3(n_483),
.B1(n_8),
.B2(n_9),
.C(n_7),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_490),
.A2(n_486),
.B(n_8),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_492),
.B(n_491),
.Y(n_493)
);

AO21x1_ASAP7_75t_L g494 ( 
.A1(n_493),
.A2(n_8),
.B(n_9),
.Y(n_494)
);


endmodule