module fake_ariane_793_n_2618 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_543, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_2618);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_2618;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_2370;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_762;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2599;
wire n_699;
wire n_590;
wire n_727;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_2516;
wire n_2555;
wire n_1969;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1373;
wire n_1081;
wire n_742;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1769;
wire n_1632;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1524;
wire n_1476;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_2606;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_907;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_2425;
wire n_1952;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_2372;
wire n_1806;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_2081;
wire n_937;
wire n_1474;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_2590;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_573;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_217),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_93),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_292),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_37),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_132),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_8),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_397),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_257),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_388),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_213),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_209),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_86),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_358),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_150),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_347),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_480),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_409),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_157),
.Y(n_566)
);

CKINVDCx14_ASAP7_75t_R g567 ( 
.A(n_417),
.Y(n_567)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_209),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_445),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_421),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_288),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_418),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_523),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_467),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_539),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_289),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_99),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_199),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_466),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_403),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_493),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_529),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_99),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_126),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_483),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_35),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_522),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_247),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_530),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_75),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_257),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_504),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_481),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_266),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_440),
.Y(n_595)
);

BUFx5_ASAP7_75t_L g596 ( 
.A(n_21),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_176),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_149),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_322),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_116),
.Y(n_600)
);

CKINVDCx16_ASAP7_75t_R g601 ( 
.A(n_521),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_377),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_528),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_301),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_494),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_118),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_159),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_136),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_174),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_305),
.Y(n_610)
);

BUFx8_ASAP7_75t_SL g611 ( 
.A(n_488),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_309),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_73),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_4),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_526),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_0),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_176),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_189),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_380),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_47),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_492),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_24),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_537),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_312),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_267),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_296),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_25),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_216),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_461),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_474),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_124),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_213),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_540),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_517),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_453),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_543),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_106),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_26),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_305),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_166),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_267),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_422),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_344),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_374),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_148),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_541),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_486),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_471),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_235),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_30),
.Y(n_650)
);

BUFx2_ASAP7_75t_SL g651 ( 
.A(n_166),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_531),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_510),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_98),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_278),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_318),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_274),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_379),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_534),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_336),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_291),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_160),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_345),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_524),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_321),
.Y(n_665)
);

CKINVDCx16_ASAP7_75t_R g666 ( 
.A(n_348),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_69),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_459),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_61),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_533),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_386),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_147),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_169),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_203),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_266),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_35),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_52),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_357),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_463),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_13),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_536),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_143),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_425),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_465),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_68),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_410),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_272),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_39),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_487),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_262),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_89),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_424),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_172),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_14),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_491),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_442),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_154),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_299),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_138),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_146),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_268),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_271),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_104),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_206),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_484),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_384),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_366),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_255),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_121),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_65),
.Y(n_710)
);

BUFx2_ASAP7_75t_SL g711 ( 
.A(n_285),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_200),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_50),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_346),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_446),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_28),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_353),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_26),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_44),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_42),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_406),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_443),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_498),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_67),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_90),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_485),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_329),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_289),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_293),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_398),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_381),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_283),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_297),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_518),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_544),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_532),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_341),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_535),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_407),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_162),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_323),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_331),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_360),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_98),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_170),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_460),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_262),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_61),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_426),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_137),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_25),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_538),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_354),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_525),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_215),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_432),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_110),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_527),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_1),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_330),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_448),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_240),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_255),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_214),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_519),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_78),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_236),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_205),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_502),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_542),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_288),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_428),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_79),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_50),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_239),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_520),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_415),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_52),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_350),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_598),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_598),
.Y(n_781)
);

CKINVDCx14_ASAP7_75t_R g782 ( 
.A(n_567),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_618),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_568),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_618),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_560),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_611),
.Y(n_787)
);

NOR2xp67_ASAP7_75t_L g788 ( 
.A(n_732),
.B(n_0),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_578),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_676),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_676),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_693),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_693),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_699),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_568),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_699),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_601),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_766),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_661),
.Y(n_799)
);

BUFx10_ASAP7_75t_L g800 ( 
.A(n_602),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_596),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_766),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_596),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_611),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_596),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_666),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_596),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_596),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_596),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_596),
.Y(n_810)
);

NOR2xp67_ASAP7_75t_L g811 ( 
.A(n_558),
.B(n_1),
.Y(n_811)
);

NOR2xp67_ASAP7_75t_L g812 ( 
.A(n_558),
.B(n_2),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_560),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_550),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_557),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_559),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_562),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_576),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_571),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_586),
.Y(n_820)
);

INVxp33_ASAP7_75t_L g821 ( 
.A(n_626),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_549),
.Y(n_822)
);

INVxp33_ASAP7_75t_SL g823 ( 
.A(n_658),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_590),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_551),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_591),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_597),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_604),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_606),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_571),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_617),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_754),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_613),
.Y(n_833)
);

BUFx2_ASAP7_75t_SL g834 ( 
.A(n_575),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_622),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_777),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_661),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_567),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_627),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_594),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_723),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_628),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_723),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_661),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_632),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_639),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_641),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_645),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_654),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_655),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_552),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_657),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_669),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_672),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_677),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_690),
.Y(n_856)
);

BUFx5_ASAP7_75t_L g857 ( 
.A(n_561),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_701),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_575),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_704),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_716),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_661),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_594),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_718),
.Y(n_864)
);

INVxp33_ASAP7_75t_L g865 ( 
.A(n_626),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_682),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_575),
.Y(n_867)
);

INVxp67_ASAP7_75t_SL g868 ( 
.A(n_682),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_651),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_719),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_724),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_725),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_682),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_595),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_595),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_744),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_553),
.Y(n_877)
);

BUFx2_ASAP7_75t_SL g878 ( 
.A(n_595),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_751),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_735),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_763),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_764),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_844),
.Y(n_883)
);

NOR2xp67_ASAP7_75t_L g884 ( 
.A(n_787),
.B(n_563),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_866),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_804),
.B(n_555),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_868),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_803),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_805),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_808),
.Y(n_890)
);

CKINVDCx16_ASAP7_75t_R g891 ( 
.A(n_831),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_809),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_782),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_799),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_841),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_810),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_786),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_786),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_869),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_814),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_841),
.Y(n_901)
);

INVxp67_ASAP7_75t_SL g902 ( 
.A(n_821),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_819),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_816),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_819),
.Y(n_905)
);

NOR2xp67_ASAP7_75t_L g906 ( 
.A(n_838),
.B(n_564),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_782),
.B(n_572),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_817),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_818),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_840),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_843),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_843),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_838),
.B(n_574),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_789),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_840),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_813),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_834),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_L g918 ( 
.A(n_859),
.B(n_570),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_797),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_797),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_830),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_806),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_795),
.B(n_617),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_801),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_820),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_806),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_859),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_823),
.B(n_580),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_867),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_863),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_824),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_867),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_826),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_874),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_827),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_874),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_832),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_878),
.Y(n_938)
);

XNOR2x1_ASAP7_75t_L g939 ( 
.A(n_832),
.B(n_608),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_828),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_875),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_875),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_880),
.Y(n_943)
);

INVxp33_ASAP7_75t_SL g944 ( 
.A(n_784),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_880),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_829),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_833),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_902),
.B(n_815),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_900),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_924),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_904),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_897),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_924),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_928),
.B(n_784),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_908),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_899),
.B(n_836),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_909),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_888),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_913),
.B(n_823),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_895),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_889),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_925),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_894),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_923),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_931),
.B(n_821),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_933),
.B(n_865),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_935),
.B(n_865),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_914),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_927),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_890),
.B(n_836),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_940),
.Y(n_971)
);

OA21x2_ASAP7_75t_L g972 ( 
.A1(n_892),
.A2(n_807),
.B(n_801),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_946),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_947),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_896),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_929),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_932),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_883),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_885),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_894),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_887),
.B(n_802),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_901),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_894),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_907),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_906),
.A2(n_807),
.B(n_799),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_918),
.B(n_857),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_917),
.B(n_815),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_893),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_911),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_938),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_897),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_884),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_893),
.B(n_780),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_934),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_912),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_886),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_937),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_936),
.B(n_835),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_945),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_941),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_942),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_898),
.Y(n_1002)
);

AND3x2_ASAP7_75t_L g1003 ( 
.A(n_891),
.B(n_877),
.C(n_825),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_943),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_919),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_944),
.B(n_857),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_920),
.Y(n_1007)
);

NAND3xp33_ASAP7_75t_L g1008 ( 
.A(n_922),
.B(n_851),
.C(n_822),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_926),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_944),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_939),
.B(n_781),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_939),
.B(n_783),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_916),
.B(n_839),
.Y(n_1013)
);

NOR2x1_ASAP7_75t_L g1014 ( 
.A(n_916),
.B(n_842),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_921),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_930),
.Y(n_1016)
);

XNOR2xp5_ASAP7_75t_L g1017 ( 
.A(n_921),
.B(n_667),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_930),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_898),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_903),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_903),
.B(n_800),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_905),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_905),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_910),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_910),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_915),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_915),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_895),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_900),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_900),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_900),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_902),
.B(n_857),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_914),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_924),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_900),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_924),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_972),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_972),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_972),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1034),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_984),
.B(n_857),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_998),
.B(n_800),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1034),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_958),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_950),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_958),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_965),
.B(n_800),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_998),
.B(n_788),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_950),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_961),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_961),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_1016),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_975),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_965),
.B(n_785),
.Y(n_1054)
);

BUFx4f_ASAP7_75t_L g1055 ( 
.A(n_1010),
.Y(n_1055)
);

BUFx8_ASAP7_75t_SL g1056 ( 
.A(n_988),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_1032),
.A2(n_623),
.B(n_621),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_975),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_983),
.Y(n_1059)
);

AND3x2_ASAP7_75t_L g1060 ( 
.A(n_982),
.B(n_708),
.C(n_667),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_959),
.B(n_708),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_985),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_950),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_959),
.B(n_556),
.C(n_554),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_985),
.Y(n_1065)
);

AND3x2_ASAP7_75t_L g1066 ( 
.A(n_989),
.B(n_733),
.C(n_767),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_954),
.B(n_733),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_956),
.B(n_566),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_963),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_963),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_948),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_966),
.B(n_790),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_998),
.B(n_577),
.Y(n_1073)
);

BUFx10_ASAP7_75t_L g1074 ( 
.A(n_1007),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_1016),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_950),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_963),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_948),
.B(n_1006),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_978),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_953),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_953),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_953),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_953),
.Y(n_1083)
);

OAI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_969),
.A2(n_976),
.B1(n_977),
.B2(n_1007),
.Y(n_1084)
);

INVxp33_ASAP7_75t_L g1085 ( 
.A(n_1017),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_966),
.B(n_791),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_963),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_994),
.B(n_583),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_980),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_980),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_980),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_980),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_949),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1036),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_948),
.B(n_857),
.Y(n_1095)
);

AO21x2_ASAP7_75t_L g1096 ( 
.A1(n_986),
.A2(n_970),
.B(n_955),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_1036),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_951),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_994),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_957),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_L g1101 ( 
.A1(n_962),
.A2(n_634),
.B(n_629),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_971),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_994),
.B(n_584),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_973),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_994),
.B(n_999),
.Y(n_1105)
);

OAI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_969),
.A2(n_811),
.B1(n_812),
.B2(n_767),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_974),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1029),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1000),
.B(n_588),
.Y(n_1109)
);

CKINVDCx6p67_ASAP7_75t_R g1110 ( 
.A(n_988),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_964),
.A2(n_857),
.B1(n_653),
.B2(n_660),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_967),
.B(n_857),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1030),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1031),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1035),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_979),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_967),
.B(n_569),
.Y(n_1117)
);

AOI21x1_ASAP7_75t_L g1118 ( 
.A1(n_996),
.A2(n_668),
.B(n_646),
.Y(n_1118)
);

CKINVDCx6p67_ASAP7_75t_R g1119 ( 
.A(n_1026),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_981),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_981),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_993),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_987),
.B(n_635),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_990),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_1005),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_992),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_L g1127 ( 
.A1(n_993),
.A2(n_696),
.B(n_671),
.Y(n_1127)
);

BUFx8_ASAP7_75t_SL g1128 ( 
.A(n_952),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_964),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_987),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_999),
.B(n_600),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1013),
.B(n_792),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_987),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_997),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_997),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1008),
.A2(n_726),
.B(n_705),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1001),
.A2(n_736),
.B(n_734),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1011),
.B(n_607),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1004),
.B(n_1009),
.Y(n_1139)
);

INVx5_ASAP7_75t_L g1140 ( 
.A(n_999),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1013),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1013),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1026),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1011),
.Y(n_1144)
);

CKINVDCx6p67_ASAP7_75t_R g1145 ( 
.A(n_1010),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_968),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1012),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_968),
.B(n_793),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1012),
.B(n_609),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1009),
.Y(n_1150)
);

INVxp33_ASAP7_75t_SL g1151 ( 
.A(n_976),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1014),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1010),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1010),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_999),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1005),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1005),
.Y(n_1157)
);

AND3x2_ASAP7_75t_L g1158 ( 
.A(n_960),
.B(n_846),
.C(n_845),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1005),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_995),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1003),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1015),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_977),
.Y(n_1163)
);

NOR2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1033),
.B(n_876),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1015),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1033),
.B(n_610),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1018),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1018),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1018),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1018),
.Y(n_1170)
);

INVx11_ASAP7_75t_L g1171 ( 
.A(n_1028),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1027),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1027),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1027),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1050),
.Y(n_1175)
);

INVx4_ASAP7_75t_L g1176 ( 
.A(n_1145),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1171),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1056),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1050),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1040),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1056),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_1145),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1045),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1116),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1067),
.B(n_1021),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1049),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1116),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1055),
.B(n_1023),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1045),
.Y(n_1189)
);

AND2x6_ASAP7_75t_L g1190 ( 
.A(n_1099),
.B(n_1027),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1071),
.B(n_1068),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1071),
.B(n_778),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1171),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_1099),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1040),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1061),
.B(n_1020),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1052),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1151),
.B(n_1022),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_1075),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1079),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1162),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1162),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1045),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1165),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1125),
.B(n_1023),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1128),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1151),
.B(n_1146),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1165),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1148),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1043),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1117),
.B(n_612),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1134),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1134),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1093),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1093),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1055),
.B(n_1023),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1100),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1128),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1055),
.B(n_1025),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1110),
.Y(n_1220)
);

NAND2xp33_ASAP7_75t_L g1221 ( 
.A(n_1099),
.B(n_614),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1045),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1140),
.B(n_1025),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1140),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1110),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1047),
.B(n_1025),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1099),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1049),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1043),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1100),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1107),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1148),
.Y(n_1232)
);

INVx4_ASAP7_75t_SL g1233 ( 
.A(n_1099),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1074),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1140),
.B(n_1024),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1107),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1084),
.B(n_1019),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1140),
.B(n_616),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1113),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1044),
.Y(n_1240)
);

AND2x6_ASAP7_75t_L g1241 ( 
.A(n_1125),
.B(n_565),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1143),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1140),
.B(n_1139),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1074),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1049),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1135),
.B(n_620),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1074),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1113),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1047),
.B(n_952),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1122),
.B(n_625),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1144),
.B(n_991),
.Y(n_1251)
);

INVx1_ASAP7_75t_SL g1252 ( 
.A(n_1119),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1122),
.B(n_1160),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1044),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1144),
.B(n_991),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1135),
.B(n_631),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1160),
.B(n_1002),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1078),
.B(n_637),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1172),
.B(n_1002),
.Y(n_1259)
);

INVx4_ASAP7_75t_L g1260 ( 
.A(n_1119),
.Y(n_1260)
);

INVx4_ASAP7_75t_L g1261 ( 
.A(n_1172),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1114),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1083),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1141),
.B(n_711),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1083),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1163),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1114),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1153),
.B(n_638),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1098),
.Y(n_1269)
);

OAI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1138),
.A2(n_640),
.B1(n_650),
.B2(n_649),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1163),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1046),
.Y(n_1272)
);

AND2x6_ASAP7_75t_L g1273 ( 
.A(n_1062),
.B(n_565),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1046),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1153),
.B(n_847),
.Y(n_1275)
);

NOR3xp33_ASAP7_75t_L g1276 ( 
.A(n_1073),
.B(n_673),
.C(n_662),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1163),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1051),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1153),
.B(n_848),
.Y(n_1279)
);

AO22x2_ASAP7_75t_L g1280 ( 
.A1(n_1147),
.A2(n_882),
.B1(n_850),
.B2(n_852),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1098),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1154),
.B(n_674),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1083),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1045),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1097),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1147),
.B(n_794),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1051),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1154),
.B(n_675),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1135),
.B(n_680),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1102),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1164),
.B(n_860),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1141),
.B(n_849),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1053),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1155),
.B(n_685),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1120),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1102),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1053),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1108),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1108),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_1120),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1115),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1155),
.B(n_687),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1097),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1161),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1121),
.B(n_796),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1142),
.B(n_853),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1059),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1097),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1167),
.B(n_688),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1158),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1115),
.Y(n_1311)
);

NAND2xp33_ASAP7_75t_SL g1312 ( 
.A(n_1156),
.B(n_691),
.Y(n_1312)
);

AND2x6_ASAP7_75t_L g1313 ( 
.A(n_1062),
.B(n_582),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1063),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1167),
.B(n_694),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1104),
.A2(n_698),
.B1(n_702),
.B2(n_700),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1058),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1121),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1157),
.B(n_703),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1161),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1168),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1132),
.B(n_1149),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1077),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1058),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1168),
.B(n_710),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1169),
.B(n_1170),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1104),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1059),
.Y(n_1328)
);

CKINVDCx6p67_ASAP7_75t_R g1329 ( 
.A(n_1042),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1169),
.B(n_712),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_1094),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1104),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1094),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1157),
.B(n_713),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1077),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1132),
.B(n_798),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1063),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1133),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1076),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1076),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1170),
.B(n_720),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1173),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1133),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1159),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1080),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1142),
.A2(n_735),
.B1(n_617),
.B2(n_697),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1159),
.B(n_729),
.Y(n_1347)
);

BUFx4f_ASAP7_75t_L g1348 ( 
.A(n_1161),
.Y(n_1348)
);

BUFx10_ASAP7_75t_L g1349 ( 
.A(n_1109),
.Y(n_1349)
);

BUFx10_ASAP7_75t_L g1350 ( 
.A(n_1060),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1173),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1080),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1124),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1065),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1130),
.A2(n_735),
.B1(n_697),
.B2(n_740),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1156),
.B(n_745),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1081),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1054),
.B(n_854),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1081),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1065),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1082),
.Y(n_1361)
);

INVx4_ASAP7_75t_L g1362 ( 
.A(n_1077),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1130),
.A2(n_697),
.B1(n_748),
.B2(n_747),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1112),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1037),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1082),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1037),
.Y(n_1367)
);

AND2x6_ASAP7_75t_L g1368 ( 
.A(n_1038),
.B(n_582),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1038),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1089),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1054),
.B(n_750),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1089),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1150),
.B(n_755),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1090),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1090),
.Y(n_1375)
);

OR2x6_ASAP7_75t_L g1376 ( 
.A(n_1174),
.B(n_855),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1129),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1307),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1214),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1215),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1196),
.B(n_1129),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1322),
.B(n_1300),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1217),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1328),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1175),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1230),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1349),
.B(n_1197),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1231),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1185),
.B(n_1085),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1236),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1239),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1248),
.A2(n_1064),
.B1(n_1111),
.B2(n_1041),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1318),
.B(n_1072),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1349),
.B(n_1106),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1260),
.B(n_1176),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1175),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1358),
.B(n_1072),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1249),
.B(n_1086),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1257),
.A2(n_1198),
.B1(n_1237),
.B2(n_1232),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1199),
.B(n_1174),
.Y(n_1400)
);

NAND2xp33_ASAP7_75t_SL g1401 ( 
.A(n_1277),
.B(n_1105),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1295),
.B(n_1209),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1191),
.A2(n_1095),
.B(n_1126),
.C(n_1086),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1179),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1253),
.B(n_1048),
.C(n_1088),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1262),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1207),
.B(n_1166),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1251),
.B(n_1123),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1255),
.B(n_1103),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1226),
.B(n_1152),
.Y(n_1410)
);

NAND2x1_ASAP7_75t_L g1411 ( 
.A(n_1224),
.B(n_1091),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1336),
.B(n_1152),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1292),
.B(n_1096),
.Y(n_1413)
);

AND2x4_ASAP7_75t_SL g1414 ( 
.A(n_1176),
.B(n_1091),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1292),
.B(n_1096),
.Y(n_1415)
);

NOR3xp33_ASAP7_75t_L g1416 ( 
.A(n_1270),
.B(n_1131),
.C(n_1127),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1242),
.A2(n_1066),
.B1(n_1070),
.B2(n_1069),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1206),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1177),
.A2(n_1070),
.B1(n_1087),
.B2(n_1069),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1348),
.B(n_1092),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1179),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1306),
.B(n_1096),
.Y(n_1422)
);

AND2x6_ASAP7_75t_L g1423 ( 
.A(n_1327),
.B(n_1039),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1193),
.B(n_1087),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1259),
.A2(n_1280),
.B1(n_1306),
.B2(n_1187),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1267),
.B(n_1092),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1200),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1212),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1259),
.B(n_856),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1280),
.B(n_858),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1371),
.B(n_861),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1264),
.B(n_864),
.Y(n_1432)
);

NOR3xp33_ASAP7_75t_L g1433 ( 
.A(n_1276),
.B(n_1127),
.C(n_1136),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1213),
.Y(n_1434)
);

BUFx10_ASAP7_75t_L g1435 ( 
.A(n_1178),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1180),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1266),
.B(n_1136),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1348),
.B(n_1137),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1182),
.B(n_1137),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1286),
.B(n_870),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1205),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1260),
.B(n_1182),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1305),
.B(n_871),
.Y(n_1443)
);

NAND2xp33_ASAP7_75t_L g1444 ( 
.A(n_1194),
.B(n_1039),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1353),
.B(n_872),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1194),
.B(n_1118),
.Y(n_1446)
);

OAI22x1_ASAP7_75t_SL g1447 ( 
.A1(n_1181),
.A2(n_759),
.B1(n_762),
.B2(n_757),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1195),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1184),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_L g1450 ( 
.A(n_1194),
.B(n_768),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1211),
.B(n_1252),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1291),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1320),
.B(n_1118),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1275),
.B(n_879),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_1220),
.Y(n_1455)
);

NAND2x1p5_ASAP7_75t_L g1456 ( 
.A(n_1227),
.B(n_1101),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1264),
.B(n_1057),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1210),
.Y(n_1458)
);

A2O1A1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1332),
.A2(n_738),
.B(n_739),
.C(n_737),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1229),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1227),
.B(n_771),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1227),
.B(n_1205),
.Y(n_1462)
);

A2O1A1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1309),
.A2(n_746),
.B(n_756),
.C(n_741),
.Y(n_1463)
);

AO22x2_ASAP7_75t_L g1464 ( 
.A1(n_1269),
.A2(n_881),
.B1(n_681),
.B2(n_686),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1281),
.A2(n_774),
.B1(n_775),
.B2(n_773),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1240),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1225),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1275),
.B(n_1101),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1354),
.A2(n_1360),
.B1(n_1324),
.B2(n_1317),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1279),
.B(n_1290),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1218),
.A2(n_709),
.B1(n_728),
.B2(n_682),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1329),
.B(n_1057),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1279),
.B(n_799),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1296),
.B(n_709),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1258),
.B(n_573),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1298),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1261),
.B(n_579),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1254),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1377),
.B(n_581),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1299),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1301),
.B(n_709),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1311),
.A2(n_728),
.B1(n_709),
.B2(n_761),
.Y(n_1482)
);

AND2x2_ASAP7_75t_SL g1483 ( 
.A(n_1261),
.B(n_1221),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1272),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_SL g1485 ( 
.A(n_1234),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1274),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1244),
.B(n_752),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1201),
.Y(n_1488)
);

NAND3xp33_ASAP7_75t_L g1489 ( 
.A(n_1364),
.B(n_728),
.C(n_769),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1190),
.B(n_728),
.Y(n_1490)
);

BUFx5_ASAP7_75t_L g1491 ( 
.A(n_1354),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_SL g1492 ( 
.A(n_1247),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1202),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1190),
.B(n_837),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1190),
.B(n_837),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1271),
.B(n_758),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1190),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1233),
.B(n_1224),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1376),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1188),
.B(n_585),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1315),
.B(n_862),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1338),
.A2(n_770),
.B1(n_670),
.B2(n_686),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1216),
.B(n_587),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1278),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1219),
.B(n_589),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1233),
.B(n_779),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1312),
.A2(n_593),
.B1(n_599),
.B2(n_592),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1287),
.Y(n_1508)
);

INVx8_ASAP7_75t_L g1509 ( 
.A(n_1241),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1204),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1208),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1364),
.A2(n_681),
.B(n_670),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1372),
.B(n_727),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1250),
.B(n_603),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1293),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1373),
.B(n_605),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1297),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1360),
.A2(n_753),
.B(n_743),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1333),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1246),
.A2(n_753),
.B(n_743),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1325),
.B(n_862),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1365),
.B(n_873),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1365),
.B(n_873),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1330),
.B(n_2),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1372),
.B(n_760),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1341),
.B(n_3),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1192),
.B(n_3),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1343),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1376),
.B(n_4),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1374),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1183),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1321),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1339),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_SL g1534 ( 
.A(n_1241),
.B(n_619),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1372),
.B(n_776),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1316),
.B(n_624),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1350),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1375),
.B(n_772),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1342),
.B(n_1367),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1367),
.B(n_5),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1304),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1183),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1351),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1310),
.A2(n_749),
.B1(n_615),
.B2(n_633),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1223),
.B(n_630),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1357),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1369),
.B(n_5),
.Y(n_1547)
);

NOR3xp33_ASAP7_75t_L g1548 ( 
.A(n_1282),
.B(n_765),
.C(n_642),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1359),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1361),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1303),
.B(n_636),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1303),
.B(n_643),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1308),
.B(n_644),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1369),
.B(n_6),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1350),
.A2(n_749),
.B1(n_615),
.B2(n_648),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1375),
.B(n_647),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1326),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1331),
.B(n_6),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1308),
.B(n_652),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1375),
.B(n_656),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1241),
.B(n_7),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1241),
.B(n_7),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1256),
.B(n_8),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1323),
.B(n_659),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1370),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1370),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1289),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_L g1568 ( 
.A(n_1344),
.B(n_663),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1288),
.B(n_664),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1346),
.B(n_9),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1356),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1243),
.B(n_749),
.C(n_615),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1363),
.B(n_10),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1323),
.B(n_11),
.Y(n_1574)
);

NOR4xp25_ASAP7_75t_SL g1575 ( 
.A(n_1238),
.B(n_1235),
.C(n_1268),
.D(n_1294),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1355),
.A2(n_615),
.B1(n_749),
.B2(n_678),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1186),
.A2(n_679),
.B(n_683),
.C(n_665),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1302),
.A2(n_689),
.B1(n_692),
.B2(n_684),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1319),
.A2(n_706),
.B1(n_707),
.B2(n_695),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1334),
.B(n_714),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1314),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1314),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1314),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1335),
.B(n_12),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1335),
.B(n_715),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1362),
.B(n_12),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1362),
.B(n_13),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1395),
.B(n_1186),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1397),
.B(n_1337),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1399),
.B(n_1347),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1395),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1378),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1398),
.B(n_1337),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1389),
.A2(n_1313),
.B1(n_1273),
.B2(n_1245),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1429),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1451),
.B(n_1285),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1418),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1453),
.B(n_1285),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1382),
.B(n_1408),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1435),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1536),
.A2(n_1313),
.B1(n_1273),
.B2(n_1245),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1509),
.B(n_1337),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1499),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1443),
.B(n_1340),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1384),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1427),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1587),
.B(n_1228),
.Y(n_1607)
);

INVx5_ASAP7_75t_L g1608 ( 
.A(n_1509),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1587),
.B(n_1228),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1409),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1435),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1394),
.B(n_1340),
.Y(n_1612)
);

AO22x1_ASAP7_75t_L g1613 ( 
.A1(n_1573),
.A2(n_1537),
.B1(n_1442),
.B2(n_1472),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1379),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1524),
.A2(n_1526),
.B1(n_1407),
.B2(n_1405),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1440),
.B(n_1340),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1444),
.A2(n_1284),
.B(n_1265),
.Y(n_1617)
);

O2A1O1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1463),
.A2(n_1265),
.B(n_1283),
.C(n_1263),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1528),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1380),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1383),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1455),
.A2(n_1273),
.B1(n_1313),
.B2(n_1283),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1442),
.B(n_1263),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1405),
.A2(n_1284),
.B1(n_1189),
.B2(n_1203),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1386),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1393),
.B(n_1345),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1483),
.B(n_1183),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1388),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1390),
.Y(n_1629)
);

NOR3xp33_ASAP7_75t_SL g1630 ( 
.A(n_1401),
.B(n_721),
.C(n_717),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1498),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1436),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1402),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1391),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1567),
.A2(n_1563),
.B1(n_1431),
.B2(n_1381),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1454),
.B(n_1345),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1410),
.B(n_1345),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1412),
.B(n_1352),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1541),
.Y(n_1639)
);

CKINVDCx11_ASAP7_75t_R g1640 ( 
.A(n_1441),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1406),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1467),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1428),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1498),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1441),
.A2(n_1313),
.B1(n_1273),
.B2(n_1352),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1557),
.B(n_1352),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1471),
.A2(n_730),
.B1(n_731),
.B2(n_722),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1532),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1452),
.A2(n_1366),
.B1(n_1368),
.B2(n_1189),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1434),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1449),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1485),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1425),
.B(n_1366),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1543),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1531),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1387),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1430),
.B(n_1366),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1385),
.B(n_1189),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1396),
.B(n_1203),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1531),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1476),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1414),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1424),
.B(n_1203),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1432),
.B(n_14),
.Y(n_1664)
);

INVx4_ASAP7_75t_L g1665 ( 
.A(n_1485),
.Y(n_1665)
);

NAND2xp33_ASAP7_75t_SL g1666 ( 
.A(n_1492),
.B(n_1222),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1529),
.B(n_1222),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1582),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1480),
.Y(n_1669)
);

BUFx3_ASAP7_75t_L g1670 ( 
.A(n_1583),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1488),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1404),
.B(n_1222),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1421),
.B(n_1368),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_R g1674 ( 
.A(n_1492),
.B(n_1368),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1448),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1546),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1447),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1581),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1531),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1493),
.Y(n_1680)
);

A2O1A1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1416),
.A2(n_1520),
.B(n_1403),
.C(n_1527),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1542),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1510),
.Y(n_1683)
);

BUFx12f_ASAP7_75t_L g1684 ( 
.A(n_1542),
.Y(n_1684)
);

NOR2x1_ASAP7_75t_L g1685 ( 
.A(n_1450),
.B(n_1368),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1514),
.B(n_742),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1417),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1462),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1570),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1458),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1511),
.Y(n_1691)
);

NAND2x2_ASAP7_75t_L g1692 ( 
.A(n_1574),
.B(n_15),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1460),
.Y(n_1693)
);

NOR3xp33_ASAP7_75t_L g1694 ( 
.A(n_1571),
.B(n_16),
.C(n_17),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1437),
.A2(n_1479),
.B1(n_1475),
.B2(n_1569),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1466),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1516),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1470),
.B(n_18),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1445),
.B(n_19),
.Y(n_1699)
);

INVx8_ASAP7_75t_L g1700 ( 
.A(n_1509),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1478),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1497),
.B(n_548),
.Y(n_1702)
);

INVx5_ASAP7_75t_L g1703 ( 
.A(n_1423),
.Y(n_1703)
);

NOR3xp33_ASAP7_75t_SL g1704 ( 
.A(n_1487),
.B(n_20),
.C(n_21),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1539),
.B(n_22),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1473),
.B(n_22),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1515),
.B(n_23),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1420),
.B(n_547),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1423),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1517),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1519),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1530),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1464),
.B(n_23),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1534),
.B(n_24),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1400),
.B(n_311),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1533),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1549),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1464),
.B(n_27),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1465),
.B(n_1580),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1534),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1496),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1484),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1568),
.B(n_29),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1486),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1550),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1584),
.Y(n_1726)
);

NAND3xp33_ASAP7_75t_SL g1727 ( 
.A(n_1575),
.B(n_30),
.C(n_31),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1504),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1508),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1500),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1426),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1469),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1419),
.B(n_32),
.Y(n_1733)
);

OR2x6_ASAP7_75t_L g1734 ( 
.A(n_1461),
.B(n_33),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1551),
.B(n_34),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1552),
.B(n_34),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1469),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1540),
.Y(n_1738)
);

AND2x6_ASAP7_75t_L g1739 ( 
.A(n_1561),
.B(n_1562),
.Y(n_1739)
);

NOR2x2_ASAP7_75t_L g1740 ( 
.A(n_1565),
.B(n_36),
.Y(n_1740)
);

AND2x4_ASAP7_75t_SL g1741 ( 
.A(n_1566),
.B(n_313),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1558),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1506),
.Y(n_1743)
);

A2O1A1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1520),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1553),
.B(n_38),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1559),
.B(n_39),
.Y(n_1746)
);

INVx4_ASAP7_75t_L g1747 ( 
.A(n_1423),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1413),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1503),
.A2(n_1505),
.B1(n_1545),
.B2(n_1507),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1415),
.B(n_40),
.Y(n_1750)
);

BUFx4f_ASAP7_75t_L g1751 ( 
.A(n_1423),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1586),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1422),
.B(n_41),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1494),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1490),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1457),
.B(n_43),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1547),
.B(n_43),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1491),
.B(n_44),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1554),
.B(n_45),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1555),
.B(n_45),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1522),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1456),
.Y(n_1762)
);

NOR3xp33_ASAP7_75t_SL g1763 ( 
.A(n_1477),
.B(n_46),
.C(n_47),
.Y(n_1763)
);

AND3x1_ASAP7_75t_L g1764 ( 
.A(n_1548),
.B(n_46),
.C(n_48),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1522),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1523),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1491),
.B(n_48),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1523),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1512),
.B(n_49),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1513),
.B(n_546),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1491),
.B(n_49),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1411),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1491),
.B(n_51),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1502),
.B(n_51),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1501),
.B(n_53),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1512),
.B(n_53),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1521),
.B(n_54),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_1575),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1576),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1495),
.Y(n_1780)
);

OAI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1392),
.A2(n_55),
.B(n_56),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1474),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1456),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1481),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1491),
.B(n_57),
.Y(n_1785)
);

NAND2x1p5_ASAP7_75t_L g1786 ( 
.A(n_1608),
.B(n_1525),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1695),
.B(n_1438),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1681),
.A2(n_1518),
.B(n_1439),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1749),
.B(n_1468),
.Y(n_1789)
);

CKINVDCx10_ASAP7_75t_R g1790 ( 
.A(n_1734),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1610),
.B(n_1535),
.Y(n_1791)
);

O2A1O1Ixp33_ASAP7_75t_L g1792 ( 
.A1(n_1615),
.A2(n_1459),
.B(n_1392),
.C(n_1577),
.Y(n_1792)
);

O2A1O1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1781),
.A2(n_1518),
.B(n_1433),
.C(n_1538),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1616),
.B(n_1556),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1751),
.A2(n_1446),
.B(n_1489),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1606),
.Y(n_1796)
);

BUFx12f_ASAP7_75t_L g1797 ( 
.A(n_1652),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1686),
.B(n_1560),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1635),
.B(n_1489),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1639),
.B(n_1564),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1751),
.A2(n_1572),
.B(n_1585),
.Y(n_1801)
);

O2A1O1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1590),
.A2(n_1579),
.B(n_1578),
.C(n_1544),
.Y(n_1802)
);

XOR2x2_ASAP7_75t_SL g1803 ( 
.A(n_1740),
.B(n_57),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1599),
.B(n_58),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1595),
.B(n_58),
.Y(n_1805)
);

O2A1O1Ixp5_ASAP7_75t_L g1806 ( 
.A1(n_1714),
.A2(n_1572),
.B(n_1482),
.C(n_62),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1617),
.A2(n_59),
.B(n_60),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1607),
.A2(n_59),
.B(n_60),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1664),
.B(n_62),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1726),
.B(n_63),
.Y(n_1810)
);

OR2x6_ASAP7_75t_SL g1811 ( 
.A(n_1778),
.B(n_1677),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1633),
.B(n_63),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1591),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1719),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1609),
.A2(n_64),
.B(n_66),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1597),
.B(n_67),
.Y(n_1816)
);

OR2x6_ASAP7_75t_L g1817 ( 
.A(n_1700),
.B(n_1613),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1591),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1614),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1598),
.A2(n_68),
.B(n_69),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1713),
.A2(n_1718),
.B1(n_1694),
.B2(n_1764),
.C(n_1736),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1663),
.B(n_70),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1676),
.B(n_1593),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1591),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1721),
.B(n_70),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1640),
.B(n_71),
.Y(n_1826)
);

OAI22x1_ASAP7_75t_L g1827 ( 
.A1(n_1697),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1827)
);

OA22x2_ASAP7_75t_L g1828 ( 
.A1(n_1687),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1647),
.A2(n_77),
.B1(n_74),
.B2(n_76),
.Y(n_1829)
);

AOI21x1_ASAP7_75t_L g1830 ( 
.A1(n_1756),
.A2(n_315),
.B(n_314),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1619),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1727),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1832)
);

OAI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1735),
.A2(n_79),
.B(n_80),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1700),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1703),
.A2(n_80),
.B(n_81),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1703),
.A2(n_81),
.B(n_82),
.Y(n_1836)
);

A2O1A1Ixp33_ASAP7_75t_L g1837 ( 
.A1(n_1745),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1604),
.B(n_83),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_1684),
.Y(n_1839)
);

AOI22x1_ASAP7_75t_L g1840 ( 
.A1(n_1642),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_R g1841 ( 
.A(n_1666),
.B(n_316),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1731),
.B(n_85),
.Y(n_1842)
);

O2A1O1Ixp33_ASAP7_75t_SL g1843 ( 
.A1(n_1746),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1760),
.A2(n_90),
.B1(n_87),
.B2(n_88),
.Y(n_1844)
);

OAI21x1_ASAP7_75t_L g1845 ( 
.A1(n_1782),
.A2(n_319),
.B(n_317),
.Y(n_1845)
);

A2O1A1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1730),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1703),
.A2(n_91),
.B(n_92),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1732),
.A2(n_94),
.B(n_95),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1742),
.B(n_94),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1603),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_SL g1851 ( 
.A(n_1665),
.B(n_320),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1770),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1752),
.B(n_96),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1737),
.A2(n_97),
.B(n_100),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1620),
.B(n_100),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1769),
.A2(n_101),
.B(n_102),
.Y(n_1856)
);

INVx5_ASAP7_75t_L g1857 ( 
.A(n_1709),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1596),
.B(n_101),
.Y(n_1858)
);

AOI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1784),
.A2(n_325),
.B(n_324),
.Y(n_1859)
);

NOR3xp33_ASAP7_75t_L g1860 ( 
.A(n_1744),
.B(n_1733),
.C(n_1757),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1621),
.B(n_1625),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1653),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1628),
.B(n_103),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1678),
.B(n_105),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1629),
.B(n_105),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_R g1866 ( 
.A(n_1631),
.B(n_326),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1709),
.B(n_106),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1592),
.Y(n_1868)
);

BUFx4f_ASAP7_75t_L g1869 ( 
.A(n_1655),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1634),
.B(n_107),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1631),
.B(n_107),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1588),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1709),
.B(n_1622),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1648),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1655),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1776),
.A2(n_108),
.B(n_109),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1656),
.B(n_108),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1720),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1605),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1654),
.Y(n_1880)
);

O2A1O1Ixp33_ASAP7_75t_L g1881 ( 
.A1(n_1759),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1641),
.B(n_112),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1774),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1594),
.B(n_114),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1643),
.B(n_115),
.Y(n_1885)
);

INVx6_ASAP7_75t_L g1886 ( 
.A(n_1665),
.Y(n_1886)
);

AOI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1747),
.A2(n_116),
.B(n_117),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1702),
.B(n_117),
.Y(n_1888)
);

NOR2x1_ASAP7_75t_L g1889 ( 
.A(n_1785),
.B(n_118),
.Y(n_1889)
);

NOR3xp33_ASAP7_75t_L g1890 ( 
.A(n_1689),
.B(n_119),
.C(n_120),
.Y(n_1890)
);

A2O1A1Ixp33_ASAP7_75t_SL g1891 ( 
.A1(n_1772),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1650),
.B(n_122),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1747),
.A2(n_122),
.B(n_123),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1588),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1646),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1632),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1601),
.A2(n_1618),
.B(n_1627),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1758),
.A2(n_1771),
.B(n_1767),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1773),
.A2(n_123),
.B(n_124),
.Y(n_1899)
);

A2O1A1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1770),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_1900)
);

NOR2xp67_ASAP7_75t_L g1901 ( 
.A(n_1600),
.B(n_327),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1667),
.B(n_125),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1675),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1624),
.A2(n_127),
.B(n_128),
.Y(n_1904)
);

INVxp67_ASAP7_75t_L g1905 ( 
.A(n_1637),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1738),
.A2(n_1777),
.B(n_1702),
.Y(n_1906)
);

AOI21x1_ASAP7_75t_L g1907 ( 
.A1(n_1750),
.A2(n_332),
.B(n_328),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1705),
.B(n_128),
.Y(n_1908)
);

AOI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1765),
.A2(n_1766),
.B(n_1753),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1779),
.A2(n_129),
.B(n_130),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_SL g1911 ( 
.A1(n_1723),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1911)
);

BUFx2_ASAP7_75t_SL g1912 ( 
.A(n_1611),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1651),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1626),
.B(n_131),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1674),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1612),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1661),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1589),
.A2(n_133),
.B(n_134),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1669),
.B(n_135),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1772),
.A2(n_135),
.B(n_136),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1645),
.A2(n_137),
.B(n_138),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_SL g1922 ( 
.A(n_1608),
.B(n_1623),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1671),
.B(n_139),
.Y(n_1923)
);

A2O1A1Ixp33_ASAP7_75t_L g1924 ( 
.A1(n_1699),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_1924)
);

BUFx12f_ASAP7_75t_L g1925 ( 
.A(n_1655),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1734),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1658),
.A2(n_142),
.B(n_143),
.Y(n_1927)
);

OAI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1698),
.A2(n_144),
.B(n_145),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1659),
.A2(n_144),
.B(n_145),
.Y(n_1929)
);

AOI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1748),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.C(n_149),
.Y(n_1930)
);

AO32x1_ASAP7_75t_L g1931 ( 
.A1(n_1680),
.A2(n_152),
.A3(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1644),
.B(n_151),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1683),
.Y(n_1933)
);

O2A1O1Ixp5_ASAP7_75t_L g1934 ( 
.A1(n_1707),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1691),
.B(n_155),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1672),
.A2(n_155),
.B(n_156),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1685),
.A2(n_156),
.B(n_157),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1704),
.B(n_158),
.Y(n_1938)
);

AND2x6_ASAP7_75t_L g1939 ( 
.A(n_1783),
.B(n_333),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1710),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1660),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1636),
.B(n_158),
.Y(n_1942)
);

AOI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1673),
.A2(n_159),
.B(n_160),
.Y(n_1943)
);

AOI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1761),
.A2(n_161),
.B(n_162),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1623),
.B(n_161),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1775),
.A2(n_163),
.B(n_164),
.Y(n_1946)
);

A2O1A1Ixp33_ASAP7_75t_L g1947 ( 
.A1(n_1763),
.A2(n_165),
.B(n_163),
.C(n_164),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1657),
.B(n_165),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1644),
.B(n_167),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1668),
.Y(n_1950)
);

AOI221xp5_ASAP7_75t_L g1951 ( 
.A1(n_1743),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.C(n_170),
.Y(n_1951)
);

INVx3_ASAP7_75t_L g1952 ( 
.A(n_1660),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1692),
.A2(n_172),
.B1(n_168),
.B2(n_171),
.Y(n_1953)
);

OAI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1630),
.A2(n_174),
.B1(n_171),
.B2(n_173),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1717),
.B(n_173),
.Y(n_1955)
);

O2A1O1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1706),
.A2(n_1688),
.B(n_1638),
.C(n_1682),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1670),
.B(n_175),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1711),
.B(n_175),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1660),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1712),
.B(n_177),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1690),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_1961)
);

NAND3xp33_ASAP7_75t_L g1962 ( 
.A(n_1821),
.B(n_1715),
.C(n_1708),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1823),
.B(n_1716),
.Y(n_1963)
);

AOI21xp33_ASAP7_75t_L g1964 ( 
.A1(n_1792),
.A2(n_1754),
.B(n_1715),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1834),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1831),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1850),
.Y(n_1967)
);

NAND2x1p5_ASAP7_75t_L g1968 ( 
.A(n_1869),
.B(n_1608),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1834),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_L g1970 ( 
.A(n_1798),
.B(n_1679),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1895),
.B(n_1725),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1957),
.B(n_1679),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1790),
.B(n_1791),
.Y(n_1973)
);

NAND3xp33_ASAP7_75t_SL g1974 ( 
.A(n_1926),
.B(n_1649),
.C(n_1755),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1796),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1809),
.B(n_1679),
.Y(n_1976)
);

AOI21xp33_ASAP7_75t_L g1977 ( 
.A1(n_1799),
.A2(n_1780),
.B(n_1708),
.Y(n_1977)
);

AOI21xp33_ASAP7_75t_L g1978 ( 
.A1(n_1793),
.A2(n_1768),
.B(n_1762),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1906),
.B(n_1783),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1905),
.B(n_1739),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1868),
.Y(n_1981)
);

OAI21x1_ASAP7_75t_L g1982 ( 
.A1(n_1788),
.A2(n_1728),
.B(n_1696),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1787),
.A2(n_1602),
.B(n_1783),
.Y(n_1983)
);

NAND3xp33_ASAP7_75t_SL g1984 ( 
.A(n_1946),
.B(n_1833),
.C(n_1890),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1898),
.A2(n_1602),
.B(n_1741),
.Y(n_1985)
);

AOI21xp33_ASAP7_75t_L g1986 ( 
.A1(n_1956),
.A2(n_1701),
.B(n_1693),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1834),
.Y(n_1987)
);

AOI21x1_ASAP7_75t_L g1988 ( 
.A1(n_1789),
.A2(n_1662),
.B(n_1722),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1861),
.B(n_1739),
.Y(n_1989)
);

INVx3_ASAP7_75t_L g1990 ( 
.A(n_1925),
.Y(n_1990)
);

NAND2x1p5_ASAP7_75t_L g1991 ( 
.A(n_1857),
.B(n_1724),
.Y(n_1991)
);

OAI21x1_ASAP7_75t_SL g1992 ( 
.A1(n_1928),
.A2(n_1729),
.B(n_1739),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1897),
.A2(n_1739),
.B(n_178),
.Y(n_1993)
);

A2O1A1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1802),
.A2(n_181),
.B(n_179),
.C(n_180),
.Y(n_1994)
);

OAI21x1_ASAP7_75t_L g1995 ( 
.A1(n_1795),
.A2(n_335),
.B(n_334),
.Y(n_1995)
);

OAI21x1_ASAP7_75t_L g1996 ( 
.A1(n_1907),
.A2(n_338),
.B(n_337),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1819),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1922),
.B(n_339),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1913),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1879),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1917),
.Y(n_2001)
);

OAI21x1_ASAP7_75t_L g2002 ( 
.A1(n_1909),
.A2(n_342),
.B(n_340),
.Y(n_2002)
);

OAI21x1_ASAP7_75t_L g2003 ( 
.A1(n_1859),
.A2(n_349),
.B(n_343),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1801),
.A2(n_180),
.B(n_181),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1857),
.B(n_351),
.Y(n_2005)
);

OAI21xp33_ASAP7_75t_L g2006 ( 
.A1(n_1814),
.A2(n_182),
.B(n_183),
.Y(n_2006)
);

BUFx4f_ASAP7_75t_L g2007 ( 
.A(n_1817),
.Y(n_2007)
);

INVxp67_ASAP7_75t_SL g2008 ( 
.A(n_1940),
.Y(n_2008)
);

NAND2x1_ASAP7_75t_L g2009 ( 
.A(n_1817),
.B(n_182),
.Y(n_2009)
);

AOI21xp33_ASAP7_75t_L g2010 ( 
.A1(n_1910),
.A2(n_183),
.B(n_184),
.Y(n_2010)
);

BUFx5_ASAP7_75t_L g2011 ( 
.A(n_1939),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1933),
.B(n_184),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1896),
.Y(n_2013)
);

AOI21xp33_ASAP7_75t_L g2014 ( 
.A1(n_1881),
.A2(n_185),
.B(n_186),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1884),
.A2(n_185),
.B(n_186),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1860),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1812),
.B(n_187),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1902),
.B(n_188),
.Y(n_2018)
);

INVx5_ASAP7_75t_L g2019 ( 
.A(n_1939),
.Y(n_2019)
);

A2O1A1Ixp33_ASAP7_75t_L g2020 ( 
.A1(n_1852),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_2020)
);

OAI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1856),
.A2(n_190),
.B(n_191),
.Y(n_2021)
);

AO21x1_ASAP7_75t_L g2022 ( 
.A1(n_1876),
.A2(n_192),
.B(n_193),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1846),
.A2(n_193),
.B(n_194),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1950),
.B(n_194),
.Y(n_2024)
);

OAI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_1900),
.A2(n_1807),
.B(n_1848),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1888),
.A2(n_195),
.B(n_196),
.Y(n_2026)
);

O2A1O1Ixp5_ASAP7_75t_L g2027 ( 
.A1(n_1878),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_1880),
.Y(n_2028)
);

AOI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1873),
.A2(n_1931),
.B(n_1851),
.Y(n_2029)
);

BUFx2_ASAP7_75t_L g2030 ( 
.A(n_1875),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1903),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1857),
.B(n_352),
.Y(n_2032)
);

AO31x2_ASAP7_75t_L g2033 ( 
.A1(n_1827),
.A2(n_1937),
.A3(n_1921),
.B(n_1943),
.Y(n_2033)
);

OAI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_1832),
.A2(n_1916),
.B1(n_1829),
.B2(n_1947),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1830),
.A2(n_356),
.B(n_355),
.Y(n_2035)
);

OAI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1854),
.A2(n_197),
.B(n_198),
.Y(n_2036)
);

OAI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1904),
.A2(n_198),
.B(n_199),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1855),
.Y(n_2038)
);

OAI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_1844),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1813),
.B(n_1824),
.Y(n_2040)
);

AOI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_1931),
.A2(n_1836),
.B(n_1835),
.Y(n_2041)
);

BUFx4f_ASAP7_75t_L g2042 ( 
.A(n_1839),
.Y(n_2042)
);

AOI21xp33_ASAP7_75t_L g2043 ( 
.A1(n_1908),
.A2(n_201),
.B(n_202),
.Y(n_2043)
);

A2O1A1Ixp33_ASAP7_75t_L g2044 ( 
.A1(n_1810),
.A2(n_205),
.B(n_203),
.C(n_204),
.Y(n_2044)
);

OAI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_1837),
.A2(n_204),
.B(n_206),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1847),
.A2(n_207),
.B(n_208),
.Y(n_2046)
);

AO21x2_ASAP7_75t_L g2047 ( 
.A1(n_1841),
.A2(n_545),
.B(n_361),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1863),
.Y(n_2048)
);

AOI21x1_ASAP7_75t_L g2049 ( 
.A1(n_1822),
.A2(n_207),
.B(n_208),
.Y(n_2049)
);

INVxp67_ASAP7_75t_L g2050 ( 
.A(n_1800),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1865),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1804),
.B(n_1842),
.Y(n_2052)
);

OAI21x1_ASAP7_75t_L g2053 ( 
.A1(n_1845),
.A2(n_362),
.B(n_359),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1914),
.Y(n_2054)
);

AOI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_1887),
.A2(n_210),
.B(n_211),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1893),
.A2(n_210),
.B(n_211),
.Y(n_2056)
);

AOI21x1_ASAP7_75t_L g2057 ( 
.A1(n_1820),
.A2(n_212),
.B(n_214),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_1867),
.A2(n_212),
.B(n_215),
.Y(n_2058)
);

OAI21x1_ASAP7_75t_L g2059 ( 
.A1(n_1918),
.A2(n_364),
.B(n_363),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1849),
.B(n_216),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1891),
.A2(n_217),
.B(n_218),
.Y(n_2061)
);

OAI21xp33_ASAP7_75t_L g2062 ( 
.A1(n_1924),
.A2(n_218),
.B(n_219),
.Y(n_2062)
);

OAI21x1_ASAP7_75t_L g2063 ( 
.A1(n_1899),
.A2(n_367),
.B(n_365),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_1843),
.A2(n_219),
.B(n_220),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1853),
.B(n_220),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_L g2066 ( 
.A1(n_1934),
.A2(n_369),
.B(n_368),
.Y(n_2066)
);

A2O1A1Ixp33_ASAP7_75t_L g2067 ( 
.A1(n_1930),
.A2(n_223),
.B(n_221),
.C(n_222),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1864),
.B(n_221),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1948),
.B(n_222),
.Y(n_2069)
);

A2O1A1Ixp33_ASAP7_75t_L g2070 ( 
.A1(n_1889),
.A2(n_225),
.B(n_223),
.C(n_224),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1794),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1942),
.B(n_1870),
.Y(n_2072)
);

BUFx3_ASAP7_75t_L g2073 ( 
.A(n_1839),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1882),
.Y(n_2074)
);

OAI21x1_ASAP7_75t_L g2075 ( 
.A1(n_1927),
.A2(n_371),
.B(n_370),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_SL g2076 ( 
.A1(n_1885),
.A2(n_224),
.B(n_225),
.Y(n_2076)
);

OAI21x1_ASAP7_75t_L g2077 ( 
.A1(n_1929),
.A2(n_373),
.B(n_372),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1892),
.B(n_226),
.Y(n_2078)
);

NAND3xp33_ASAP7_75t_L g2079 ( 
.A(n_1951),
.B(n_226),
.C(n_227),
.Y(n_2079)
);

BUFx12f_ASAP7_75t_L g2080 ( 
.A(n_1965),
.Y(n_2080)
);

BUFx2_ASAP7_75t_SL g2081 ( 
.A(n_2019),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_1962),
.A2(n_1828),
.B1(n_1825),
.B2(n_1938),
.Y(n_2082)
);

BUFx4_ASAP7_75t_SL g2083 ( 
.A(n_2073),
.Y(n_2083)
);

INVx3_ASAP7_75t_SL g2084 ( 
.A(n_1965),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_1967),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1966),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2008),
.B(n_1919),
.Y(n_2087)
);

INVx3_ASAP7_75t_L g2088 ( 
.A(n_2040),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_2030),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_2042),
.Y(n_2090)
);

INVx4_ASAP7_75t_L g2091 ( 
.A(n_2019),
.Y(n_2091)
);

NAND2x1_ASAP7_75t_L g2092 ( 
.A(n_1989),
.B(n_1886),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_2019),
.B(n_2001),
.Y(n_2093)
);

CKINVDCx20_ASAP7_75t_R g2094 ( 
.A(n_2042),
.Y(n_2094)
);

BUFx3_ASAP7_75t_L g2095 ( 
.A(n_2028),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1976),
.B(n_1826),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1975),
.Y(n_2097)
);

BUFx3_ASAP7_75t_L g2098 ( 
.A(n_1965),
.Y(n_2098)
);

CKINVDCx20_ASAP7_75t_R g2099 ( 
.A(n_1972),
.Y(n_2099)
);

BUFx2_ASAP7_75t_SL g2100 ( 
.A(n_2011),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_2040),
.B(n_1874),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_1969),
.Y(n_2102)
);

INVx4_ASAP7_75t_L g2103 ( 
.A(n_2007),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1981),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1970),
.B(n_1912),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1997),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1969),
.Y(n_2107)
);

BUFx6f_ASAP7_75t_L g2108 ( 
.A(n_1969),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_SL g2109 ( 
.A(n_2011),
.B(n_1939),
.Y(n_2109)
);

AOI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_1984),
.A2(n_1911),
.B1(n_1883),
.B2(n_1953),
.Y(n_2110)
);

NAND2x1p5_ASAP7_75t_L g2111 ( 
.A(n_2007),
.B(n_1871),
.Y(n_2111)
);

BUFx2_ASAP7_75t_SL g2112 ( 
.A(n_2011),
.Y(n_2112)
);

CKINVDCx6p67_ASAP7_75t_R g2113 ( 
.A(n_1987),
.Y(n_2113)
);

AOI22xp33_ASAP7_75t_L g2114 ( 
.A1(n_2006),
.A2(n_2034),
.B1(n_2062),
.B2(n_2023),
.Y(n_2114)
);

NAND2x1p5_ASAP7_75t_L g2115 ( 
.A(n_2032),
.B(n_1987),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1999),
.Y(n_2116)
);

BUFx2_ASAP7_75t_R g2117 ( 
.A(n_2047),
.Y(n_2117)
);

BUFx12f_ASAP7_75t_L g2118 ( 
.A(n_1987),
.Y(n_2118)
);

INVx6_ASAP7_75t_L g2119 ( 
.A(n_2011),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1971),
.Y(n_2120)
);

BUFx8_ASAP7_75t_L g2121 ( 
.A(n_2068),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_1973),
.Y(n_2122)
);

INVx1_ASAP7_75t_SL g2123 ( 
.A(n_1980),
.Y(n_2123)
);

BUFx3_ASAP7_75t_L g2124 ( 
.A(n_1990),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2000),
.Y(n_2125)
);

BUFx10_ASAP7_75t_L g2126 ( 
.A(n_2032),
.Y(n_2126)
);

BUFx2_ASAP7_75t_L g2127 ( 
.A(n_2054),
.Y(n_2127)
);

INVx1_ASAP7_75t_SL g2128 ( 
.A(n_1963),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2013),
.Y(n_2129)
);

BUFx5_ASAP7_75t_L g2130 ( 
.A(n_2038),
.Y(n_2130)
);

BUFx4_ASAP7_75t_SL g2131 ( 
.A(n_2048),
.Y(n_2131)
);

BUFx4f_ASAP7_75t_L g2132 ( 
.A(n_1968),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2050),
.B(n_1816),
.Y(n_2133)
);

AOI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_2045),
.A2(n_1840),
.B1(n_1954),
.B2(n_1944),
.Y(n_2134)
);

OAI22xp33_ASAP7_75t_L g2135 ( 
.A1(n_2016),
.A2(n_1955),
.B1(n_1803),
.B2(n_1920),
.Y(n_2135)
);

BUFx2_ASAP7_75t_L g2136 ( 
.A(n_1990),
.Y(n_2136)
);

INVx4_ASAP7_75t_L g2137 ( 
.A(n_2011),
.Y(n_2137)
);

INVx8_ASAP7_75t_L g2138 ( 
.A(n_2009),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2031),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2051),
.B(n_1923),
.Y(n_2140)
);

BUFx3_ASAP7_75t_L g2141 ( 
.A(n_2071),
.Y(n_2141)
);

OR2x6_ASAP7_75t_L g2142 ( 
.A(n_1979),
.B(n_1886),
.Y(n_2142)
);

CKINVDCx20_ASAP7_75t_R g2143 ( 
.A(n_2024),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1982),
.Y(n_2144)
);

INVx2_ASAP7_75t_SL g2145 ( 
.A(n_2074),
.Y(n_2145)
);

CKINVDCx20_ASAP7_75t_R g2146 ( 
.A(n_2017),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2052),
.B(n_1935),
.Y(n_2147)
);

NAND2x1p5_ASAP7_75t_L g2148 ( 
.A(n_1988),
.B(n_1998),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2072),
.B(n_1858),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_1983),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2012),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1992),
.Y(n_2152)
);

BUFx8_ASAP7_75t_L g2153 ( 
.A(n_2018),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1986),
.Y(n_2154)
);

OAI21x1_ASAP7_75t_L g2155 ( 
.A1(n_2148),
.A2(n_2029),
.B(n_2041),
.Y(n_2155)
);

OAI22xp33_ASAP7_75t_SL g2156 ( 
.A1(n_2109),
.A2(n_2154),
.B1(n_2150),
.B2(n_2128),
.Y(n_2156)
);

INVxp67_ASAP7_75t_SL g2157 ( 
.A(n_2087),
.Y(n_2157)
);

NOR2x1_ASAP7_75t_R g2158 ( 
.A(n_2122),
.B(n_1797),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_2085),
.Y(n_2159)
);

OA21x2_ASAP7_75t_L g2160 ( 
.A1(n_2152),
.A2(n_1978),
.B(n_1964),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2097),
.Y(n_2161)
);

CKINVDCx9p33_ASAP7_75t_R g2162 ( 
.A(n_2089),
.Y(n_2162)
);

OAI21x1_ASAP7_75t_L g2163 ( 
.A1(n_2148),
.A2(n_1993),
.B(n_1985),
.Y(n_2163)
);

OAI21x1_ASAP7_75t_L g2164 ( 
.A1(n_2144),
.A2(n_2035),
.B(n_1996),
.Y(n_2164)
);

AO32x2_ASAP7_75t_L g2165 ( 
.A1(n_2145),
.A2(n_2039),
.A3(n_2022),
.B1(n_2076),
.B2(n_1977),
.Y(n_2165)
);

AOI22x1_ASAP7_75t_L g2166 ( 
.A1(n_2136),
.A2(n_2021),
.B1(n_2064),
.B2(n_2026),
.Y(n_2166)
);

AOI21xp5_ASAP7_75t_L g2167 ( 
.A1(n_2109),
.A2(n_2025),
.B(n_1994),
.Y(n_2167)
);

OA21x2_ASAP7_75t_L g2168 ( 
.A1(n_2150),
.A2(n_2003),
.B(n_1995),
.Y(n_2168)
);

BUFx2_ASAP7_75t_L g2169 ( 
.A(n_2127),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2106),
.Y(n_2170)
);

AO32x2_ASAP7_75t_L g2171 ( 
.A1(n_2137),
.A2(n_1974),
.A3(n_2065),
.B1(n_2060),
.B2(n_2010),
.Y(n_2171)
);

AO21x2_ASAP7_75t_L g2172 ( 
.A1(n_2087),
.A2(n_2014),
.B(n_2036),
.Y(n_2172)
);

BUFx2_ASAP7_75t_R g2173 ( 
.A(n_2090),
.Y(n_2173)
);

OAI21x1_ASAP7_75t_L g2174 ( 
.A1(n_2092),
.A2(n_2002),
.B(n_2004),
.Y(n_2174)
);

OAI21x1_ASAP7_75t_L g2175 ( 
.A1(n_2140),
.A2(n_2066),
.B(n_1991),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_2093),
.B(n_1839),
.Y(n_2176)
);

OAI21x1_ASAP7_75t_L g2177 ( 
.A1(n_2140),
.A2(n_2049),
.B(n_2053),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2116),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2139),
.Y(n_2179)
);

AO31x2_ASAP7_75t_L g2180 ( 
.A1(n_2137),
.A2(n_2070),
.A3(n_2044),
.B(n_2020),
.Y(n_2180)
);

OAI21x1_ASAP7_75t_L g2181 ( 
.A1(n_2115),
.A2(n_2057),
.B(n_2059),
.Y(n_2181)
);

OR2x6_ASAP7_75t_L g2182 ( 
.A(n_2081),
.B(n_2037),
.Y(n_2182)
);

AO21x2_ASAP7_75t_L g2183 ( 
.A1(n_2151),
.A2(n_1960),
.B(n_1958),
.Y(n_2183)
);

INVx1_ASAP7_75t_SL g2184 ( 
.A(n_2123),
.Y(n_2184)
);

INVx1_ASAP7_75t_SL g2185 ( 
.A(n_2123),
.Y(n_2185)
);

AO21x2_ASAP7_75t_L g2186 ( 
.A1(n_2147),
.A2(n_2078),
.B(n_2069),
.Y(n_2186)
);

NOR2xp67_ASAP7_75t_L g2187 ( 
.A(n_2091),
.B(n_1875),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2120),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2128),
.B(n_1805),
.Y(n_2189)
);

OAI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_2114),
.A2(n_2110),
.B1(n_2082),
.B2(n_2134),
.Y(n_2190)
);

OAI21xp5_ASAP7_75t_L g2191 ( 
.A1(n_2110),
.A2(n_2027),
.B(n_2067),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_2093),
.A2(n_2005),
.B(n_2055),
.Y(n_2192)
);

AOI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_2135),
.A2(n_2079),
.B1(n_2043),
.B2(n_2015),
.Y(n_2193)
);

OAI21x1_ASAP7_75t_L g2194 ( 
.A1(n_2111),
.A2(n_2061),
.B(n_2075),
.Y(n_2194)
);

OAI21x1_ASAP7_75t_L g2195 ( 
.A1(n_2111),
.A2(n_2077),
.B(n_2063),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_2088),
.B(n_2101),
.Y(n_2196)
);

INVx3_ASAP7_75t_L g2197 ( 
.A(n_2088),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_L g2198 ( 
.A1(n_2147),
.A2(n_2046),
.B(n_2056),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2101),
.B(n_1941),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2086),
.Y(n_2200)
);

AOI21x1_ASAP7_75t_L g2201 ( 
.A1(n_2149),
.A2(n_1838),
.B(n_1901),
.Y(n_2201)
);

CKINVDCx20_ASAP7_75t_R g2202 ( 
.A(n_2094),
.Y(n_2202)
);

AOI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_2190),
.A2(n_2141),
.B1(n_2146),
.B2(n_2143),
.Y(n_2203)
);

BUFx2_ASAP7_75t_R g2204 ( 
.A(n_2169),
.Y(n_2204)
);

BUFx2_ASAP7_75t_L g2205 ( 
.A(n_2162),
.Y(n_2205)
);

INVx4_ASAP7_75t_L g2206 ( 
.A(n_2182),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2157),
.B(n_2149),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2157),
.Y(n_2208)
);

AND2x4_ASAP7_75t_L g2209 ( 
.A(n_2196),
.B(n_2095),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2186),
.B(n_2130),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2161),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2159),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2170),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2178),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2186),
.Y(n_2215)
);

INVx3_ASAP7_75t_L g2216 ( 
.A(n_2197),
.Y(n_2216)
);

OA21x2_ASAP7_75t_L g2217 ( 
.A1(n_2155),
.A2(n_2125),
.B(n_2104),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2179),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_2196),
.Y(n_2219)
);

AOI22xp33_ASAP7_75t_L g2220 ( 
.A1(n_2190),
.A2(n_2096),
.B1(n_2130),
.B2(n_2133),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2188),
.Y(n_2221)
);

CKINVDCx20_ASAP7_75t_R g2222 ( 
.A(n_2202),
.Y(n_2222)
);

BUFx2_ASAP7_75t_R g2223 ( 
.A(n_2183),
.Y(n_2223)
);

OAI21x1_ASAP7_75t_L g2224 ( 
.A1(n_2164),
.A2(n_2105),
.B(n_2129),
.Y(n_2224)
);

INVx3_ASAP7_75t_L g2225 ( 
.A(n_2197),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_2176),
.Y(n_2226)
);

OAI21x1_ASAP7_75t_L g2227 ( 
.A1(n_2224),
.A2(n_2160),
.B(n_2163),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2217),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2217),
.Y(n_2229)
);

OR2x2_ASAP7_75t_L g2230 ( 
.A(n_2207),
.B(n_2159),
.Y(n_2230)
);

BUFx2_ASAP7_75t_L g2231 ( 
.A(n_2205),
.Y(n_2231)
);

INVx3_ASAP7_75t_L g2232 ( 
.A(n_2206),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2211),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_2206),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2207),
.B(n_2184),
.Y(n_2235)
);

BUFx2_ASAP7_75t_SL g2236 ( 
.A(n_2222),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2217),
.Y(n_2237)
);

CKINVDCx20_ASAP7_75t_R g2238 ( 
.A(n_2205),
.Y(n_2238)
);

INVx3_ASAP7_75t_L g2239 ( 
.A(n_2232),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_2228),
.Y(n_2240)
);

INVx2_ASAP7_75t_SL g2241 ( 
.A(n_2232),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2228),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2229),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2233),
.Y(n_2244)
);

INVx3_ASAP7_75t_L g2245 ( 
.A(n_2232),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2244),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2245),
.B(n_2231),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2245),
.B(n_2231),
.Y(n_2248)
);

AO31x2_ASAP7_75t_L g2249 ( 
.A1(n_2240),
.A2(n_2215),
.A3(n_2237),
.B(n_2229),
.Y(n_2249)
);

HB1xp67_ASAP7_75t_L g2250 ( 
.A(n_2241),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2240),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2242),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2242),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2239),
.B(n_2234),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2243),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2246),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2251),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2249),
.Y(n_2258)
);

AND2x4_ASAP7_75t_L g2259 ( 
.A(n_2247),
.B(n_2238),
.Y(n_2259)
);

HB1xp67_ASAP7_75t_L g2260 ( 
.A(n_2250),
.Y(n_2260)
);

OR2x2_ASAP7_75t_L g2261 ( 
.A(n_2250),
.B(n_2230),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2248),
.B(n_2241),
.Y(n_2262)
);

BUFx2_ASAP7_75t_L g2263 ( 
.A(n_2254),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2254),
.B(n_2234),
.Y(n_2264)
);

HB1xp67_ASAP7_75t_L g2265 ( 
.A(n_2252),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2253),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2255),
.B(n_2234),
.Y(n_2267)
);

BUFx3_ASAP7_75t_L g2268 ( 
.A(n_2259),
.Y(n_2268)
);

NAND4xp25_ASAP7_75t_L g2269 ( 
.A(n_2263),
.B(n_2239),
.C(n_2191),
.D(n_2193),
.Y(n_2269)
);

O2A1O1Ixp33_ASAP7_75t_L g2270 ( 
.A1(n_2260),
.A2(n_2191),
.B(n_2243),
.C(n_2193),
.Y(n_2270)
);

OAI21x1_ASAP7_75t_L g2271 ( 
.A1(n_2261),
.A2(n_2239),
.B(n_2235),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2259),
.Y(n_2272)
);

OAI211xp5_ASAP7_75t_L g2273 ( 
.A1(n_2256),
.A2(n_2166),
.B(n_2206),
.C(n_1877),
.Y(n_2273)
);

BUFx3_ASAP7_75t_L g2274 ( 
.A(n_2259),
.Y(n_2274)
);

INVx4_ASAP7_75t_L g2275 ( 
.A(n_2262),
.Y(n_2275)
);

INVx2_ASAP7_75t_SL g2276 ( 
.A(n_2262),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2273),
.A2(n_2258),
.B1(n_2266),
.B2(n_2257),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_2276),
.B(n_2261),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2268),
.Y(n_2279)
);

OAI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2270),
.A2(n_2265),
.B(n_2267),
.Y(n_2280)
);

INVxp67_ASAP7_75t_L g2281 ( 
.A(n_2278),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2279),
.B(n_2269),
.Y(n_2282)
);

INVx1_ASAP7_75t_SL g2283 ( 
.A(n_2280),
.Y(n_2283)
);

HB1xp67_ASAP7_75t_L g2284 ( 
.A(n_2277),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2282),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2283),
.B(n_2274),
.Y(n_2286)
);

INVx1_ASAP7_75t_SL g2287 ( 
.A(n_2284),
.Y(n_2287)
);

BUFx2_ASAP7_75t_L g2288 ( 
.A(n_2281),
.Y(n_2288)
);

A2O1A1Ixp33_ASAP7_75t_L g2289 ( 
.A1(n_2284),
.A2(n_2273),
.B(n_2269),
.C(n_2272),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2283),
.B(n_2275),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2288),
.Y(n_2291)
);

INVx2_ASAP7_75t_SL g2292 ( 
.A(n_2286),
.Y(n_2292)
);

OAI22xp33_ASAP7_75t_L g2293 ( 
.A1(n_2287),
.A2(n_2275),
.B1(n_2258),
.B2(n_2267),
.Y(n_2293)
);

NAND4xp25_ASAP7_75t_SL g2294 ( 
.A(n_2289),
.B(n_2264),
.C(n_2271),
.D(n_2236),
.Y(n_2294)
);

AOI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2285),
.A2(n_2236),
.B1(n_2264),
.B2(n_2215),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2290),
.B(n_2235),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_SL g2297 ( 
.A(n_2287),
.B(n_2204),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2288),
.Y(n_2298)
);

O2A1O1Ixp33_ASAP7_75t_L g2299 ( 
.A1(n_2289),
.A2(n_2203),
.B(n_2182),
.C(n_2210),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2288),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2297),
.B(n_2230),
.Y(n_2301)
);

INVx1_ASAP7_75t_SL g2302 ( 
.A(n_2292),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2291),
.B(n_2298),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2300),
.B(n_2209),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2296),
.Y(n_2305)
);

INVx1_ASAP7_75t_SL g2306 ( 
.A(n_2295),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2294),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2293),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_2299),
.B(n_2209),
.Y(n_2309)
);

INVx1_ASAP7_75t_SL g2310 ( 
.A(n_2297),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_2292),
.Y(n_2311)
);

NOR2x1_ASAP7_75t_SL g2312 ( 
.A(n_2292),
.B(n_2158),
.Y(n_2312)
);

INVx1_ASAP7_75t_SL g2313 ( 
.A(n_2292),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2311),
.B(n_2153),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2311),
.Y(n_2315)
);

INVx1_ASAP7_75t_SL g2316 ( 
.A(n_2302),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2302),
.B(n_2153),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2313),
.Y(n_2318)
);

NAND2x1p5_ASAP7_75t_L g2319 ( 
.A(n_2313),
.B(n_2310),
.Y(n_2319)
);

AND2x4_ASAP7_75t_L g2320 ( 
.A(n_2304),
.B(n_2209),
.Y(n_2320)
);

INVx2_ASAP7_75t_SL g2321 ( 
.A(n_2301),
.Y(n_2321)
);

OAI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2308),
.A2(n_2173),
.B1(n_2233),
.B2(n_2220),
.Y(n_2322)
);

O2A1O1Ixp33_ASAP7_75t_SL g2323 ( 
.A1(n_2303),
.A2(n_2212),
.B(n_2131),
.C(n_2083),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2305),
.B(n_2121),
.Y(n_2324)
);

AOI22xp5_ASAP7_75t_SL g2325 ( 
.A1(n_2307),
.A2(n_1915),
.B1(n_2124),
.B2(n_2121),
.Y(n_2325)
);

NAND2xp33_ASAP7_75t_L g2326 ( 
.A(n_2306),
.B(n_2138),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2309),
.A2(n_2173),
.B1(n_2208),
.B2(n_2189),
.Y(n_2327)
);

OAI31xp33_ASAP7_75t_L g2328 ( 
.A1(n_2309),
.A2(n_2237),
.A3(n_2156),
.B(n_2167),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2319),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2316),
.B(n_2312),
.Y(n_2330)
);

OAI32xp33_ASAP7_75t_L g2331 ( 
.A1(n_2317),
.A2(n_2208),
.A3(n_1811),
.B1(n_2189),
.B2(n_2103),
.Y(n_2331)
);

AOI21xp5_ASAP7_75t_L g2332 ( 
.A1(n_2314),
.A2(n_1945),
.B(n_2058),
.Y(n_2332)
);

OAI221xp5_ASAP7_75t_SL g2333 ( 
.A1(n_2321),
.A2(n_2182),
.B1(n_2167),
.B2(n_1961),
.C(n_1815),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2320),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2318),
.B(n_2249),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2315),
.B(n_2249),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2324),
.B(n_2249),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2325),
.Y(n_2338)
);

OAI21xp33_ASAP7_75t_SL g2339 ( 
.A1(n_2328),
.A2(n_2227),
.B(n_2225),
.Y(n_2339)
);

OAI21x1_ASAP7_75t_SL g2340 ( 
.A1(n_2327),
.A2(n_2201),
.B(n_2103),
.Y(n_2340)
);

OAI221xp5_ASAP7_75t_L g2341 ( 
.A1(n_2326),
.A2(n_2132),
.B1(n_1936),
.B2(n_1808),
.C(n_2221),
.Y(n_2341)
);

NAND2x1p5_ASAP7_75t_L g2342 ( 
.A(n_2323),
.B(n_2132),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2329),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2330),
.B(n_2322),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2334),
.B(n_2227),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2342),
.B(n_2219),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2338),
.B(n_2183),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2335),
.Y(n_2348)
);

OAI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2341),
.A2(n_2223),
.B1(n_2213),
.B2(n_2214),
.Y(n_2349)
);

AND2x4_ASAP7_75t_L g2350 ( 
.A(n_2337),
.B(n_2176),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2336),
.Y(n_2351)
);

NOR2x1p5_ASAP7_75t_L g2352 ( 
.A(n_2331),
.B(n_2216),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2339),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2340),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2332),
.B(n_2221),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2333),
.B(n_2099),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2329),
.B(n_2138),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2329),
.B(n_2172),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2329),
.B(n_2219),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2329),
.B(n_2226),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2329),
.B(n_2172),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2329),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2329),
.Y(n_2363)
);

OAI221xp5_ASAP7_75t_SL g2364 ( 
.A1(n_2339),
.A2(n_1862),
.B1(n_2192),
.B2(n_1949),
.C(n_2171),
.Y(n_2364)
);

OAI21xp33_ASAP7_75t_L g2365 ( 
.A1(n_2362),
.A2(n_2226),
.B(n_2225),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2363),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_SL g2367 ( 
.A(n_2343),
.B(n_1871),
.Y(n_2367)
);

NOR3x1_ASAP7_75t_L g2368 ( 
.A(n_2344),
.B(n_227),
.C(n_228),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2350),
.B(n_2224),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_L g2370 ( 
.A(n_2350),
.B(n_2138),
.Y(n_2370)
);

NAND4xp75_ASAP7_75t_L g2371 ( 
.A(n_2351),
.B(n_2160),
.C(n_230),
.D(n_228),
.Y(n_2371)
);

NOR3xp33_ASAP7_75t_L g2372 ( 
.A(n_2348),
.B(n_1932),
.C(n_229),
.Y(n_2372)
);

NOR3xp33_ASAP7_75t_L g2373 ( 
.A(n_2353),
.B(n_1932),
.C(n_229),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2359),
.B(n_2211),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2346),
.Y(n_2375)
);

NOR3xp33_ASAP7_75t_L g2376 ( 
.A(n_2354),
.B(n_230),
.C(n_231),
.Y(n_2376)
);

OAI211xp5_ASAP7_75t_SL g2377 ( 
.A1(n_2358),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_2377)
);

NAND4xp25_ASAP7_75t_L g2378 ( 
.A(n_2357),
.B(n_2192),
.C(n_234),
.D(n_232),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2355),
.Y(n_2379)
);

OAI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2345),
.A2(n_2177),
.B(n_2198),
.Y(n_2380)
);

NAND4xp25_ASAP7_75t_L g2381 ( 
.A(n_2360),
.B(n_235),
.C(n_233),
.D(n_234),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2356),
.B(n_2226),
.Y(n_2382)
);

AOI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_2361),
.A2(n_2214),
.B(n_2213),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2347),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2352),
.Y(n_2385)
);

BUFx2_ASAP7_75t_L g2386 ( 
.A(n_2349),
.Y(n_2386)
);

NOR3xp33_ASAP7_75t_L g2387 ( 
.A(n_2364),
.B(n_236),
.C(n_237),
.Y(n_2387)
);

AOI21xp33_ASAP7_75t_SL g2388 ( 
.A1(n_2353),
.A2(n_237),
.B(n_238),
.Y(n_2388)
);

OAI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2344),
.A2(n_2194),
.B(n_2174),
.Y(n_2389)
);

NAND4xp25_ASAP7_75t_L g2390 ( 
.A(n_2343),
.B(n_240),
.C(n_238),
.D(n_239),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2350),
.B(n_2218),
.Y(n_2391)
);

NAND5xp2_ASAP7_75t_L g2392 ( 
.A(n_2343),
.B(n_1786),
.C(n_242),
.D(n_243),
.E(n_244),
.Y(n_2392)
);

NOR3xp33_ASAP7_75t_L g2393 ( 
.A(n_2362),
.B(n_241),
.C(n_242),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_SL g2394 ( 
.A(n_2362),
.B(n_2080),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2350),
.B(n_2218),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2362),
.Y(n_2396)
);

NOR2x1_ASAP7_75t_SL g2397 ( 
.A(n_2362),
.B(n_2118),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2350),
.B(n_2217),
.Y(n_2398)
);

AOI22xp5_ASAP7_75t_L g2399 ( 
.A1(n_2353),
.A2(n_2185),
.B1(n_2184),
.B2(n_2130),
.Y(n_2399)
);

NAND3xp33_ASAP7_75t_L g2400 ( 
.A(n_2348),
.B(n_241),
.C(n_243),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2368),
.B(n_2185),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2366),
.Y(n_2402)
);

BUFx3_ASAP7_75t_L g2403 ( 
.A(n_2396),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2400),
.Y(n_2404)
);

NOR3xp33_ASAP7_75t_L g2405 ( 
.A(n_2384),
.B(n_244),
.C(n_245),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2392),
.B(n_245),
.Y(n_2406)
);

NOR2x1_ASAP7_75t_L g2407 ( 
.A(n_2375),
.B(n_246),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2397),
.B(n_2394),
.Y(n_2408)
);

AOI211xp5_ASAP7_75t_L g2409 ( 
.A1(n_2388),
.A2(n_1866),
.B(n_248),
.C(n_246),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2400),
.Y(n_2410)
);

AOI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2381),
.A2(n_247),
.B(n_248),
.Y(n_2411)
);

OAI21xp33_ASAP7_75t_L g2412 ( 
.A1(n_2378),
.A2(n_2367),
.B(n_2365),
.Y(n_2412)
);

AOI221x1_ASAP7_75t_L g2413 ( 
.A1(n_2385),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.C(n_252),
.Y(n_2413)
);

INVx2_ASAP7_75t_SL g2414 ( 
.A(n_2382),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2393),
.B(n_2168),
.Y(n_2415)
);

NAND3xp33_ASAP7_75t_L g2416 ( 
.A(n_2376),
.B(n_249),
.C(n_250),
.Y(n_2416)
);

AOI211xp5_ASAP7_75t_SL g2417 ( 
.A1(n_2379),
.A2(n_253),
.B(n_251),
.C(n_252),
.Y(n_2417)
);

OAI21xp33_ASAP7_75t_SL g2418 ( 
.A1(n_2399),
.A2(n_2162),
.B(n_2216),
.Y(n_2418)
);

AND2x2_ASAP7_75t_SL g2419 ( 
.A(n_2373),
.B(n_253),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_SL g2420 ( 
.A(n_2390),
.B(n_2386),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2377),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2372),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2370),
.B(n_254),
.Y(n_2423)
);

NOR2x1_ASAP7_75t_L g2424 ( 
.A(n_2374),
.B(n_254),
.Y(n_2424)
);

OAI21xp33_ASAP7_75t_L g2425 ( 
.A1(n_2387),
.A2(n_2225),
.B(n_2216),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2391),
.B(n_256),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2395),
.Y(n_2427)
);

NAND3xp33_ASAP7_75t_L g2428 ( 
.A(n_2389),
.B(n_256),
.C(n_258),
.Y(n_2428)
);

INVx2_ASAP7_75t_SL g2429 ( 
.A(n_2369),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2371),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2383),
.B(n_2168),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2407),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2424),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2403),
.Y(n_2434)
);

OAI21xp33_ASAP7_75t_SL g2435 ( 
.A1(n_2408),
.A2(n_2380),
.B(n_2398),
.Y(n_2435)
);

INVx2_ASAP7_75t_SL g2436 ( 
.A(n_2402),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2406),
.B(n_2199),
.Y(n_2437)
);

NOR3xp33_ASAP7_75t_L g2438 ( 
.A(n_2414),
.B(n_258),
.C(n_259),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2417),
.B(n_259),
.Y(n_2439)
);

OAI33xp33_ASAP7_75t_L g2440 ( 
.A1(n_2430),
.A2(n_260),
.A3(n_261),
.B1(n_263),
.B2(n_264),
.B3(n_265),
.Y(n_2440)
);

AOI221xp5_ASAP7_75t_L g2441 ( 
.A1(n_2412),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.C(n_264),
.Y(n_2441)
);

NAND4xp75_ASAP7_75t_L g2442 ( 
.A(n_2404),
.B(n_269),
.C(n_265),
.D(n_268),
.Y(n_2442)
);

OA22x2_ASAP7_75t_L g2443 ( 
.A1(n_2413),
.A2(n_2084),
.B1(n_2175),
.B2(n_2181),
.Y(n_2443)
);

AOI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_2427),
.A2(n_1939),
.B1(n_2130),
.B2(n_2113),
.Y(n_2444)
);

NAND3xp33_ASAP7_75t_L g2445 ( 
.A(n_2420),
.B(n_2410),
.C(n_2405),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2421),
.Y(n_2446)
);

OAI322xp33_ASAP7_75t_L g2447 ( 
.A1(n_2429),
.A2(n_269),
.A3(n_270),
.B1(n_271),
.B2(n_272),
.C1(n_273),
.C2(n_274),
.Y(n_2447)
);

OAI22xp5_ASAP7_75t_L g2448 ( 
.A1(n_2428),
.A2(n_2117),
.B1(n_2142),
.B2(n_2098),
.Y(n_2448)
);

NOR3x1_ASAP7_75t_L g2449 ( 
.A(n_2416),
.B(n_2422),
.C(n_2401),
.Y(n_2449)
);

NOR2xp33_ASAP7_75t_R g2450 ( 
.A(n_2426),
.B(n_270),
.Y(n_2450)
);

AOI221xp5_ASAP7_75t_L g2451 ( 
.A1(n_2411),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.C(n_277),
.Y(n_2451)
);

NAND4xp75_ASAP7_75t_L g2452 ( 
.A(n_2419),
.B(n_277),
.C(n_275),
.D(n_276),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2409),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2423),
.Y(n_2454)
);

OAI21xp33_ASAP7_75t_L g2455 ( 
.A1(n_2425),
.A2(n_2102),
.B(n_2117),
.Y(n_2455)
);

OAI211xp5_ASAP7_75t_SL g2456 ( 
.A1(n_2418),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_2456)
);

OAI21xp33_ASAP7_75t_SL g2457 ( 
.A1(n_2431),
.A2(n_2195),
.B(n_279),
.Y(n_2457)
);

AOI21xp33_ASAP7_75t_L g2458 ( 
.A1(n_2415),
.A2(n_280),
.B(n_281),
.Y(n_2458)
);

AOI22xp5_ASAP7_75t_L g2459 ( 
.A1(n_2418),
.A2(n_2130),
.B1(n_2142),
.B2(n_2108),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_2403),
.B(n_2107),
.Y(n_2460)
);

NAND2xp33_ASAP7_75t_L g2461 ( 
.A(n_2408),
.B(n_281),
.Y(n_2461)
);

OAI21xp5_ASAP7_75t_SL g2462 ( 
.A1(n_2408),
.A2(n_282),
.B(n_283),
.Y(n_2462)
);

AOI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_2402),
.A2(n_2142),
.B1(n_2108),
.B2(n_2107),
.Y(n_2463)
);

AOI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_2414),
.A2(n_282),
.B(n_284),
.Y(n_2464)
);

NAND4xp25_ASAP7_75t_SL g2465 ( 
.A(n_2408),
.B(n_284),
.C(n_285),
.D(n_286),
.Y(n_2465)
);

INVx1_ASAP7_75t_SL g2466 ( 
.A(n_2403),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_2403),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2407),
.Y(n_2468)
);

AOI211xp5_ASAP7_75t_L g2469 ( 
.A1(n_2402),
.A2(n_286),
.B(n_287),
.C(n_290),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2407),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2407),
.Y(n_2471)
);

AOI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2414),
.A2(n_287),
.B(n_290),
.Y(n_2472)
);

OAI22xp33_ASAP7_75t_SL g2473 ( 
.A1(n_2420),
.A2(n_2119),
.B1(n_2171),
.B2(n_2165),
.Y(n_2473)
);

AOI22xp5_ASAP7_75t_L g2474 ( 
.A1(n_2436),
.A2(n_2108),
.B1(n_2107),
.B2(n_2187),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2467),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2432),
.Y(n_2476)
);

AOI22xp5_ASAP7_75t_L g2477 ( 
.A1(n_2466),
.A2(n_2119),
.B1(n_2126),
.B2(n_2112),
.Y(n_2477)
);

OAI21xp33_ASAP7_75t_SL g2478 ( 
.A1(n_2434),
.A2(n_291),
.B(n_292),
.Y(n_2478)
);

OAI22xp5_ASAP7_75t_L g2479 ( 
.A1(n_2459),
.A2(n_2091),
.B1(n_2100),
.B2(n_2165),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2468),
.Y(n_2480)
);

OAI22xp5_ASAP7_75t_SL g2481 ( 
.A1(n_2439),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_2481)
);

AOI22xp5_ASAP7_75t_L g2482 ( 
.A1(n_2435),
.A2(n_2126),
.B1(n_2165),
.B2(n_2171),
.Y(n_2482)
);

AO22x2_ASAP7_75t_L g2483 ( 
.A1(n_2470),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_2483)
);

AOI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_2446),
.A2(n_2165),
.B1(n_2171),
.B2(n_1959),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2471),
.Y(n_2485)
);

AO22x2_ASAP7_75t_L g2486 ( 
.A1(n_2433),
.A2(n_2452),
.B1(n_2445),
.B2(n_2454),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2461),
.Y(n_2487)
);

AOI22xp5_ASAP7_75t_L g2488 ( 
.A1(n_2437),
.A2(n_2438),
.B1(n_2457),
.B2(n_2455),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2442),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2460),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2462),
.Y(n_2491)
);

NOR4xp25_ASAP7_75t_L g2492 ( 
.A(n_2456),
.B(n_297),
.C(n_298),
.D(n_299),
.Y(n_2492)
);

NOR2x1_ASAP7_75t_L g2493 ( 
.A(n_2465),
.B(n_298),
.Y(n_2493)
);

AOI22xp5_ASAP7_75t_L g2494 ( 
.A1(n_2453),
.A2(n_1959),
.B1(n_1952),
.B2(n_1941),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2450),
.Y(n_2495)
);

HB1xp67_ASAP7_75t_L g2496 ( 
.A(n_2449),
.Y(n_2496)
);

AOI22xp5_ASAP7_75t_L g2497 ( 
.A1(n_2451),
.A2(n_1952),
.B1(n_1818),
.B2(n_2200),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2443),
.Y(n_2498)
);

AOI22xp5_ASAP7_75t_L g2499 ( 
.A1(n_2440),
.A2(n_1818),
.B1(n_301),
.B2(n_302),
.Y(n_2499)
);

INVxp67_ASAP7_75t_SL g2500 ( 
.A(n_2469),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2464),
.B(n_300),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2447),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_L g2503 ( 
.A(n_2458),
.B(n_300),
.Y(n_2503)
);

NOR2x1_ASAP7_75t_L g2504 ( 
.A(n_2472),
.B(n_302),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2441),
.B(n_303),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2448),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2463),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2444),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2473),
.Y(n_2509)
);

A2O1A1Ixp33_ASAP7_75t_SL g2510 ( 
.A1(n_2476),
.A2(n_303),
.B(n_304),
.C(n_306),
.Y(n_2510)
);

OAI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_2496),
.A2(n_1806),
.B(n_304),
.Y(n_2511)
);

OR2x2_ASAP7_75t_L g2512 ( 
.A(n_2492),
.B(n_306),
.Y(n_2512)
);

AOI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2480),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2475),
.B(n_307),
.Y(n_2514)
);

AOI221xp5_ASAP7_75t_L g2515 ( 
.A1(n_2485),
.A2(n_2509),
.B1(n_2498),
.B2(n_2486),
.C(n_2502),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2495),
.B(n_308),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2487),
.B(n_310),
.Y(n_2517)
);

NAND3xp33_ASAP7_75t_L g2518 ( 
.A(n_2489),
.B(n_310),
.C(n_1818),
.Y(n_2518)
);

BUFx2_ASAP7_75t_L g2519 ( 
.A(n_2478),
.Y(n_2519)
);

NOR3xp33_ASAP7_75t_L g2520 ( 
.A(n_2490),
.B(n_375),
.C(n_376),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2483),
.Y(n_2521)
);

NOR3xp33_ASAP7_75t_L g2522 ( 
.A(n_2481),
.B(n_378),
.C(n_382),
.Y(n_2522)
);

NAND3xp33_ASAP7_75t_L g2523 ( 
.A(n_2491),
.B(n_383),
.C(n_385),
.Y(n_2523)
);

AOI211x1_ASAP7_75t_SL g2524 ( 
.A1(n_2505),
.A2(n_387),
.B(n_389),
.C(n_390),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2486),
.B(n_2504),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2483),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2493),
.B(n_391),
.Y(n_2527)
);

NOR3xp33_ASAP7_75t_L g2528 ( 
.A(n_2500),
.B(n_392),
.C(n_393),
.Y(n_2528)
);

AOI21xp33_ASAP7_75t_L g2529 ( 
.A1(n_2503),
.A2(n_394),
.B(n_395),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2501),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_L g2531 ( 
.A(n_2488),
.B(n_396),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_2506),
.B(n_399),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2499),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_SL g2534 ( 
.A(n_2507),
.B(n_1872),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2474),
.B(n_2180),
.Y(n_2535)
);

NOR2x1_ASAP7_75t_L g2536 ( 
.A(n_2508),
.B(n_400),
.Y(n_2536)
);

NOR3xp33_ASAP7_75t_L g2537 ( 
.A(n_2494),
.B(n_401),
.C(n_402),
.Y(n_2537)
);

AOI21xp5_ASAP7_75t_L g2538 ( 
.A1(n_2479),
.A2(n_404),
.B(n_405),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_2497),
.B(n_1872),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2477),
.B(n_408),
.Y(n_2540)
);

AOI21xp5_ASAP7_75t_L g2541 ( 
.A1(n_2482),
.A2(n_411),
.B(n_412),
.Y(n_2541)
);

HB1xp67_ASAP7_75t_L g2542 ( 
.A(n_2484),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2496),
.Y(n_2543)
);

NOR2x1_ASAP7_75t_L g2544 ( 
.A(n_2525),
.B(n_2543),
.Y(n_2544)
);

NOR2x1_ASAP7_75t_L g2545 ( 
.A(n_2521),
.B(n_2526),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2519),
.B(n_2180),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_2512),
.B(n_2180),
.Y(n_2547)
);

NOR2x1_ASAP7_75t_L g2548 ( 
.A(n_2530),
.B(n_413),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_2515),
.B(n_414),
.Y(n_2549)
);

NAND4xp25_ASAP7_75t_L g2550 ( 
.A(n_2524),
.B(n_416),
.C(n_419),
.D(n_420),
.Y(n_2550)
);

AOI21xp33_ASAP7_75t_SL g2551 ( 
.A1(n_2527),
.A2(n_423),
.B(n_427),
.Y(n_2551)
);

AND4x1_ASAP7_75t_L g2552 ( 
.A(n_2531),
.B(n_429),
.C(n_430),
.D(n_431),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2536),
.B(n_433),
.Y(n_2553)
);

AND2x2_ASAP7_75t_L g2554 ( 
.A(n_2532),
.B(n_2033),
.Y(n_2554)
);

INVx1_ASAP7_75t_SL g2555 ( 
.A(n_2517),
.Y(n_2555)
);

NAND4xp25_ASAP7_75t_L g2556 ( 
.A(n_2510),
.B(n_434),
.C(n_435),
.D(n_436),
.Y(n_2556)
);

NAND4xp75_ASAP7_75t_L g2557 ( 
.A(n_2533),
.B(n_437),
.C(n_438),
.D(n_439),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_2513),
.B(n_1872),
.Y(n_2558)
);

NAND4xp25_ASAP7_75t_L g2559 ( 
.A(n_2522),
.B(n_441),
.C(n_444),
.D(n_447),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2542),
.B(n_449),
.Y(n_2560)
);

XOR2x2_ASAP7_75t_L g2561 ( 
.A(n_2518),
.B(n_450),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2514),
.Y(n_2562)
);

NAND3x1_ASAP7_75t_L g2563 ( 
.A(n_2516),
.B(n_451),
.C(n_452),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2541),
.B(n_454),
.Y(n_2564)
);

INVx1_ASAP7_75t_SL g2565 ( 
.A(n_2553),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2544),
.Y(n_2566)
);

NOR2x1p5_ASAP7_75t_L g2567 ( 
.A(n_2556),
.B(n_2523),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2548),
.Y(n_2568)
);

NAND3xp33_ASAP7_75t_L g2569 ( 
.A(n_2545),
.B(n_2529),
.C(n_2528),
.Y(n_2569)
);

OR2x2_ASAP7_75t_L g2570 ( 
.A(n_2555),
.B(n_2534),
.Y(n_2570)
);

NOR3x1_ASAP7_75t_L g2571 ( 
.A(n_2560),
.B(n_2540),
.C(n_2511),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2562),
.B(n_2538),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2563),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2561),
.Y(n_2574)
);

AOI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_2549),
.A2(n_2537),
.B1(n_2520),
.B2(n_2535),
.Y(n_2575)
);

NOR3xp33_ASAP7_75t_L g2576 ( 
.A(n_2551),
.B(n_2539),
.C(n_456),
.Y(n_2576)
);

NOR3xp33_ASAP7_75t_L g2577 ( 
.A(n_2564),
.B(n_455),
.C(n_457),
.Y(n_2577)
);

AOI221xp5_ASAP7_75t_L g2578 ( 
.A1(n_2559),
.A2(n_458),
.B1(n_462),
.B2(n_464),
.C(n_468),
.Y(n_2578)
);

BUFx2_ASAP7_75t_L g2579 ( 
.A(n_2546),
.Y(n_2579)
);

XOR2x1_ASAP7_75t_L g2580 ( 
.A(n_2547),
.B(n_469),
.Y(n_2580)
);

NAND4xp75_ASAP7_75t_L g2581 ( 
.A(n_2566),
.B(n_2558),
.C(n_2554),
.D(n_2552),
.Y(n_2581)
);

NOR3xp33_ASAP7_75t_L g2582 ( 
.A(n_2579),
.B(n_2550),
.C(n_2557),
.Y(n_2582)
);

NOR2x1_ASAP7_75t_L g2583 ( 
.A(n_2569),
.B(n_470),
.Y(n_2583)
);

NOR3xp33_ASAP7_75t_SL g2584 ( 
.A(n_2574),
.B(n_472),
.C(n_473),
.Y(n_2584)
);

INVx1_ASAP7_75t_SL g2585 ( 
.A(n_2580),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2568),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2573),
.Y(n_2587)
);

NAND3xp33_ASAP7_75t_L g2588 ( 
.A(n_2570),
.B(n_475),
.C(n_476),
.Y(n_2588)
);

NOR3xp33_ASAP7_75t_L g2589 ( 
.A(n_2565),
.B(n_477),
.C(n_478),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2567),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2585),
.B(n_2571),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2590),
.Y(n_2592)
);

XOR2xp5_ASAP7_75t_L g2593 ( 
.A(n_2586),
.B(n_2572),
.Y(n_2593)
);

OAI22x1_ASAP7_75t_SL g2594 ( 
.A1(n_2587),
.A2(n_2575),
.B1(n_2576),
.B2(n_2577),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2581),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_SL g2596 ( 
.A(n_2592),
.B(n_2582),
.Y(n_2596)
);

OAI22x1_ASAP7_75t_L g2597 ( 
.A1(n_2593),
.A2(n_2583),
.B1(n_2588),
.B2(n_2584),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2591),
.Y(n_2598)
);

NOR2xp33_ASAP7_75t_L g2599 ( 
.A(n_2595),
.B(n_2589),
.Y(n_2599)
);

BUFx4f_ASAP7_75t_L g2600 ( 
.A(n_2594),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2600),
.Y(n_2601)
);

XOR2x1_ASAP7_75t_L g2602 ( 
.A(n_2598),
.B(n_2596),
.Y(n_2602)
);

HB1xp67_ASAP7_75t_L g2603 ( 
.A(n_2597),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2602),
.Y(n_2604)
);

XNOR2xp5_ASAP7_75t_L g2605 ( 
.A(n_2601),
.B(n_2599),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2603),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2606),
.B(n_2604),
.Y(n_2607)
);

OR2x2_ASAP7_75t_L g2608 ( 
.A(n_2605),
.B(n_2578),
.Y(n_2608)
);

OAI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2606),
.A2(n_1894),
.B1(n_482),
.B2(n_489),
.Y(n_2609)
);

OAI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2607),
.A2(n_479),
.B1(n_490),
.B2(n_495),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2610),
.Y(n_2611)
);

AOI221xp5_ASAP7_75t_L g2612 ( 
.A1(n_2611),
.A2(n_2608),
.B1(n_2609),
.B2(n_499),
.C(n_500),
.Y(n_2612)
);

AOI22xp5_ASAP7_75t_L g2613 ( 
.A1(n_2612),
.A2(n_496),
.B1(n_497),
.B2(n_501),
.Y(n_2613)
);

AOI21xp5_ASAP7_75t_L g2614 ( 
.A1(n_2613),
.A2(n_503),
.B(n_505),
.Y(n_2614)
);

XNOR2xp5_ASAP7_75t_L g2615 ( 
.A(n_2614),
.B(n_506),
.Y(n_2615)
);

AOI221xp5_ASAP7_75t_L g2616 ( 
.A1(n_2615),
.A2(n_507),
.B1(n_508),
.B2(n_509),
.C(n_511),
.Y(n_2616)
);

AOI22xp5_ASAP7_75t_L g2617 ( 
.A1(n_2616),
.A2(n_1894),
.B1(n_513),
.B2(n_514),
.Y(n_2617)
);

AOI211xp5_ASAP7_75t_L g2618 ( 
.A1(n_2617),
.A2(n_512),
.B(n_515),
.C(n_516),
.Y(n_2618)
);


endmodule