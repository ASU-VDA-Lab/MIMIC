module fake_jpeg_25497_n_167 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_10),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_33),
.B(n_35),
.Y(n_48)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_6),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_7),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_16),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_20),
.B1(n_15),
.B2(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_59),
.B1(n_24),
.B2(n_18),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_20),
.B1(n_15),
.B2(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_31),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_69),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_31),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_76),
.B1(n_87),
.B2(n_19),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_24),
.B1(n_18),
.B2(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_84),
.Y(n_100)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_61),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_23),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_90),
.Y(n_101)
);

AOI22x1_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_61),
.B1(n_63),
.B2(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_29),
.B1(n_25),
.B2(n_23),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_3),
.B(n_4),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_4),
.B(n_5),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_31),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_21),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_4),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_95),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_54),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_98),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_102),
.B1(n_81),
.B2(n_75),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_52),
.B1(n_57),
.B2(n_19),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_72),
.B1(n_84),
.B2(n_75),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_52),
.C(n_19),
.Y(n_98)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_17),
.A3(n_38),
.B1(n_9),
.B2(n_8),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_106),
.B(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_77),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_17),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_113),
.B(n_115),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_70),
.B1(n_89),
.B2(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_105),
.B1(n_95),
.B2(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_108),
.B(n_81),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_89),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_79),
.B1(n_74),
.B2(n_118),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_98),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_125),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_108),
.B(n_106),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_136),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_112),
.C(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_137),
.B(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_113),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_143),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_123),
.C(n_114),
.Y(n_140)
);

OA21x2_ASAP7_75t_SL g151 ( 
.A1(n_140),
.A2(n_141),
.B(n_132),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_111),
.B(n_109),
.C(n_79),
.D(n_17),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_111),
.C(n_109),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_128),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_128),
.B1(n_129),
.B2(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_149),
.B(n_142),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_157),
.B(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_117),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_140),
.B(n_144),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_152),
.C(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_161),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_126),
.B1(n_130),
.B2(n_8),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_160),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_162),
.A2(n_13),
.B(n_83),
.C(n_163),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_83),
.C(n_13),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_83),
.Y(n_167)
);


endmodule