module fake_jpeg_17468_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_0),
.B(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_33),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NAND2x1_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_19),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_16),
.B1(n_30),
.B2(n_24),
.Y(n_70)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_60),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_16),
.B1(n_29),
.B2(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_16),
.B1(n_29),
.B2(n_30),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_67),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_29),
.B1(n_38),
.B2(n_16),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_30),
.B1(n_18),
.B2(n_17),
.Y(n_90)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_22),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_69),
.B(n_87),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_28),
.B1(n_33),
.B2(n_32),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_42),
.B1(n_20),
.B2(n_19),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_25),
.B1(n_24),
.B2(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_76),
.B1(n_82),
.B2(n_86),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_28),
.B1(n_17),
.B2(n_32),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

OAI22x1_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_19),
.B1(n_27),
.B2(n_26),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_89),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_45),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_25),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_19),
.B(n_49),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_19),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_31),
.B1(n_18),
.B2(n_27),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_46),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_48),
.C(n_44),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_106),
.C(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_44),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_101),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_96),
.B(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_109),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_48),
.C(n_20),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_66),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_51),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_114),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_48),
.C(n_20),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_51),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_19),
.B(n_80),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_53),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_80),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_82),
.B1(n_69),
.B2(n_90),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_122),
.A2(n_96),
.B1(n_103),
.B2(n_115),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_139),
.Y(n_175)
);

OAI22x1_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_82),
.B1(n_74),
.B2(n_92),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_142),
.B1(n_113),
.B2(n_112),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_74),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_128),
.A2(n_132),
.B(n_147),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_72),
.B(n_74),
.Y(n_132)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_93),
.A2(n_47),
.B1(n_88),
.B2(n_74),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_97),
.B1(n_104),
.B2(n_106),
.Y(n_152)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_47),
.B1(n_91),
.B2(n_88),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_47),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_57),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_88),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_127),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_150),
.A2(n_177),
.B1(n_50),
.B2(n_144),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_117),
.A3(n_97),
.B1(n_95),
.B2(n_109),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_151),
.B(n_153),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_156),
.B1(n_158),
.B2(n_164),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_106),
.C(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_101),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_178),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_104),
.B1(n_99),
.B2(n_98),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_131),
.B1(n_122),
.B2(n_121),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_125),
.B1(n_123),
.B2(n_137),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_117),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_98),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_129),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_114),
.B1(n_111),
.B2(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_105),
.B(n_100),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_172),
.B(n_31),
.Y(n_196)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_171),
.B(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_170),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_48),
.B(n_57),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_123),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_13),
.B(n_11),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_176),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_64),
.B1(n_119),
.B2(n_83),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_121),
.B1(n_134),
.B2(n_146),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_186),
.B1(n_192),
.B2(n_162),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_161),
.A2(n_131),
.B(n_126),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_182),
.A2(n_187),
.B(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_203),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_145),
.B1(n_129),
.B2(n_134),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_138),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_198),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_151),
.A2(n_119),
.B1(n_53),
.B2(n_54),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_144),
.B(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_200),
.B1(n_164),
.B2(n_166),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_31),
.Y(n_197)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_31),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_26),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_162),
.C(n_171),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_170),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_149),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_167),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_176),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_159),
.B1(n_202),
.B2(n_194),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_196),
.B1(n_191),
.B2(n_190),
.Y(n_235)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_218),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_185),
.B(n_178),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_179),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_155),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_214),
.C(n_216),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_157),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_156),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_224),
.C(n_186),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_163),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_225),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_165),
.C(n_149),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_197),
.B(n_173),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_189),
.A2(n_163),
.B1(n_144),
.B2(n_3),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_8),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_187),
.A2(n_26),
.B(n_2),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_181),
.B(n_179),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_180),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_237),
.C(n_241),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_235),
.B(n_222),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_204),
.B1(n_183),
.B2(n_182),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_204),
.C(n_191),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_193),
.C(n_199),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_242),
.B(n_229),
.Y(n_255)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_247),
.C(n_249),
.Y(n_263)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_20),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_248),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_20),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_1),
.C(n_3),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_208),
.C(n_207),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_217),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_4),
.B(n_5),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_217),
.B(n_215),
.Y(n_253)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_261),
.B(n_262),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_209),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_221),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_264),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_232),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_265),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_206),
.B(n_207),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_254),
.A2(n_262),
.B1(n_258),
.B2(n_259),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_279),
.B1(n_265),
.B2(n_258),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_243),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_275),
.Y(n_288)
);

OAI221xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_244),
.B1(n_242),
.B2(n_206),
.C(n_250),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_241),
.Y(n_275)
);

OAI221xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_237),
.B1(n_235),
.B2(n_233),
.C(n_231),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_231),
.C(n_245),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_280),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_247),
.C(n_249),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_290),
.Y(n_298)
);

AOI21x1_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_264),
.B(n_267),
.Y(n_284)
);

AOI322xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_286),
.A3(n_290),
.B1(n_282),
.B2(n_285),
.C1(n_14),
.C2(n_10),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_259),
.B1(n_263),
.B2(n_212),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_277),
.A2(n_263),
.B1(n_5),
.B2(n_6),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_287),
.B(n_291),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_9),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_9),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_281),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_15),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_291),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_274),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_297),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_297),
.Y(n_304)
);

AOI21x1_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_272),
.B(n_280),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_299),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_287),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_12),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_303),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_15),
.C(n_296),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_304),
.A2(n_301),
.B(n_302),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_300),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_307),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_308),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_302),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_306),
.Y(n_311)
);


endmodule