module real_jpeg_22921_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_0),
.B(n_37),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_0),
.B(n_132),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_0),
.B(n_32),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_0),
.B(n_45),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_0),
.B(n_43),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_0),
.B(n_26),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_0),
.B(n_51),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_0),
.B(n_75),
.Y(n_295)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_2),
.B(n_43),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_2),
.B(n_26),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_3),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_3),
.B(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_3),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_3),
.B(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_3),
.B(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_3),
.B(n_17),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_3),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_3),
.B(n_32),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_4),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_4),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_4),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_4),
.B(n_37),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_4),
.B(n_32),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_4),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_7),
.B(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_7),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_7),
.B(n_37),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_7),
.B(n_32),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx8_ASAP7_75t_SL g52 ( 
.A(n_9),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_10),
.B(n_32),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_10),
.B(n_37),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_10),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_10),
.B(n_45),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_10),
.B(n_43),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_10),
.B(n_26),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_10),
.B(n_51),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_10),
.B(n_55),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_12),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_12),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_12),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_12),
.B(n_37),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_12),
.B(n_32),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_12),
.B(n_45),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_12),
.B(n_43),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_12),
.B(n_26),
.Y(n_308)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_14),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_14),
.B(n_37),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_14),
.B(n_32),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_14),
.B(n_45),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_14),
.B(n_43),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_14),
.B(n_26),
.Y(n_264)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_14),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_14),
.B(n_75),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_15),
.B(n_26),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_15),
.B(n_51),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_15),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_15),
.B(n_37),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_16),
.B(n_45),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_16),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_16),
.B(n_37),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_16),
.B(n_43),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_16),
.B(n_26),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_16),
.B(n_51),
.Y(n_212)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_17),
.Y(n_133)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_17),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_117),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_88),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_21),
.A2(n_22),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.C(n_64),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_23),
.B(n_358),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.C(n_47),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_24),
.B(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_29),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_25),
.B(n_31),
.C(n_34),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_39),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_30),
.A2(n_31),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_31),
.B(n_80),
.C(n_83),
.Y(n_95)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_32),
.Y(n_150)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_67),
.C(n_70),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_34),
.A2(n_39),
.B1(n_67),
.B2(n_68),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_35),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_35),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_36),
.B(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_40),
.B(n_47),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.C(n_44),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_41),
.B(n_42),
.CI(n_44),
.CON(n_322),
.SN(n_322)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_43),
.Y(n_289)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g368 ( 
.A(n_47),
.Y(n_368)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.CI(n_50),
.CON(n_47),
.SN(n_47)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_49),
.C(n_50),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_53),
.A2(n_64),
.B1(n_65),
.B2(n_359),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_53),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_60),
.C(n_63),
.Y(n_93)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_58),
.B(n_149),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_62),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_73),
.C(n_76),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_66),
.B(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_67),
.A2(n_68),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_67),
.B(n_299),
.C(n_300),
.Y(n_321)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_69),
.B(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_70),
.B(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_72),
.B(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_332),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_76),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_76),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_76),
.B(n_328),
.C(n_331),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_77),
.B(n_88),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_86),
.C(n_87),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_78),
.A2(n_79),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_81),
.B(n_84),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_85),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_100),
.C(n_101),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_84),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_86),
.B(n_87),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_95),
.C(n_96),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_106),
.Y(n_105)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.CI(n_93),
.CON(n_90),
.SN(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_100),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_115),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_360),
.C(n_361),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_348),
.C(n_349),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_336),
.C(n_337),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_312),
.C(n_313),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_280),
.C(n_281),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_246),
.C(n_247),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_216),
.C(n_217),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_195),
.C(n_196),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_177),
.C(n_178),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_155),
.C(n_156),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_141),
.C(n_146),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_137),
.B2(n_138),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_139),
.C(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_131),
.Y(n_136)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_133),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_136),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.C(n_151),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_168),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_161),
.C(n_168),
.Y(n_177)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_162),
.Y(n_167)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_165),
.B(n_167),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_176),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_175),
.C(n_176),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_186),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_181),
.C(n_186),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_184),
.C(n_185),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_189),
.C(n_190),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_194),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_210),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_211),
.C(n_215),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_206),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_205),
.C(n_206),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_200),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_204),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g364 ( 
.A(n_206),
.Y(n_364)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.CI(n_209),
.CON(n_206),
.SN(n_206)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_208),
.C(n_209),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.CI(n_214),
.CON(n_211),
.SN(n_211)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_232),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_221),
.C(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_228),
.C(n_231),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g365 ( 
.A(n_223),
.Y(n_365)
);

FAx1_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.CI(n_226),
.CON(n_223),
.SN(n_223)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_224),
.B(n_225),
.C(n_226),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_239),
.C(n_244),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_239),
.B1(n_244),
.B2(n_245),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_235),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B(n_238),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_238),
.B(n_271),
.C(n_272),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_239),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_267),
.B2(n_279),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_268),
.C(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_252),
.C(n_260),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_260),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_256),
.C(n_259),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_258),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_266),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_265),
.C(n_266),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_264),
.Y(n_265)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_276),
.C(n_278),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_310),
.B2(n_311),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_282),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_301),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_301),
.C(n_310),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_293),
.C(n_294),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_288),
.C(n_290),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_300),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_295),
.Y(n_300)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_304),
.C(n_305),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_308),
.C(n_309),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_316),
.C(n_335),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_323),
.B2(n_335),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_321),
.C(n_322),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g367 ( 
.A(n_322),
.Y(n_367)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_326),
.C(n_327),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_330),
.B2(n_334),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_331),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_347),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_341),
.C(n_347),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_344),
.C(n_345),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_352),
.C(n_357),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_356),
.B2(n_357),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_362),
.Y(n_363)
);


endmodule