module fake_jpeg_28729_n_429 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_429);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_429;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_2),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_47),
.B(n_63),
.Y(n_132)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_49),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_60),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_51),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_52),
.Y(n_117)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_54),
.Y(n_148)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_55),
.Y(n_150)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_57),
.Y(n_125)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_59),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_14),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_13),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_12),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_65),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_12),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_28),
.B(n_35),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_26),
.B(n_37),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_75),
.Y(n_118)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_17),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_77),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_4),
.Y(n_137)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_35),
.B(n_2),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_85),
.Y(n_128)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_43),
.B(n_3),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_90),
.Y(n_140)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_32),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_91),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_94),
.Y(n_146)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_32),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_43),
.B(n_3),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_3),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_93),
.B1(n_68),
.B2(n_51),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_97),
.A2(n_119),
.B1(n_121),
.B2(n_76),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_114),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_56),
.A2(n_36),
.B1(n_21),
.B2(n_20),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_105),
.A2(n_106),
.B1(n_111),
.B2(n_123),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_61),
.A2(n_36),
.B1(n_21),
.B2(n_20),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_36),
.B1(n_21),
.B2(n_20),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_58),
.A2(n_46),
.B1(n_34),
.B2(n_38),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_142),
.B1(n_69),
.B2(n_54),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_62),
.A2(n_46),
.B1(n_38),
.B2(n_34),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_47),
.A2(n_38),
.B1(n_40),
.B2(n_39),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_SL g126 ( 
.A1(n_59),
.A2(n_41),
.B(n_42),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_135),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_91),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_137),
.Y(n_163)
);

OR2x4_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_37),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_53),
.A2(n_26),
.B1(n_41),
.B2(n_31),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_138),
.B1(n_52),
.B2(n_88),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_81),
.A2(n_41),
.B1(n_31),
.B2(n_6),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_71),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_142)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_67),
.B1(n_80),
.B2(n_57),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_152),
.A2(n_156),
.B1(n_165),
.B2(n_168),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_52),
.A3(n_77),
.B1(n_75),
.B2(n_48),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_155),
.B(n_162),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_55),
.B1(n_66),
.B2(n_87),
.Y(n_156)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_77),
.B1(n_75),
.B2(n_29),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_161),
.A2(n_177),
.B1(n_190),
.B2(n_112),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_164),
.A2(n_171),
.B1(n_188),
.B2(n_189),
.Y(n_228)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_59),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_170),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_121),
.A2(n_124),
.B1(n_145),
.B2(n_110),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_187),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_140),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_128),
.B(n_70),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_172),
.B(n_120),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

BUFx2_ASAP7_75t_SL g226 ( 
.A(n_173),
.Y(n_226)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_109),
.Y(n_175)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_175),
.B(n_117),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_96),
.B(n_41),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_182),
.Y(n_208)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_84),
.B1(n_91),
.B2(n_49),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_110),
.B(n_49),
.C(n_29),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_125),
.C(n_144),
.Y(n_198)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_135),
.A2(n_27),
.B1(n_5),
.B2(n_6),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_181),
.A2(n_186),
.B1(n_99),
.B2(n_192),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_100),
.B(n_27),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_184),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_125),
.A2(n_4),
.B(n_6),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_144),
.B(n_125),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_147),
.B1(n_122),
.B2(n_116),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_7),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_149),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_150),
.A2(n_8),
.B1(n_10),
.B2(n_101),
.Y(n_189)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_133),
.A2(n_8),
.B1(n_10),
.B2(n_116),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_97),
.B(n_10),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_194),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_113),
.B(n_103),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_195),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_133),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_129),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_197),
.B(n_198),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_144),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_199),
.B(n_157),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_139),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_202),
.B(n_176),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_205),
.A2(n_214),
.B(n_179),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_155),
.A2(n_98),
.B1(n_122),
.B2(n_112),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_212),
.B1(n_218),
.B2(n_231),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_158),
.A2(n_139),
.B(n_129),
.C(n_134),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_221),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_164),
.A2(n_98),
.B1(n_108),
.B2(n_134),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_156),
.A2(n_150),
.B1(n_107),
.B2(n_120),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_219),
.A2(n_154),
.B1(n_159),
.B2(n_166),
.Y(n_265)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_163),
.A2(n_99),
.B1(n_107),
.B2(n_158),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_234),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_163),
.A2(n_160),
.B1(n_192),
.B2(n_167),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_168),
.B1(n_182),
.B2(n_165),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_152),
.B(n_169),
.C(n_173),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_205),
.A2(n_185),
.B(n_175),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_236),
.A2(n_245),
.B(n_214),
.Y(n_279)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

OAI21x1_ASAP7_75t_R g292 ( 
.A1(n_237),
.A2(n_250),
.B(n_166),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_238),
.B(n_204),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_194),
.B(n_190),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_252),
.B1(n_210),
.B2(n_239),
.Y(n_278)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_195),
.B(n_194),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_207),
.B(n_170),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_246),
.B(n_247),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_206),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_197),
.Y(n_289)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_177),
.B(n_190),
.C(n_184),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_207),
.B(n_172),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_251),
.B(n_259),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_218),
.A2(n_186),
.B1(n_190),
.B2(n_151),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_178),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_213),
.Y(n_255)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_260),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_210),
.A2(n_177),
.B1(n_159),
.B2(n_180),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_258),
.A2(n_222),
.B1(n_229),
.B2(n_206),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_208),
.B(n_174),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_208),
.B(n_196),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_215),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_264),
.Y(n_284)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_200),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_221),
.B(n_191),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_266),
.B1(n_245),
.B2(n_258),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_206),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_202),
.C(n_198),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_281),
.C(n_285),
.Y(n_311)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_270),
.Y(n_305)
);

AOI32xp33_ASAP7_75t_L g271 ( 
.A1(n_240),
.A2(n_248),
.A3(n_263),
.B1(n_236),
.B2(n_253),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_279),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_247),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_278),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_264),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_275),
.B(n_290),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_279),
.A2(n_289),
.B(n_240),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_227),
.C(n_220),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_232),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_204),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_253),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_162),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_291),
.A2(n_293),
.B1(n_225),
.B2(n_250),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_265),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_251),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_297),
.B(n_316),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_300),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_243),
.B1(n_252),
.B2(n_239),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_301),
.A2(n_318),
.B1(n_274),
.B2(n_267),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_302),
.B(n_303),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_263),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_314),
.C(n_289),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_259),
.Y(n_306)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_272),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_317),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_313),
.B(n_225),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_260),
.Y(n_310)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_310),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_241),
.Y(n_312)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_253),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_315),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_283),
.B(n_238),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_284),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_320),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_292),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_253),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_312),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_299),
.A2(n_293),
.B1(n_283),
.B2(n_285),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_323),
.A2(n_325),
.B1(n_313),
.B2(n_316),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_328),
.C(n_329),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_299),
.A2(n_236),
.B1(n_250),
.B2(n_241),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_289),
.C(n_254),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_254),
.C(n_287),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_331),
.A2(n_333),
.B1(n_341),
.B2(n_320),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_286),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_337),
.C(n_338),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_301),
.A2(n_272),
.B1(n_277),
.B2(n_276),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_298),
.A2(n_249),
.B1(n_244),
.B2(n_242),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_334),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_262),
.C(n_256),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_303),
.B(n_235),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_320),
.A2(n_270),
.B1(n_268),
.B2(n_229),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_321),
.B(n_237),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_344),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_345),
.A2(n_296),
.B(n_305),
.Y(n_362)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_346),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_300),
.Y(n_347)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_347),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_330),
.A2(n_309),
.B(n_313),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_349),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_306),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_351),
.Y(n_371)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_355),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_336),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_308),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_357),
.Y(n_369)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_341),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_345),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_358),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_340),
.B(n_307),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_364),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_310),
.C(n_319),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_337),
.C(n_329),
.Y(n_370)
);

O2A1O1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_362),
.A2(n_363),
.B(n_343),
.C(n_342),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_325),
.A2(n_296),
.B(n_315),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_331),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_201),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_323),
.Y(n_377)
);

INVx2_ASAP7_75t_R g368 ( 
.A(n_348),
.Y(n_368)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_368),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_370),
.B(n_377),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_324),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_376),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_354),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_378),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_328),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_381),
.C(n_353),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_338),
.C(n_339),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_379),
.B(n_355),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_389),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_372),
.Y(n_384)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_384),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_387),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_353),
.C(n_339),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_371),
.B(n_352),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_372),
.B(n_370),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_392),
.Y(n_401)
);

NAND3xp33_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_359),
.C(n_358),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_366),
.B(n_373),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_393),
.A2(n_394),
.B(n_369),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_362),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_386),
.A2(n_363),
.B(n_374),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_397),
.B(n_404),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_380),
.C(n_376),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_400),
.C(n_388),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_375),
.C(n_367),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_349),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_402),
.B(n_405),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_384),
.A2(n_364),
.B1(n_357),
.B2(n_356),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_378),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_346),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_392),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_408),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_401),
.B(n_382),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_411),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_395),
.A2(n_361),
.B1(n_400),
.B2(n_405),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_344),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_413),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_407),
.A2(n_403),
.B1(n_399),
.B2(n_402),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_414),
.B(n_416),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_409),
.B(n_398),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_410),
.A2(n_209),
.B(n_224),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_419),
.A2(n_407),
.B(n_224),
.Y(n_421)
);

AOI321xp33_ASAP7_75t_SL g425 ( 
.A1(n_421),
.A2(n_417),
.A3(n_237),
.B1(n_201),
.B2(n_203),
.C(n_213),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_209),
.C(n_229),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_422),
.B(n_423),
.Y(n_424)
);

INVxp33_ASAP7_75t_SL g423 ( 
.A(n_415),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_425),
.A2(n_203),
.B(n_420),
.Y(n_426)
);

BUFx24_ASAP7_75t_SL g427 ( 
.A(n_426),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_427),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_428),
.A2(n_424),
.B(n_417),
.Y(n_429)
);


endmodule