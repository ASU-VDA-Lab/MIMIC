module real_aes_2886_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_56;
wire n_34;
wire n_55;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_53;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_37;
wire n_51;
wire n_54;
wire n_35;
wire n_42;
wire n_45;
wire n_39;
wire n_27;
wire n_23;
wire n_50;
wire n_38;
wire n_29;
wire n_20;
wire n_52;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx20_ASAP7_75t_R g43 ( .A(n_0), .Y(n_43) );
CKINVDCx20_ASAP7_75t_R g56 ( .A(n_1), .Y(n_56) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_2), .Y(n_24) );
NOR3xp33_ASAP7_75t_SL g22 ( .A(n_3), .B(n_7), .C(n_23), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_4), .Y(n_23) );
CKINVDCx20_ASAP7_75t_R g52 ( .A(n_5), .Y(n_52) );
NOR2xp33_ASAP7_75t_R g20 ( .A(n_6), .B(n_21), .Y(n_20) );
NAND3xp33_ASAP7_75t_SL g39 ( .A(n_6), .B(n_40), .C(n_41), .Y(n_39) );
NOR2xp33_ASAP7_75t_R g31 ( .A(n_8), .B(n_11), .Y(n_31) );
CKINVDCx20_ASAP7_75t_R g42 ( .A(n_8), .Y(n_42) );
AOI221xp5_ASAP7_75t_SL g44 ( .A1(n_9), .A2(n_13), .B1(n_45), .B2(n_46), .C(n_50), .Y(n_44) );
NOR2xp33_ASAP7_75t_R g29 ( .A(n_10), .B(n_30), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g40 ( .A(n_10), .Y(n_40) );
NAND2xp33_ASAP7_75t_SL g34 ( .A(n_11), .B(n_35), .Y(n_34) );
NOR2xp33_ASAP7_75t_R g45 ( .A(n_11), .B(n_36), .Y(n_45) );
NAND2xp33_ASAP7_75t_SL g47 ( .A(n_11), .B(n_48), .Y(n_47) );
CKINVDCx20_ASAP7_75t_R g55 ( .A(n_11), .Y(n_55) );
HB1xp67_ASAP7_75t_L g33 ( .A(n_12), .Y(n_33) );
CKINVDCx20_ASAP7_75t_R g25 ( .A(n_14), .Y(n_25) );
NAND2xp33_ASAP7_75t_SL g49 ( .A(n_14), .B(n_38), .Y(n_49) );
NAND2xp33_ASAP7_75t_SL g51 ( .A(n_14), .B(n_20), .Y(n_51) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_15), .Y(n_27) );
NOR2xp33_ASAP7_75t_R g41 ( .A(n_15), .B(n_42), .Y(n_41) );
OAI221xp5_ASAP7_75t_SL g16 ( .A1(n_17), .A2(n_32), .B1(n_34), .B2(n_43), .C(n_44), .Y(n_16) );
NAND2xp33_ASAP7_75t_SL g17 ( .A(n_18), .B(n_26), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
NAND2xp33_ASAP7_75t_SL g19 ( .A(n_20), .B(n_25), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g38 ( .A(n_21), .Y(n_38) );
NAND2xp33_ASAP7_75t_SL g21 ( .A(n_22), .B(n_24), .Y(n_21) );
NAND2xp33_ASAP7_75t_SL g37 ( .A(n_25), .B(n_38), .Y(n_37) );
CKINVDCx20_ASAP7_75t_R g53 ( .A(n_26), .Y(n_53) );
NOR2xp33_ASAP7_75t_R g26 ( .A(n_27), .B(n_28), .Y(n_26) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_29), .Y(n_28) );
CKINVDCx14_ASAP7_75t_R g30 ( .A(n_31), .Y(n_30) );
CKINVDCx20_ASAP7_75t_R g32 ( .A(n_33), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g35 ( .A(n_36), .Y(n_35) );
OR2x2_ASAP7_75t_L g36 ( .A(n_37), .B(n_39), .Y(n_36) );
NOR2xp33_ASAP7_75t_R g48 ( .A(n_39), .B(n_49), .Y(n_48) );
CKINVDCx14_ASAP7_75t_R g46 ( .A(n_47), .Y(n_46) );
NAND2xp33_ASAP7_75t_SL g54 ( .A(n_48), .B(n_55), .Y(n_54) );
OAI32xp33_ASAP7_75t_L g50 ( .A1(n_51), .A2(n_52), .A3(n_53), .B1(n_54), .B2(n_56), .Y(n_50) );
endmodule