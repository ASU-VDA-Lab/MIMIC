module fake_jpeg_6859_n_250 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_0),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_18),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_34),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_27),
.B1(n_25),
.B2(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_61),
.B1(n_21),
.B2(n_32),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_64),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_27),
.B1(n_25),
.B2(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_23),
.B1(n_19),
.B2(n_35),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_70),
.B1(n_23),
.B2(n_32),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_33),
.B1(n_20),
.B2(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_88),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_SL g73 ( 
.A1(n_70),
.A2(n_33),
.B(n_43),
.C(n_45),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_50),
.B(n_60),
.Y(n_96)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_42),
.Y(n_76)
);

OAI211xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_62),
.B(n_63),
.C(n_68),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_78),
.B1(n_89),
.B2(n_68),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_21),
.B1(n_32),
.B2(n_29),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_66),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_26),
.B1(n_31),
.B2(n_16),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_93),
.Y(n_109)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_56),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_98),
.B(n_101),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_73),
.B1(n_87),
.B2(n_84),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_107),
.B1(n_80),
.B2(n_94),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_67),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_85),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_64),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_111),
.C(n_56),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_53),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_106),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_69),
.B1(n_50),
.B2(n_65),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_118),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_88),
.B1(n_80),
.B2(n_93),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_59),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_59),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_116),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_72),
.B(n_14),
.Y(n_116)
);

BUFx4f_ASAP7_75t_SL g117 ( 
.A(n_81),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_86),
.A2(n_56),
.B1(n_42),
.B2(n_31),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_132),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_112),
.B1(n_98),
.B2(n_97),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_85),
.B(n_90),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_129),
.B(n_96),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_133),
.B(n_142),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_31),
.B(n_81),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_0),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_14),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_109),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_26),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_108),
.B(n_1),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_120),
.B(n_140),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_156),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_129),
.B1(n_132),
.B2(n_134),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_95),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_97),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_103),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_158),
.C(n_165),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_97),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_95),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_97),
.B1(n_112),
.B2(n_98),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_133),
.B(n_142),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_163),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_105),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_117),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_116),
.C(n_110),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_171),
.B1(n_182),
.B2(n_187),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_151),
.B(n_146),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_122),
.B1(n_126),
.B2(n_138),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_122),
.B1(n_126),
.B2(n_130),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_183),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_179),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_136),
.B1(n_130),
.B2(n_139),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_109),
.B(n_135),
.C(n_113),
.D(n_117),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_110),
.C(n_104),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_185),
.C(n_167),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_102),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_197),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_154),
.B1(n_156),
.B2(n_151),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_181),
.B1(n_175),
.B2(n_184),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_194),
.Y(n_208)
);

XOR2x2_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_147),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_201),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_169),
.B(n_155),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_204),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_202),
.C(n_165),
.Y(n_215)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_180),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_153),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_208),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_187),
.B1(n_180),
.B2(n_177),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_217),
.B1(n_191),
.B2(n_196),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_210),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_176),
.B1(n_166),
.B2(n_161),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_195),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_216),
.C(n_200),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_174),
.C(n_2),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_219),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_221),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_189),
.C(n_202),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_224),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_192),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_192),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_225),
.A2(n_226),
.B(n_1),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_203),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_212),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_213),
.B1(n_214),
.B2(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_230),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_217),
.B(n_216),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_232),
.B(n_6),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_227),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_7),
.Y(n_243)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_224),
.B(n_9),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_239),
.B(n_240),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_231),
.Y(n_239)
);

AOI21x1_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_13),
.B(n_9),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_241),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_7),
.C(n_9),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_237),
.C(n_11),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_10),
.B(n_11),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_247),
.B(n_10),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_13),
.Y(n_250)
);


endmodule