module fake_netlist_1_1959_n_721 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_721);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_721;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_17), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_31), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_46), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_24), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_14), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_8), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_55), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_0), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_15), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_1), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_9), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_68), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_49), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_39), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_57), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_25), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_58), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_42), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_78), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_61), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_45), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_75), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_34), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_12), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_19), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_43), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_14), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_23), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_59), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_76), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_37), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_54), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_35), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_23), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_48), .Y(n_115) );
INVxp33_ASAP7_75t_SL g116 ( .A(n_52), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_5), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_51), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_73), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_70), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_64), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_22), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_17), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_13), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_4), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_36), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_29), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_8), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_82), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_124), .B(n_0), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_124), .B(n_1), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_97), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_97), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_80), .B(n_2), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_80), .B(n_2), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_109), .B(n_3), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_93), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_93), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_94), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_95), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_95), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_84), .B(n_3), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_96), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_96), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_98), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_85), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_98), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_99), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_99), .Y(n_155) );
INVxp67_ASAP7_75t_L g156 ( .A(n_84), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_100), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_100), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_103), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_103), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_126), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
CKINVDCx11_ASAP7_75t_R g163 ( .A(n_101), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_87), .B(n_4), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_127), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_85), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g167 ( .A1(n_87), .A2(n_6), .B1(n_7), .B2(n_9), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_127), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_106), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_111), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_113), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_118), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_119), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_130), .B(n_128), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_134), .B(n_120), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_130), .B(n_128), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_133), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
INVx4_ASAP7_75t_L g183 ( .A(n_134), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_130), .B(n_102), .Y(n_184) );
INVxp67_ASAP7_75t_L g185 ( .A(n_131), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_133), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_134), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_133), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_163), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_136), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_156), .B(n_121), .Y(n_193) );
AND2x6_ASAP7_75t_L g194 ( .A(n_136), .B(n_125), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_156), .B(n_92), .Y(n_195) );
INVxp67_ASAP7_75t_L g196 ( .A(n_131), .Y(n_196) );
OAI22xp33_ASAP7_75t_SL g197 ( .A1(n_166), .A2(n_108), .B1(n_105), .B2(n_90), .Y(n_197) );
OR2x6_ASAP7_75t_L g198 ( .A(n_131), .B(n_125), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_129), .B(n_123), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_136), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_129), .B(n_91), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_135), .B(n_123), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_135), .B(n_112), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_136), .B(n_89), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_133), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_133), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_137), .B(n_116), .Y(n_207) );
AND2x6_ASAP7_75t_L g208 ( .A(n_136), .B(n_89), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_151), .Y(n_209) );
INVx5_ASAP7_75t_L g210 ( .A(n_145), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_133), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_145), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_137), .B(n_112), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_140), .B(n_92), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_140), .B(n_146), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_145), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_151), .Y(n_217) );
NAND3xp33_ASAP7_75t_L g218 ( .A(n_141), .B(n_88), .C(n_117), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_151), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_146), .B(n_114), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_145), .Y(n_221) );
OAI22xp33_ASAP7_75t_L g222 ( .A1(n_141), .A2(n_122), .B1(n_107), .B2(n_104), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_158), .B(n_115), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_158), .B(n_159), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_159), .B(n_110), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_145), .Y(n_226) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_148), .A2(n_81), .B(n_40), .Y(n_227) );
NAND3xp33_ASAP7_75t_SL g228 ( .A(n_148), .B(n_10), .C(n_11), .Y(n_228) );
INVxp67_ASAP7_75t_SL g229 ( .A(n_151), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_161), .B(n_10), .Y(n_230) );
OAI221xp5_ASAP7_75t_L g231 ( .A1(n_164), .A2(n_11), .B1(n_12), .B2(n_13), .C(n_15), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_161), .A2(n_16), .B1(n_18), .B2(n_19), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_168), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_171), .A2(n_16), .B1(n_18), .B2(n_20), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_168), .B(n_20), .Y(n_235) );
OAI21xp33_ASAP7_75t_SL g236 ( .A1(n_175), .A2(n_164), .B(n_168), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_194), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_213), .B(n_168), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_217), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_217), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_183), .Y(n_241) );
NOR2x1p5_ASAP7_75t_L g242 ( .A(n_190), .B(n_166), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_213), .B(n_173), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_217), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_194), .A2(n_173), .B1(n_171), .B2(n_172), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_233), .Y(n_246) );
AND3x1_ASAP7_75t_L g247 ( .A(n_232), .B(n_170), .C(n_172), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_229), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_190), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_194), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_184), .A2(n_173), .B1(n_171), .B2(n_167), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_215), .Y(n_252) );
INVx5_ASAP7_75t_L g253 ( .A(n_194), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_215), .B(n_173), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_215), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_209), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_214), .B(n_173), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_198), .B(n_172), .Y(n_258) );
BUFx4f_ASAP7_75t_L g259 ( .A(n_194), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_214), .B(n_171), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_194), .Y(n_261) );
INVxp33_ASAP7_75t_L g262 ( .A(n_177), .Y(n_262) );
BUFx4f_ASAP7_75t_SL g263 ( .A(n_182), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_184), .A2(n_171), .B1(n_167), .B2(n_170), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_208), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_187), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_187), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_183), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_187), .Y(n_269) );
INVx4_ASAP7_75t_L g270 ( .A(n_208), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_209), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_219), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_219), .Y(n_273) );
BUFx12f_ASAP7_75t_L g274 ( .A(n_198), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_200), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_183), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_193), .B(n_170), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_221), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_207), .B(n_150), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_198), .B(n_150), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_198), .B(n_174), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_188), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_188), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_185), .B(n_150), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_208), .A2(n_230), .B1(n_204), .B2(n_179), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_182), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_221), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_208), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_196), .A2(n_154), .B1(n_165), .B2(n_162), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_203), .B(n_154), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_188), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_174), .B(n_154), .Y(n_292) );
INVx4_ASAP7_75t_L g293 ( .A(n_208), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_174), .B(n_155), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_179), .B(n_155), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_179), .B(n_155), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_191), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_191), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_208), .A2(n_138), .B1(n_165), .B2(n_162), .Y(n_299) );
NOR2x1_ASAP7_75t_L g300 ( .A(n_218), .B(n_138), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_226), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_178), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_178), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_277), .A2(n_178), .B(n_191), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_266), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_281), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_270), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_263), .Y(n_308) );
NAND2x1_ASAP7_75t_L g309 ( .A(n_270), .B(n_204), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_236), .A2(n_197), .B(n_222), .C(n_231), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_281), .A2(n_204), .B1(n_228), .B2(n_230), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_281), .B(n_199), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_262), .A2(n_199), .B1(n_202), .B2(n_220), .C(n_201), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_290), .A2(n_224), .B(n_195), .Y(n_314) );
OAI21x1_ASAP7_75t_SL g315 ( .A1(n_302), .A2(n_225), .B(n_223), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_280), .B(n_202), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_302), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_280), .B(n_235), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_270), .B(n_234), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_266), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_237), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_267), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
OR2x2_ASAP7_75t_SL g324 ( .A(n_274), .B(n_138), .Y(n_324) );
INVx4_ASAP7_75t_L g325 ( .A(n_293), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_303), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_274), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_293), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_285), .A2(n_139), .B1(n_142), .B2(n_143), .Y(n_329) );
BUFx4_ASAP7_75t_SL g330 ( .A(n_249), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_267), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_280), .B(n_227), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_280), .B(n_157), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_237), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_250), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_269), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_286), .Y(n_337) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_236), .A2(n_157), .B(n_165), .C(n_162), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_250), .Y(n_339) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_259), .B(n_144), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_286), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_258), .A2(n_227), .B1(n_169), .B2(n_142), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_261), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_303), .A2(n_144), .B1(n_157), .B2(n_160), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_258), .B(n_227), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_258), .B(n_160), .Y(n_346) );
O2A1O1Ixp33_ASAP7_75t_L g347 ( .A1(n_295), .A2(n_139), .B(n_142), .C(n_143), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_258), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_249), .Y(n_349) );
NOR2x1_ASAP7_75t_L g350 ( .A(n_261), .B(n_160), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_269), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_292), .B(n_139), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_246), .Y(n_353) );
NOR2xp33_ASAP7_75t_SL g354 ( .A(n_259), .B(n_143), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_265), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_265), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_246), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_253), .B(n_169), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_353), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_337), .A2(n_292), .B1(n_294), .B2(n_259), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_305), .Y(n_361) );
NAND3xp33_ASAP7_75t_SL g362 ( .A(n_349), .B(n_251), .C(n_264), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_312), .B(n_292), .Y(n_363) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_341), .A2(n_288), .B1(n_255), .B2(n_252), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_305), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_328), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_342), .A2(n_275), .B(n_243), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_SL g368 ( .A1(n_310), .A2(n_284), .B(n_245), .C(n_279), .Y(n_368) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_308), .A2(n_288), .B1(n_255), .B2(n_252), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_319), .A2(n_242), .B1(n_294), .B2(n_248), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_305), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_330), .Y(n_372) );
AO22x2_ASAP7_75t_L g373 ( .A1(n_315), .A2(n_247), .B1(n_294), .B2(n_275), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_327), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_327), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_340), .A2(n_296), .B1(n_299), .B2(n_289), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_353), .Y(n_377) );
OR2x6_ASAP7_75t_L g378 ( .A(n_306), .B(n_238), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_351), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_325), .B(n_253), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_319), .A2(n_242), .B1(n_248), .B2(n_298), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_319), .A2(n_283), .B1(n_298), .B2(n_297), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g383 ( .A1(n_306), .A2(n_257), .B1(n_260), .B2(n_253), .Y(n_383) );
NOR2x1_ASAP7_75t_R g384 ( .A(n_319), .B(n_253), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_315), .A2(n_253), .B1(n_291), .B2(n_241), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_325), .B(n_253), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_328), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_340), .A2(n_272), .B1(n_271), .B2(n_254), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_348), .A2(n_276), .B1(n_297), .B2(n_283), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_324), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_357), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_312), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_361), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_373), .A2(n_324), .B1(n_348), .B2(n_318), .Y(n_395) );
AO21x1_ASAP7_75t_L g396 ( .A1(n_367), .A2(n_345), .B(n_332), .Y(n_396) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_362), .A2(n_313), .B(n_316), .C(n_329), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
OR2x6_ASAP7_75t_L g399 ( .A(n_378), .B(n_317), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_361), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_373), .A2(n_340), .B1(n_357), .B2(n_311), .Y(n_402) );
BUFx8_ASAP7_75t_SL g403 ( .A(n_372), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_379), .B(n_316), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_373), .A2(n_300), .B1(n_352), .B2(n_333), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_373), .A2(n_300), .B1(n_352), .B2(n_333), .Y(n_406) );
OR2x2_ASAP7_75t_SL g407 ( .A(n_359), .B(n_144), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_379), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_365), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_370), .A2(n_322), .B1(n_336), .B2(n_320), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_390), .A2(n_354), .B1(n_326), .B2(n_317), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_378), .A2(n_326), .B1(n_346), .B2(n_344), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_381), .A2(n_320), .B1(n_336), .B2(n_322), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_375), .A2(n_354), .B1(n_325), .B2(n_328), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_365), .B(n_351), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_371), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_386), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_371), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_374), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_378), .Y(n_420) );
AOI322xp5_ASAP7_75t_L g421 ( .A1(n_359), .A2(n_132), .A3(n_331), .B1(n_309), .B2(n_21), .C1(n_22), .C2(n_153), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_386), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_397), .B(n_393), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_398), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_408), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_398), .B(n_392), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_399), .A2(n_378), .B1(n_392), .B2(n_377), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_397), .A2(n_382), .B1(n_363), .B2(n_338), .C(n_391), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_400), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_415), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_399), .A2(n_378), .B1(n_391), .B2(n_377), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_415), .B(n_367), .Y(n_432) );
NAND4xp25_ASAP7_75t_L g433 ( .A(n_421), .B(n_368), .C(n_360), .D(n_314), .Y(n_433) );
OAI211xp5_ASAP7_75t_L g434 ( .A1(n_421), .A2(n_372), .B(n_385), .C(n_389), .Y(n_434) );
AND2x4_ASAP7_75t_SL g435 ( .A(n_399), .B(n_386), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_404), .B(n_364), .Y(n_436) );
OAI22xp33_ASAP7_75t_L g437 ( .A1(n_399), .A2(n_376), .B1(n_388), .B2(n_369), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_402), .A2(n_383), .B1(n_331), .B2(n_350), .Y(n_438) );
AOI33xp33_ASAP7_75t_L g439 ( .A1(n_405), .A2(n_406), .A3(n_410), .B1(n_132), .B2(n_413), .B3(n_411), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_400), .B(n_366), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_401), .B(n_366), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_401), .B(n_409), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_414), .B(n_366), .Y(n_443) );
OAI31xp33_ASAP7_75t_SL g444 ( .A1(n_395), .A2(n_384), .A3(n_386), .B(n_350), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_412), .A2(n_347), .B(n_304), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_404), .B(n_384), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_394), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_422), .B(n_387), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_419), .B(n_309), .Y(n_449) );
OAI22xp33_ASAP7_75t_L g450 ( .A1(n_399), .A2(n_380), .B1(n_325), .B2(n_387), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_409), .B(n_387), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_420), .A2(n_169), .B1(n_132), .B2(n_149), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_420), .A2(n_169), .B1(n_149), .B2(n_153), .Y(n_453) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_396), .A2(n_186), .B(n_189), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_422), .A2(n_169), .B1(n_149), .B2(n_153), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_396), .A2(n_149), .B1(n_147), .B2(n_153), .C(n_169), .Y(n_456) );
OAI31xp33_ASAP7_75t_SL g457 ( .A1(n_416), .A2(n_271), .A3(n_272), .B(n_240), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_447), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_424), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_430), .B(n_416), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_447), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_424), .B(n_418), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_442), .B(n_418), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_442), .B(n_408), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_423), .B(n_394), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_426), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_432), .B(n_429), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_429), .B(n_407), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_444), .B(n_422), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_432), .B(n_407), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g471 ( .A1(n_431), .A2(n_435), .B1(n_427), .B2(n_434), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_425), .B(n_422), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_425), .B(n_417), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_425), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_447), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_426), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_431), .A2(n_417), .B1(n_380), .B2(n_339), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_440), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_440), .B(n_147), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_451), .B(n_147), .Y(n_480) );
OAI321xp33_ASAP7_75t_L g481 ( .A1(n_427), .A2(n_147), .A3(n_149), .B1(n_153), .B2(n_169), .C(n_380), .Y(n_481) );
AOI222xp33_ASAP7_75t_L g482 ( .A1(n_428), .A2(n_153), .B1(n_149), .B2(n_147), .C1(n_21), .C2(n_403), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_454), .Y(n_483) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_447), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_451), .B(n_147), .Y(n_485) );
NAND5xp2_ASAP7_75t_L g486 ( .A(n_444), .B(n_276), .C(n_240), .D(n_192), .E(n_212), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_448), .B(n_153), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_441), .B(n_149), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_448), .B(n_147), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_454), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_441), .B(n_26), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_454), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_454), .Y(n_493) );
OAI31xp33_ASAP7_75t_L g494 ( .A1(n_437), .A2(n_307), .A3(n_323), .B(n_241), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_436), .B(n_343), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_439), .B(n_343), .Y(n_496) );
OAI221xp5_ASAP7_75t_L g497 ( .A1(n_449), .A2(n_358), .B1(n_355), .B2(n_323), .C(n_307), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g498 ( .A1(n_433), .A2(n_192), .B1(n_176), .B2(n_212), .C(n_226), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_447), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_448), .B(n_27), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_446), .B(n_355), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_448), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_435), .Y(n_504) );
AOI222xp33_ASAP7_75t_L g505 ( .A1(n_435), .A2(n_321), .B1(n_339), .B2(n_335), .C1(n_334), .C2(n_307), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_445), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_445), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_482), .B(n_457), .C(n_433), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_467), .B(n_438), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_466), .B(n_457), .Y(n_511) );
AOI33xp33_ASAP7_75t_L g512 ( .A1(n_471), .A2(n_459), .A3(n_467), .B1(n_476), .B2(n_507), .B3(n_506), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_502), .B(n_456), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_464), .B(n_450), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_464), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_462), .Y(n_516) );
NAND4xp25_ASAP7_75t_L g517 ( .A(n_482), .B(n_453), .C(n_452), .D(n_455), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_463), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_478), .B(n_189), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_462), .Y(n_520) );
AOI31xp33_ASAP7_75t_L g521 ( .A1(n_469), .A2(n_28), .A3(n_30), .B(n_32), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_502), .B(n_211), .Y(n_522) );
NOR2xp33_ASAP7_75t_SL g523 ( .A(n_494), .B(n_328), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_476), .B(n_186), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_460), .B(n_211), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_474), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_486), .A2(n_356), .B1(n_343), .B2(n_339), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_474), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_468), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_501), .B(n_33), .Y(n_530) );
AOI211xp5_ASAP7_75t_L g531 ( .A1(n_486), .A2(n_176), .B(n_181), .C(n_180), .Y(n_531) );
NAND2x1_ASAP7_75t_L g532 ( .A(n_477), .B(n_328), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_465), .B(n_205), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_470), .B(n_506), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_470), .B(n_205), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_468), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_477), .A2(n_307), .B1(n_323), .B2(n_335), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_487), .B(n_206), .C(n_181), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_507), .B(n_206), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_473), .B(n_206), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_474), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_472), .B(n_206), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_472), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_473), .B(n_206), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_479), .B(n_181), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_479), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_485), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_483), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_485), .B(n_181), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_504), .B(n_181), .Y(n_551) );
INVx3_ASAP7_75t_SL g552 ( .A(n_500), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_504), .B(n_180), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_480), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_504), .B(n_38), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_483), .B(n_180), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_480), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_503), .B(n_180), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_492), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_488), .B(n_180), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_503), .B(n_226), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_488), .B(n_226), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_492), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_490), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_491), .B(n_226), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_490), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_518), .B(n_529), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_552), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_536), .B(n_503), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_546), .Y(n_570) );
AOI21xp33_ASAP7_75t_SL g571 ( .A1(n_552), .A2(n_494), .B(n_500), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_509), .B(n_481), .C(n_489), .Y(n_572) );
NAND4xp75_ASAP7_75t_L g573 ( .A(n_511), .B(n_491), .C(n_496), .D(n_495), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_530), .B(n_500), .Y(n_574) );
NAND2x1_ASAP7_75t_L g575 ( .A(n_521), .B(n_500), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_515), .B(n_493), .Y(n_576) );
OR3x2_ASAP7_75t_L g577 ( .A(n_517), .B(n_493), .C(n_481), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_534), .B(n_461), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_546), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_534), .B(n_487), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_543), .B(n_461), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_516), .B(n_489), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_531), .A2(n_487), .B1(n_489), .B2(n_505), .Y(n_583) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_538), .B(n_487), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_520), .B(n_489), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_510), .B(n_499), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_510), .B(n_484), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_554), .B(n_475), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_547), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_549), .B(n_475), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_549), .B(n_475), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_564), .B(n_475), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_508), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_508), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_564), .B(n_458), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_566), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_566), .B(n_458), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_533), .A2(n_497), .B(n_505), .C(n_498), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_526), .B(n_458), .Y(n_599) );
OAI31xp33_ASAP7_75t_L g600 ( .A1(n_523), .A2(n_323), .A3(n_335), .B(n_334), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_532), .B(n_41), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_526), .B(n_541), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_541), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_548), .Y(n_604) );
NAND4xp25_ASAP7_75t_L g605 ( .A(n_512), .B(n_216), .C(n_334), .D(n_321), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_532), .A2(n_356), .B(n_343), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_557), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_512), .B(n_210), .C(n_216), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_535), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_559), .B(n_44), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_514), .B(n_47), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_559), .B(n_50), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_539), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_563), .B(n_53), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_563), .B(n_56), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_535), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_528), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_513), .B(n_62), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_513), .A2(n_216), .B1(n_210), .B2(n_256), .C(n_273), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_528), .B(n_63), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_604), .B(n_539), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_586), .B(n_561), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_589), .B(n_542), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_578), .B(n_556), .Y(n_624) );
AOI221x1_ASAP7_75t_L g625 ( .A1(n_572), .A2(n_555), .B1(n_525), .B2(n_524), .C(n_565), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_594), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_607), .B(n_542), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_587), .B(n_561), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_594), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_567), .B(n_556), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_575), .A2(n_522), .B1(n_553), .B2(n_551), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_596), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_609), .B(n_522), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_576), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_570), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_576), .B(n_558), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_616), .B(n_558), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_593), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_578), .B(n_519), .Y(n_639) );
AOI21xp33_ASAP7_75t_SL g640 ( .A1(n_568), .A2(n_537), .B(n_519), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_570), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_602), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_571), .A2(n_540), .B1(n_544), .B2(n_550), .C(n_545), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_569), .B(n_553), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_581), .B(n_551), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_584), .B(n_560), .Y(n_646) );
NAND2x1p5_ASAP7_75t_L g647 ( .A(n_575), .B(n_562), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_602), .B(n_527), .Y(n_648) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_605), .B(n_256), .C(n_273), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_603), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_581), .B(n_65), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_580), .B(n_66), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_613), .B(n_67), .Y(n_653) );
INVxp67_ASAP7_75t_SL g654 ( .A(n_579), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_577), .A2(n_356), .B1(n_343), .B2(n_321), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_582), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_618), .A2(n_241), .B(n_268), .C(n_291), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_585), .B(n_69), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_608), .A2(n_210), .B(n_291), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_598), .A2(n_282), .B(n_268), .C(n_301), .Y(n_660) );
AOI22x1_ASAP7_75t_L g661 ( .A1(n_568), .A2(n_356), .B1(n_72), .B2(n_74), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_591), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_573), .B(n_71), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_591), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_573), .B(n_77), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_595), .Y(n_666) );
OAI211xp5_ASAP7_75t_SL g667 ( .A1(n_583), .A2(n_268), .B(n_282), .C(n_278), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_595), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_590), .B(n_79), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_601), .B(n_356), .Y(n_670) );
XNOR2x1_ASAP7_75t_L g671 ( .A(n_597), .B(n_282), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_590), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_574), .A2(n_239), .B(n_244), .C(n_301), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_577), .A2(n_210), .B1(n_278), .B2(n_287), .Y(n_674) );
OAI21xp33_ASAP7_75t_SL g675 ( .A1(n_600), .A2(n_239), .B(n_244), .Y(n_675) );
NOR3x1_ASAP7_75t_L g676 ( .A(n_588), .B(n_210), .C(n_287), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_592), .Y(n_677) );
OAI211xp5_ASAP7_75t_L g678 ( .A1(n_611), .A2(n_597), .B(n_619), .C(n_592), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_599), .B(n_617), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_601), .A2(n_606), .B(n_615), .Y(n_680) );
OAI221xp5_ASAP7_75t_SL g681 ( .A1(n_599), .A2(n_610), .B1(n_612), .B2(n_614), .C(n_615), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_579), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_610), .Y(n_683) );
AOI222xp33_ASAP7_75t_L g684 ( .A1(n_634), .A2(n_656), .B1(n_672), .B2(n_643), .C1(n_667), .C2(n_668), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_630), .Y(n_685) );
OAI21xp5_ASAP7_75t_L g686 ( .A1(n_647), .A2(n_631), .B(n_675), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_647), .A2(n_681), .B1(n_672), .B2(n_678), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_648), .A2(n_665), .B1(n_663), .B2(n_646), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_651), .Y(n_689) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_663), .B(n_665), .Y(n_690) );
AOI21xp33_ASAP7_75t_L g691 ( .A1(n_660), .A2(n_646), .B(n_657), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_676), .B(n_666), .Y(n_692) );
AOI22x1_ASAP7_75t_L g693 ( .A1(n_680), .A2(n_651), .B1(n_659), .B2(n_654), .Y(n_693) );
AOI321xp33_ASAP7_75t_L g694 ( .A1(n_640), .A2(n_674), .A3(n_623), .B1(n_649), .B2(n_627), .C(n_633), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_649), .A2(n_673), .B(n_624), .C(n_642), .Y(n_695) );
OA22x2_ASAP7_75t_L g696 ( .A1(n_625), .A2(n_664), .B1(n_662), .B2(n_670), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_679), .Y(n_697) );
AOI31xp33_ASAP7_75t_L g698 ( .A1(n_671), .A2(n_652), .A3(n_655), .B(n_601), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_684), .B(n_624), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_687), .A2(n_677), .B1(n_638), .B2(n_632), .C(n_650), .Y(n_700) );
AOI211xp5_ASAP7_75t_L g701 ( .A1(n_695), .A2(n_652), .B(n_669), .C(n_653), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_691), .A2(n_629), .B1(n_626), .B2(n_639), .C(n_621), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_692), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_693), .A2(n_683), .B1(n_628), .B2(n_622), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_686), .A2(n_654), .B(n_661), .Y(n_705) );
OAI211xp5_ASAP7_75t_L g706 ( .A1(n_694), .A2(n_658), .B(n_644), .C(n_637), .Y(n_706) );
NOR3xp33_ASAP7_75t_L g707 ( .A(n_700), .B(n_690), .C(n_698), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_703), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_699), .A2(n_696), .B1(n_688), .B2(n_685), .Y(n_709) );
OA22x2_ASAP7_75t_L g710 ( .A1(n_706), .A2(n_692), .B1(n_689), .B2(n_696), .Y(n_710) );
BUFx2_ASAP7_75t_L g711 ( .A(n_702), .Y(n_711) );
AO22x2_ASAP7_75t_L g712 ( .A1(n_709), .A2(n_705), .B1(n_697), .B2(n_704), .Y(n_712) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_711), .A2(n_701), .B1(n_645), .B2(n_682), .Y(n_713) );
NAND5xp2_ASAP7_75t_L g714 ( .A(n_707), .B(n_612), .C(n_614), .D(n_620), .E(n_645), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_712), .A2(n_710), .B1(n_708), .B2(n_636), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_713), .A2(n_635), .B(n_641), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_715), .A2(n_714), .B(n_620), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_716), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_718), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_719), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_720), .A2(n_717), .B1(n_635), .B2(n_641), .Y(n_721) );
endmodule