module real_jpeg_25816_n_19 (n_17, n_123, n_8, n_116, n_0, n_2, n_125, n_10, n_9, n_12, n_124, n_6, n_121, n_11, n_14, n_7, n_117, n_18, n_3, n_119, n_5, n_4, n_115, n_122, n_1, n_118, n_16, n_15, n_13, n_120, n_19);

input n_17;
input n_123;
input n_8;
input n_116;
input n_0;
input n_2;
input n_125;
input n_10;
input n_9;
input n_12;
input n_124;
input n_6;
input n_121;
input n_11;
input n_14;
input n_7;
input n_117;
input n_18;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_118;
input n_16;
input n_15;
input n_13;
input n_120;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_1),
.B(n_93),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_2),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_4),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_5),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_7),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_8),
.B(n_66),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_9),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_33),
.C(n_110),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_13),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_13),
.B(n_83),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_14),
.B(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_15),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_15),
.B(n_99),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_16),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_17),
.B(n_35),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_22),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_26),
.B(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_28),
.B(n_106),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_29),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_29),
.B(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B(n_109),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_103),
.B(n_108),
.Y(n_37)
);

OAI321xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_92),
.A3(n_98),
.B1(n_101),
.B2(n_102),
.C(n_115),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_86),
.B(n_91),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_82),
.B(n_85),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_76),
.B(n_81),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_49),
.B(n_75),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_69),
.B(n_74),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_65),
.B(n_68),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_57),
.B(n_64),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_71),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_78),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_79),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_87),
.B(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_116),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_117),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_118),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_119),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_120),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_121),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_122),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_123),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_124),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_125),
.Y(n_100)
);


endmodule