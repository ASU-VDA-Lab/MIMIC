module real_aes_3777_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_1106, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_1105, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_1106;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_1105;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_357;
wire n_635;
wire n_673;
wire n_386;
wire n_1067;
wire n_518;
wire n_792;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_948;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_815;
wire n_638;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_892;
wire n_370;
wire n_994;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_1086;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_1081;
wire n_973;
wire n_1084;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1103;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_1079;
wire n_843;
wire n_810;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_749;
wire n_358;
wire n_385;
wire n_663;
wire n_1056;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_314;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_359;
wire n_456;
wire n_717;
wire n_982;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_307;
wire n_1101;
wire n_601;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_1061;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_0), .A2(n_23), .B1(n_659), .B2(n_660), .Y(n_658) );
INVx1_ASAP7_75t_SL g598 ( .A(n_1), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_1), .A2(n_50), .B1(n_839), .B2(n_843), .Y(n_838) );
INVx1_ASAP7_75t_L g654 ( .A(n_2), .Y(n_654) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_3), .Y(n_825) );
AND2x4_ASAP7_75t_L g833 ( .A(n_3), .B(n_834), .Y(n_833) );
AND2x4_ASAP7_75t_L g842 ( .A(n_3), .B(n_289), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_4), .A2(n_111), .B1(n_517), .B2(n_518), .Y(n_546) );
XOR2x2_ASAP7_75t_L g423 ( .A(n_5), .B(n_424), .Y(n_423) );
XNOR2xp5_ASAP7_75t_L g491 ( .A(n_5), .B(n_424), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_6), .A2(n_189), .B1(n_502), .B2(n_1087), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_7), .A2(n_155), .B1(n_363), .B2(n_634), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_8), .A2(n_182), .B1(n_514), .B2(n_515), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_9), .A2(n_122), .B1(n_857), .B2(n_858), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_10), .A2(n_121), .B1(n_749), .B2(n_750), .Y(n_748) );
AOI21xp33_ASAP7_75t_SL g1070 ( .A1(n_11), .A2(n_801), .B(n_1071), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_12), .A2(n_277), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI21xp33_ASAP7_75t_SL g661 ( .A1(n_13), .A2(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g615 ( .A(n_14), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_15), .A2(n_237), .B1(n_331), .B2(n_431), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_16), .A2(n_691), .B(n_692), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_17), .A2(n_257), .B1(n_502), .B2(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g437 ( .A(n_18), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_19), .A2(n_31), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g707 ( .A(n_20), .Y(n_707) );
AO22x1_ASAP7_75t_L g522 ( .A1(n_21), .A2(n_166), .B1(n_523), .B2(n_524), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_22), .A2(n_157), .B1(n_362), .B2(n_763), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_24), .A2(n_261), .B1(n_447), .B2(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_25), .A2(n_211), .B1(n_427), .B2(n_634), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_26), .A2(n_125), .B1(n_383), .B2(n_392), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_27), .A2(n_167), .B1(n_431), .B2(n_482), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_28), .A2(n_232), .B1(n_434), .B2(n_764), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_29), .A2(n_268), .B1(n_564), .B2(n_565), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_30), .A2(n_72), .B1(n_503), .B2(n_505), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_32), .A2(n_115), .B1(n_753), .B2(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g450 ( .A(n_33), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_34), .A2(n_141), .B1(n_336), .B2(n_763), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_35), .A2(n_116), .B1(n_832), .B2(n_836), .Y(n_831) );
INVx1_ASAP7_75t_L g912 ( .A(n_36), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_37), .A2(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g327 ( .A(n_38), .Y(n_327) );
INVxp67_ASAP7_75t_L g391 ( .A(n_38), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_38), .B(n_224), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_39), .A2(n_234), .B1(n_406), .B2(n_641), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_40), .A2(n_79), .B1(n_336), .B2(n_567), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_41), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_42), .A2(n_100), .B1(n_413), .B2(n_416), .Y(n_412) );
AOI21xp33_ASAP7_75t_SL g465 ( .A1(n_43), .A2(n_439), .B(n_466), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_44), .A2(n_124), .B1(n_839), .B2(n_843), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_45), .A2(n_278), .B1(n_847), .B2(n_868), .Y(n_913) );
AO22x1_ASAP7_75t_L g516 ( .A1(n_46), .A2(n_158), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_47), .A2(n_78), .B1(n_500), .B2(n_508), .C(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_48), .B(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_49), .A2(n_97), .B1(n_404), .B2(n_409), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g323 ( .A(n_51), .B(n_312), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_52), .A2(n_179), .B1(n_673), .B2(n_753), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_53), .A2(n_285), .B1(n_443), .B2(n_473), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_54), .A2(n_245), .B1(n_506), .B2(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_SL g582 ( .A(n_55), .Y(n_582) );
OAI21x1_ASAP7_75t_L g529 ( .A1(n_56), .A2(n_530), .B(n_547), .Y(n_529) );
NAND4xp25_ASAP7_75t_L g547 ( .A(n_56), .B(n_531), .C(n_535), .D(n_543), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_57), .A2(n_82), .B1(n_801), .B2(n_802), .C(n_803), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_58), .A2(n_204), .B1(n_305), .B2(n_331), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_59), .A2(n_269), .B1(n_447), .B2(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g1072 ( .A(n_60), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_61), .A2(n_225), .B1(n_410), .B2(n_587), .Y(n_668) );
NAND2xp33_ASAP7_75t_L g710 ( .A(n_62), .B(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_63), .A2(n_202), .B1(n_356), .B2(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_64), .A2(n_133), .B1(n_857), .B2(n_858), .Y(n_918) );
INVx1_ASAP7_75t_L g585 ( .A(n_65), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_66), .A2(n_262), .B1(n_523), .B2(n_524), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_67), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g823 ( .A(n_68), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_69), .A2(n_138), .B1(n_434), .B2(n_1061), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_70), .A2(n_233), .B1(n_443), .B2(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_71), .A2(n_194), .B1(n_673), .B2(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g736 ( .A(n_73), .Y(n_736) );
INVx1_ASAP7_75t_L g620 ( .A(n_74), .Y(n_620) );
INVx1_ASAP7_75t_SL g835 ( .A(n_75), .Y(n_835) );
AND2x4_ASAP7_75t_L g837 ( .A(n_75), .B(n_823), .Y(n_837) );
INVx1_ASAP7_75t_L g841 ( .A(n_75), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_76), .A2(n_218), .B1(n_515), .B2(n_521), .Y(n_1094) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_77), .A2(n_81), .B1(n_431), .B2(n_432), .Y(n_810) );
XNOR2x1_ASAP7_75t_L g687 ( .A(n_80), .B(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_83), .A2(n_173), .B1(n_363), .B2(n_545), .Y(n_544) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_84), .Y(n_312) );
XOR2x2_ASAP7_75t_L g552 ( .A(n_85), .B(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_86), .A2(n_205), .B1(n_505), .B2(n_506), .Y(n_542) );
INVx1_ASAP7_75t_L g723 ( .A(n_87), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_88), .A2(n_215), .B1(n_502), .B2(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_89), .B(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_90), .A2(n_176), .B1(n_839), .B2(n_843), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_91), .A2(n_198), .B1(n_502), .B2(n_503), .Y(n_541) );
INVx1_ASAP7_75t_L g579 ( .A(n_92), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_93), .A2(n_280), .B1(n_514), .B2(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g865 ( .A(n_94), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_95), .A2(n_259), .B1(n_369), .B2(n_373), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_96), .B(n_503), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_98), .A2(n_109), .B1(n_783), .B2(n_784), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_99), .A2(n_290), .B1(n_832), .B2(n_836), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_101), .A2(n_241), .B1(n_545), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_102), .A2(n_265), .B1(n_646), .B2(n_807), .Y(n_1069) );
INVx1_ASAP7_75t_L g313 ( .A(n_103), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_103), .B(n_223), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_104), .A2(n_190), .B1(n_518), .B2(n_520), .Y(n_1096) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_105), .A2(n_117), .B1(n_832), .B2(n_836), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_106), .A2(n_180), .B1(n_490), .B2(n_671), .Y(n_701) );
INVx1_ASAP7_75t_L g538 ( .A(n_107), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_108), .A2(n_113), .B1(n_434), .B2(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_110), .A2(n_135), .B1(n_771), .B2(n_772), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_112), .A2(n_174), .B1(n_363), .B2(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g741 ( .A(n_114), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_118), .A2(n_247), .B1(n_431), .B2(n_432), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_119), .A2(n_214), .B1(n_431), .B2(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g510 ( .A(n_120), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_123), .A2(n_203), .B1(n_520), .B2(n_521), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g774 ( .A1(n_126), .A2(n_159), .B1(n_592), .B2(n_775), .C(n_777), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g791 ( .A1(n_126), .A2(n_159), .B1(n_592), .B2(n_775), .C(n_777), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_127), .A2(n_231), .B1(n_839), .B2(n_847), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_128), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_129), .A2(n_216), .B1(n_342), .B2(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g664 ( .A(n_130), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_131), .A2(n_193), .B1(n_514), .B2(n_517), .Y(n_1095) );
INVxp33_ASAP7_75t_SL g871 ( .A(n_132), .Y(n_871) );
INVx1_ASAP7_75t_L g649 ( .A(n_134), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_136), .A2(n_144), .B1(n_368), .B2(n_372), .Y(n_367) );
XNOR2x1_ASAP7_75t_L g630 ( .A(n_137), .B(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_139), .A2(n_200), .B1(n_331), .B2(n_431), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_140), .A2(n_267), .B1(n_410), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_142), .A2(n_178), .B1(n_854), .B2(n_855), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_143), .A2(n_286), .B1(n_434), .B2(n_567), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_145), .A2(n_154), .B1(n_481), .B2(n_482), .Y(n_480) );
AO22x1_ASAP7_75t_L g519 ( .A1(n_146), .A2(n_284), .B1(n_520), .B2(n_521), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_147), .A2(n_210), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g448 ( .A(n_148), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_149), .A2(n_164), .B1(n_305), .B2(n_330), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_150), .A2(n_228), .B1(n_517), .B2(n_518), .Y(n_717) );
INVx1_ASAP7_75t_L g561 ( .A(n_151), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_152), .A2(n_249), .B1(n_427), .B2(n_634), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_153), .A2(n_254), .B1(n_812), .B2(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g617 ( .A(n_156), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_160), .A2(n_291), .B1(n_404), .B2(n_409), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_161), .A2(n_165), .B1(n_476), .B2(n_478), .Y(n_475) );
INVx1_ASAP7_75t_L g557 ( .A(n_162), .Y(n_557) );
AOI21xp33_ASAP7_75t_SL g577 ( .A1(n_163), .A2(n_439), .B(n_578), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_168), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_169), .A2(n_185), .B1(n_514), .B2(n_515), .Y(n_716) );
INVx1_ASAP7_75t_L g869 ( .A(n_170), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_171), .A2(n_283), .B1(n_427), .B2(n_634), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_172), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g1090 ( .A(n_175), .Y(n_1090) );
INVx1_ASAP7_75t_L g746 ( .A(n_177), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g1073 ( .A(n_178), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_178), .A2(n_1079), .B1(n_1099), .B2(n_1101), .Y(n_1078) );
XNOR2x2_ASAP7_75t_L g496 ( .A(n_181), .B(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g1056 ( .A1(n_183), .A2(n_244), .B1(n_490), .B2(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g735 ( .A(n_184), .Y(n_735) );
INVx1_ASAP7_75t_L g613 ( .A(n_186), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_187), .A2(n_264), .B1(n_342), .B2(n_434), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_188), .A2(n_239), .B1(n_646), .B2(n_647), .C(n_648), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_191), .A2(n_260), .B1(n_383), .B2(n_455), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_192), .A2(n_273), .B1(n_517), .B2(n_518), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_195), .B(n_455), .Y(n_695) );
OA22x2_ASAP7_75t_L g318 ( .A1(n_196), .A2(n_224), .B1(n_312), .B2(n_316), .Y(n_318) );
INVx1_ASAP7_75t_L g349 ( .A(n_196), .Y(n_349) );
INVx1_ASAP7_75t_L g445 ( .A(n_197), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_199), .B(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_201), .A2(n_272), .B1(n_336), .B2(n_342), .Y(n_335) );
INVx1_ASAP7_75t_L g570 ( .A(n_206), .Y(n_570) );
AOI21xp5_ASAP7_75t_SL g611 ( .A1(n_207), .A2(n_508), .B(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_208), .A2(n_226), .B1(n_523), .B2(n_524), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_209), .A2(n_221), .B1(n_564), .B2(n_565), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_212), .A2(n_287), .B1(n_854), .B2(n_855), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_213), .A2(n_271), .B1(n_305), .B2(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g467 ( .A(n_217), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_219), .A2(n_253), .B1(n_429), .B2(n_490), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_220), .A2(n_275), .B1(n_410), .B2(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_222), .B(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g329 ( .A(n_223), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_223), .B(n_347), .Y(n_401) );
OAI21xp33_ASAP7_75t_L g350 ( .A1(n_224), .A2(n_248), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g609 ( .A(n_227), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_229), .A2(n_274), .B1(n_514), .B2(n_515), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_230), .A2(n_243), .B1(n_523), .B2(n_524), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_231), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g882 ( .A1(n_235), .A2(n_258), .B1(n_832), .B2(n_836), .Y(n_882) );
INVx1_ASAP7_75t_L g911 ( .A(n_236), .Y(n_911) );
INVx1_ASAP7_75t_L g458 ( .A(n_238), .Y(n_458) );
INVx1_ASAP7_75t_SL g589 ( .A(n_240), .Y(n_589) );
INVxp67_ASAP7_75t_SL g779 ( .A(n_242), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_246), .A2(n_293), .B1(n_520), .B2(n_521), .Y(n_720) );
INVx1_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_248), .B(n_281), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g693 ( .A(n_250), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_251), .B(n_1067), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_252), .A2(n_296), .B1(n_369), .B2(n_429), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_255), .A2(n_266), .B1(n_587), .B2(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g743 ( .A(n_256), .Y(n_743) );
INVx1_ASAP7_75t_SL g569 ( .A(n_263), .Y(n_569) );
AOI21xp33_ASAP7_75t_L g1088 ( .A1(n_270), .A2(n_505), .B(n_1089), .Y(n_1088) );
AOI21xp33_ASAP7_75t_SL g721 ( .A1(n_276), .A2(n_508), .B(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_278), .Y(n_419) );
INVx1_ASAP7_75t_L g778 ( .A(n_279), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_281), .B(n_322), .Y(n_321) );
XNOR2x1_ASAP7_75t_L g731 ( .A(n_282), .B(n_732), .Y(n_731) );
INVxp33_ASAP7_75t_L g863 ( .A(n_288), .Y(n_863) );
INVx1_ASAP7_75t_L g834 ( .A(n_289), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_292), .Y(n_804) );
INVx1_ASAP7_75t_L g441 ( .A(n_294), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_295), .A2(n_1080), .B1(n_1081), .B2(n_1098), .Y(n_1079) );
CKINVDCx5p33_ASAP7_75t_R g1080 ( .A(n_295), .Y(n_1080) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_625), .B(n_817), .C(n_826), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_298), .A2(n_625), .B(n_818), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B1(n_492), .B2(n_493), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
XNOR2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_422), .Y(n_300) );
AO211x2_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_365), .B(n_420), .C(n_421), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_352), .Y(n_302) );
AO22x2_ASAP7_75t_L g421 ( .A1(n_303), .A2(n_366), .B1(n_419), .B2(n_1106), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_304), .B(n_335), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_306), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
INVx2_ASAP7_75t_L g757 ( .A(n_306), .Y(n_757) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx12f_ASAP7_75t_L g431 ( .A(n_307), .Y(n_431) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_307), .Y(n_481) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_319), .Y(n_307) );
AND2x2_ASAP7_75t_L g332 ( .A(n_308), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g357 ( .A(n_308), .B(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g364 ( .A(n_308), .B(n_339), .Y(n_364) );
AND2x4_ASAP7_75t_L g520 ( .A(n_308), .B(n_339), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_308), .B(n_371), .Y(n_521) );
AND2x4_ASAP7_75t_L g523 ( .A(n_308), .B(n_319), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_308), .B(n_333), .Y(n_524) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_317), .Y(n_308) );
AND2x2_ASAP7_75t_L g408 ( .A(n_309), .B(n_318), .Y(n_408) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g338 ( .A(n_310), .B(n_318), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
NAND2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx2_ASAP7_75t_L g316 ( .A(n_312), .Y(n_316) );
INVx3_ASAP7_75t_L g322 ( .A(n_312), .Y(n_322) );
NAND2xp33_ASAP7_75t_L g328 ( .A(n_312), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g351 ( .A(n_312), .Y(n_351) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_312), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_313), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
OAI21xp5_ASAP7_75t_L g390 ( .A1(n_315), .A2(n_351), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g389 ( .A(n_318), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g407 ( .A(n_319), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g411 ( .A(n_319), .B(n_338), .Y(n_411) );
AND2x4_ASAP7_75t_L g502 ( .A(n_319), .B(n_338), .Y(n_502) );
AND2x4_ASAP7_75t_L g505 ( .A(n_319), .B(n_408), .Y(n_505) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .Y(n_319) );
INVx2_ASAP7_75t_L g334 ( .A(n_320), .Y(n_334) );
AND2x4_ASAP7_75t_L g339 ( .A(n_320), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g359 ( .A(n_320), .B(n_341), .Y(n_359) );
AND2x2_ASAP7_75t_L g385 ( .A(n_320), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_322), .B(n_327), .Y(n_326) );
INVxp67_ASAP7_75t_L g347 ( .A(n_322), .Y(n_347) );
NAND3xp33_ASAP7_75t_L g400 ( .A(n_323), .B(n_346), .C(n_401), .Y(n_400) );
AND2x4_ASAP7_75t_L g333 ( .A(n_324), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g341 ( .A(n_325), .Y(n_341) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_332), .Y(n_432) );
BUFx5_ASAP7_75t_L g482 ( .A(n_332), .Y(n_482) );
INVx1_ASAP7_75t_L g761 ( .A(n_332), .Y(n_761) );
AND2x2_ASAP7_75t_L g381 ( .A(n_333), .B(n_338), .Y(n_381) );
AND2x4_ASAP7_75t_L g415 ( .A(n_333), .B(n_408), .Y(n_415) );
AND2x4_ASAP7_75t_L g418 ( .A(n_333), .B(n_345), .Y(n_418) );
AND2x2_ASAP7_75t_L g500 ( .A(n_333), .B(n_338), .Y(n_500) );
AND2x4_ASAP7_75t_L g506 ( .A(n_333), .B(n_345), .Y(n_506) );
AND2x2_ASAP7_75t_L g508 ( .A(n_333), .B(n_408), .Y(n_508) );
BUFx8_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_337), .Y(n_434) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
AND2x4_ASAP7_75t_L g370 ( .A(n_338), .B(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g514 ( .A(n_338), .B(n_358), .Y(n_514) );
AND2x4_ASAP7_75t_L g517 ( .A(n_338), .B(n_339), .Y(n_517) );
AND2x2_ASAP7_75t_L g674 ( .A(n_338), .B(n_339), .Y(n_674) );
AND2x4_ASAP7_75t_L g344 ( .A(n_339), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g518 ( .A(n_339), .B(n_345), .Y(n_518) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx4_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g484 ( .A(n_343), .Y(n_484) );
INVx4_ASAP7_75t_L g567 ( .A(n_343), .Y(n_567) );
INVx1_ASAP7_75t_L g677 ( .A(n_343), .Y(n_677) );
INVx4_ASAP7_75t_L g764 ( .A(n_343), .Y(n_764) );
INVx1_ASAP7_75t_L g1061 ( .A(n_343), .Y(n_1061) );
INVx8_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g375 ( .A(n_345), .B(n_358), .Y(n_375) );
AND2x4_ASAP7_75t_L g515 ( .A(n_345), .B(n_358), .Y(n_515) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_350), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AO22x1_ASAP7_75t_L g420 ( .A1(n_352), .A2(n_402), .B1(n_419), .B2(n_1105), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_360), .B2(n_361), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_357), .Y(n_488) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_357), .Y(n_545) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_357), .Y(n_634) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g371 ( .A(n_359), .Y(n_371) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx12f_ASAP7_75t_L g564 ( .A(n_363), .Y(n_564) );
BUFx12f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_364), .Y(n_427) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_364), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_402), .C(n_419), .Y(n_365) );
NAND2x1_ASAP7_75t_L g366 ( .A(n_367), .B(n_376), .Y(n_366) );
INVx1_ASAP7_75t_L g556 ( .A(n_368), .Y(n_556) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_370), .Y(n_490) );
BUFx12f_ASAP7_75t_L g675 ( .A(n_370), .Y(n_675) );
BUFx6f_ASAP7_75t_L g812 ( .A(n_370), .Y(n_812) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g560 ( .A(n_373), .Y(n_560) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx3_ASAP7_75t_L g534 ( .A(n_374), .Y(n_534) );
INVx5_ASAP7_75t_L g671 ( .A(n_374), .Y(n_671) );
INVx2_ASAP7_75t_L g813 ( .A(n_374), .Y(n_813) );
INVx1_ASAP7_75t_L g1057 ( .A(n_374), .Y(n_1057) );
INVx6_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx12f_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
OA21x2_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_382), .Y(n_376) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g453 ( .A(n_381), .Y(n_453) );
INVx2_ASAP7_75t_L g464 ( .A(n_381), .Y(n_464) );
BUFx4f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx5_ASAP7_75t_L g474 ( .A(n_384), .Y(n_474) );
BUFx2_ASAP7_75t_L g660 ( .A(n_384), .Y(n_660) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_389), .Y(n_384) );
AND2x4_ASAP7_75t_L g503 ( .A(n_385), .B(n_389), .Y(n_503) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_385), .B(n_389), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g396 ( .A(n_387), .Y(n_396) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx4_ASAP7_75t_L g455 ( .A(n_393), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_393), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g1089 ( .A(n_393), .B(n_1090), .Y(n_1089) );
INVx4_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx3_ASAP7_75t_L g539 ( .A(n_394), .Y(n_539) );
INVx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_395), .Y(n_470) );
AO21x2_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_400), .Y(n_395) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_397), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_412), .Y(n_402) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_405), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_734) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g440 ( .A(n_407), .Y(n_440) );
BUFx3_ASAP7_75t_L g659 ( .A(n_407), .Y(n_659) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_407), .Y(n_801) );
BUFx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g590 ( .A(n_410), .Y(n_590) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx3_ASAP7_75t_L g443 ( .A(n_411), .Y(n_443) );
INVx2_ASAP7_75t_L g644 ( .A(n_411), .Y(n_644) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx3_ASAP7_75t_L g584 ( .A(n_414), .Y(n_584) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g447 ( .A(n_415), .Y(n_447) );
INVx2_ASAP7_75t_L g477 ( .A(n_415), .Y(n_477) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_415), .Y(n_662) );
BUFx6f_ASAP7_75t_L g1085 ( .A(n_415), .Y(n_1085) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_417), .A2(n_445), .B1(n_446), .B2(n_448), .Y(n_444) );
INVx3_ASAP7_75t_L g697 ( .A(n_417), .Y(n_697) );
INVx2_ASAP7_75t_L g807 ( .A(n_417), .Y(n_807) );
INVx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_418), .Y(n_478) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_418), .Y(n_587) );
AOI22x1_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_456), .B1(n_457), .B2(n_491), .Y(n_422) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_435), .Y(n_424) );
AND4x1_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .C(n_430), .D(n_433), .Y(n_425) );
BUFx3_ASAP7_75t_L g784 ( .A(n_429), .Y(n_784) );
INVx1_ASAP7_75t_L g571 ( .A(n_432), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_444), .C(n_449), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_441), .B2(n_442), .Y(n_436) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g699 ( .A(n_440), .Y(n_699) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B(n_454), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g776 ( .A(n_453), .Y(n_776) );
INVx2_ASAP7_75t_L g802 ( .A(n_453), .Y(n_802) );
INVx3_ASAP7_75t_SL g1067 ( .A(n_453), .Y(n_1067) );
INVx2_ASAP7_75t_L g1092 ( .A(n_453), .Y(n_1092) );
INVx2_ASAP7_75t_L g580 ( .A(n_455), .Y(n_580) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
XNOR2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
NOR4xp75_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .C(n_479), .D(n_485), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .Y(n_460) );
INVx1_ASAP7_75t_L g747 ( .A(n_462), .Y(n_747) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g667 ( .A(n_463), .Y(n_667) );
INVx2_ASAP7_75t_L g691 ( .A(n_463), .Y(n_691) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g576 ( .A(n_464), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_470), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_SL g651 ( .A(n_470), .Y(n_651) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_470), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g592 ( .A(n_474), .Y(n_592) );
INVx4_ASAP7_75t_L g641 ( .A(n_474), .Y(n_641) );
INVx3_ASAP7_75t_L g749 ( .A(n_474), .Y(n_749) );
INVx2_ASAP7_75t_L g1065 ( .A(n_474), .Y(n_1065) );
INVx2_ASAP7_75t_L g742 ( .A(n_476), .Y(n_742) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_SL g646 ( .A(n_477), .Y(n_646) );
INVx4_ASAP7_75t_L g744 ( .A(n_478), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_480), .B(n_483), .Y(n_479) );
BUFx3_ASAP7_75t_L g788 ( .A(n_482), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_486), .B(n_489), .Y(n_485) );
BUFx3_ASAP7_75t_L g565 ( .A(n_488), .Y(n_565) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
XOR2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_550), .Y(n_493) );
AO22x2_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_525), .B1(n_548), .B2(n_549), .Y(n_494) );
INVx2_ASAP7_75t_L g548 ( .A(n_495), .Y(n_548) );
BUFx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_511), .Y(n_497) );
AND4x1_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .C(n_504), .D(n_507), .Y(n_498) );
INVx2_ASAP7_75t_L g610 ( .A(n_500), .Y(n_610) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_500), .Y(n_711) );
INVx1_ASAP7_75t_L g621 ( .A(n_502), .Y(n_621) );
INVx4_ASAP7_75t_L g694 ( .A(n_503), .Y(n_694) );
INVx2_ASAP7_75t_L g616 ( .A(n_505), .Y(n_616) );
INVx2_ASAP7_75t_L g618 ( .A(n_506), .Y(n_618) );
NOR4xp25_ASAP7_75t_L g511 ( .A(n_512), .B(n_516), .C(n_519), .D(n_522), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g549 ( .A(n_527), .Y(n_549) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND3x1_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .C(n_543), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_540), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx4_ASAP7_75t_L g750 ( .A(n_539), .Y(n_750) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_593), .B1(n_623), .B2(n_624), .Y(n_550) );
INVx2_ASAP7_75t_L g623 ( .A(n_551), .Y(n_623) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_572), .Y(n_553) );
NOR3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_562), .C(n_568), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_558), .B2(n_561), .Y(n_555) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g754 ( .A(n_560), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_563), .B(n_566), .Y(n_562) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_581), .C(n_588), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_574), .B(n_577), .Y(n_573) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B1(n_585), .B2(n_586), .Y(n_581) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx3_ASAP7_75t_L g772 ( .A(n_587), .Y(n_772) );
OAI21xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g624 ( .A(n_595), .Y(n_624) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OA22x2_ASAP7_75t_L g795 ( .A1(n_596), .A2(n_796), .B1(n_815), .B2(n_816), .Y(n_795) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
XNOR2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
XNOR2xp5_ASAP7_75t_L g816 ( .A(n_598), .B(n_599), .Y(n_816) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_607), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_614), .C(n_619), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_611), .Y(n_608) );
INVx2_ASAP7_75t_L g647 ( .A(n_610), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B1(n_617), .B2(n_618), .Y(n_614) );
INVxp67_ASAP7_75t_L g713 ( .A(n_618), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g619 ( .A1(n_620), .A2(n_621), .B(n_622), .Y(n_619) );
XNOR2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_728), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_685), .B1(n_726), .B2(n_727), .Y(n_626) );
INVx2_ASAP7_75t_L g726 ( .A(n_627), .Y(n_726) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
XNOR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_652), .Y(n_629) );
NAND4xp75_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .C(n_639), .D(n_645), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
BUFx3_ASAP7_75t_L g783 ( .A(n_634), .Y(n_783) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx6f_ASAP7_75t_L g739 ( .A(n_644), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NOR2xp33_ASAP7_75t_R g777 ( .A(n_650), .B(n_778), .Y(n_777) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
OAI21x1_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B(n_679), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_653), .B(n_668), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_654), .Y(n_653) );
NOR2xp67_ASAP7_75t_L g655 ( .A(n_656), .B(n_669), .Y(n_655) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_666), .C(n_668), .Y(n_656) );
INVx1_ASAP7_75t_L g683 ( .A(n_657), .Y(n_683) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_661), .Y(n_657) );
BUFx3_ASAP7_75t_L g771 ( .A(n_662), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_665), .B(n_723), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_665), .B(n_804), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g1071 ( .A(n_665), .B(n_1072), .Y(n_1071) );
INVxp67_ASAP7_75t_L g681 ( .A(n_666), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_669), .Y(n_684) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .C(n_676), .D(n_678), .Y(n_669) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx3_ASAP7_75t_L g753 ( .A(n_675), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_684), .Y(n_679) );
NOR3xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .C(n_683), .Y(n_680) );
INVx1_ASAP7_75t_L g727 ( .A(n_685), .Y(n_727) );
BUFx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OA22x2_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_705), .B1(n_724), .B2(n_725), .Y(n_686) );
INVx1_ASAP7_75t_L g725 ( .A(n_687), .Y(n_725) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_700), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_696), .C(n_698), .Y(n_689) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B(n_695), .Y(n_692) );
NAND4xp25_ASAP7_75t_SL g700 ( .A(n_701), .B(n_702), .C(n_703), .D(n_704), .Y(n_700) );
INVx3_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_706), .Y(n_724) );
XNOR2x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
NOR2x1_ASAP7_75t_L g708 ( .A(n_709), .B(n_715), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .C(n_714), .Y(n_709) );
NAND4xp25_ASAP7_75t_SL g715 ( .A(n_716), .B(n_717), .C(n_718), .D(n_721), .Y(n_715) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
XOR2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_794), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_765), .B1(n_792), .B2(n_793), .Y(n_729) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g792 ( .A(n_731), .Y(n_792) );
AND2x4_ASAP7_75t_L g732 ( .A(n_733), .B(n_751), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_740), .C(n_745), .Y(n_733) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B1(n_743), .B2(n_744), .Y(n_740) );
OAI21xp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B(n_748), .Y(n_745) );
AND4x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_755), .C(n_756), .D(n_762), .Y(n_751) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
BUFx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_SL g793 ( .A(n_765), .Y(n_793) );
AO22x2_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_779), .B1(n_780), .B2(n_790), .Y(n_765) );
NOR3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_773), .C(n_779), .Y(n_766) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND4xp75_ASAP7_75t_SL g790 ( .A(n_768), .B(n_781), .C(n_786), .D(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AND2x2_ASAP7_75t_L g780 ( .A(n_781), .B(n_786), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .Y(n_781) );
AND2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_789), .Y(n_786) );
BUFx2_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
INVxp67_ASAP7_75t_SL g815 ( .A(n_796), .Y(n_815) );
XNOR2x1_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
OR2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_808), .Y(n_798) );
NAND3xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_805), .C(n_806), .Y(n_799) );
NAND4xp25_ASAP7_75t_SL g808 ( .A(n_809), .B(n_810), .C(n_811), .D(n_814), .Y(n_808) );
BUFx10_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_824), .C(n_825), .Y(n_820) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_821), .B(n_1076), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_821), .B(n_1077), .Y(n_1100) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
OA21x2_ASAP7_75t_L g1102 ( .A1(n_822), .A2(n_835), .B(n_1103), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AND3x4_ASAP7_75t_L g832 ( .A(n_823), .B(n_833), .C(n_835), .Y(n_832) );
AND2x2_ASAP7_75t_L g840 ( .A(n_823), .B(n_841), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g1076 ( .A(n_824), .B(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_825), .Y(n_1077) );
OAI221xp5_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_1050), .B1(n_1052), .B2(n_1074), .C(n_1078), .Y(n_826) );
AOI211x1_ASAP7_75t_SL g827 ( .A1(n_828), .A2(n_906), .B(n_920), .C(n_1028), .Y(n_827) );
OAI211xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_849), .B(n_875), .C(n_895), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_844), .Y(n_829) );
INVx1_ASAP7_75t_L g880 ( .A(n_830), .Y(n_880) );
OR2x2_ASAP7_75t_L g898 ( .A(n_830), .B(n_881), .Y(n_898) );
AND2x2_ASAP7_75t_L g937 ( .A(n_830), .B(n_881), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_830), .B(n_845), .Y(n_956) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_838), .Y(n_830) );
AND2x4_ASAP7_75t_L g836 ( .A(n_833), .B(n_837), .Y(n_836) );
AND2x4_ASAP7_75t_L g854 ( .A(n_833), .B(n_840), .Y(n_854) );
AND2x4_ASAP7_75t_L g855 ( .A(n_833), .B(n_837), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_833), .B(n_837), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g1103 ( .A(n_833), .Y(n_1103) );
AND2x2_ASAP7_75t_L g843 ( .A(n_837), .B(n_842), .Y(n_843) );
AND2x4_ASAP7_75t_L g847 ( .A(n_837), .B(n_842), .Y(n_847) );
AND2x2_ASAP7_75t_L g858 ( .A(n_837), .B(n_842), .Y(n_858) );
AND2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_842), .Y(n_839) );
AND2x2_ASAP7_75t_L g857 ( .A(n_840), .B(n_842), .Y(n_857) );
AND2x4_ASAP7_75t_L g868 ( .A(n_840), .B(n_842), .Y(n_868) );
NOR2x1_ASAP7_75t_R g892 ( .A(n_844), .B(n_893), .Y(n_892) );
AND2x2_ASAP7_75t_L g933 ( .A(n_844), .B(n_879), .Y(n_933) );
AND2x2_ASAP7_75t_L g951 ( .A(n_844), .B(n_880), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_844), .B(n_985), .Y(n_984) );
AND2x2_ASAP7_75t_L g998 ( .A(n_844), .B(n_937), .Y(n_998) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_844), .B(n_989), .Y(n_1025) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_SL g878 ( .A(n_845), .Y(n_878) );
AND2x2_ASAP7_75t_L g889 ( .A(n_845), .B(n_890), .Y(n_889) );
OR2x2_ASAP7_75t_L g926 ( .A(n_845), .B(n_891), .Y(n_926) );
AND2x2_ASAP7_75t_L g988 ( .A(n_845), .B(n_989), .Y(n_988) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_845), .B(n_898), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_845), .B(n_880), .Y(n_1030) );
AND2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_848), .Y(n_845) );
INVx2_ASAP7_75t_L g870 ( .A(n_847), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_859), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_850), .B(n_951), .Y(n_950) );
NAND2xp67_ASAP7_75t_L g1048 ( .A(n_850), .B(n_876), .Y(n_1048) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NOR2x1_ASAP7_75t_L g890 ( .A(n_851), .B(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_SL g893 ( .A(n_851), .B(n_894), .Y(n_893) );
BUFx6f_ASAP7_75t_L g904 ( .A(n_851), .Y(n_904) );
INVx2_ASAP7_75t_L g925 ( .A(n_851), .Y(n_925) );
INVx1_ASAP7_75t_L g939 ( .A(n_851), .Y(n_939) );
AND2x2_ASAP7_75t_L g981 ( .A(n_851), .B(n_860), .Y(n_981) );
AND2x2_ASAP7_75t_L g987 ( .A(n_851), .B(n_988), .Y(n_987) );
NOR2xp33_ASAP7_75t_L g993 ( .A(n_851), .B(n_930), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_851), .B(n_951), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_851), .B(n_928), .Y(n_1016) );
INVx4_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_852), .B(n_887), .Y(n_957) );
OR2x2_ASAP7_75t_L g961 ( .A(n_852), .B(n_877), .Y(n_961) );
AND2x2_ASAP7_75t_L g976 ( .A(n_852), .B(n_860), .Y(n_976) );
AND2x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_856), .Y(n_852) );
INVx3_ASAP7_75t_L g862 ( .A(n_854), .Y(n_862) );
INVx1_ASAP7_75t_L g963 ( .A(n_859), .Y(n_963) );
AND2x2_ASAP7_75t_L g859 ( .A(n_860), .B(n_872), .Y(n_859) );
INVx2_ASAP7_75t_L g887 ( .A(n_860), .Y(n_887) );
INVx1_ASAP7_75t_L g928 ( .A(n_860), .Y(n_928) );
OR2x2_ASAP7_75t_L g970 ( .A(n_860), .B(n_872), .Y(n_970) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_860), .B(n_977), .Y(n_1022) );
OR2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_866), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_861) );
OAI221xp5_ASAP7_75t_L g910 ( .A1(n_862), .A2(n_864), .B1(n_911), .B2(n_912), .C(n_913), .Y(n_910) );
BUFx2_ASAP7_75t_L g1051 ( .A(n_864), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_869), .B1(n_870), .B2(n_871), .Y(n_866) );
INVx3_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
OR2x2_ASAP7_75t_L g900 ( .A(n_872), .B(n_887), .Y(n_900) );
AND2x2_ASAP7_75t_L g905 ( .A(n_872), .B(n_887), .Y(n_905) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_872), .Y(n_940) );
OR2x2_ASAP7_75t_L g944 ( .A(n_872), .B(n_916), .Y(n_944) );
AND2x2_ASAP7_75t_L g953 ( .A(n_872), .B(n_915), .Y(n_953) );
OR2x2_ASAP7_75t_L g972 ( .A(n_872), .B(n_917), .Y(n_972) );
AND2x2_ASAP7_75t_L g977 ( .A(n_872), .B(n_916), .Y(n_977) );
INVx2_ASAP7_75t_L g1004 ( .A(n_872), .Y(n_1004) );
AND2x2_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_884), .B1(n_885), .B2(n_892), .Y(n_875) );
INVx1_ASAP7_75t_L g962 ( .A(n_876), .Y(n_962) );
AND2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_879), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g895 ( .A1(n_877), .A2(n_896), .B1(n_899), .B2(n_901), .Y(n_895) );
AND2x4_ASAP7_75t_L g896 ( .A(n_877), .B(n_897), .Y(n_896) );
AND2x2_ASAP7_75t_L g936 ( .A(n_877), .B(n_937), .Y(n_936) );
AND2x2_ASAP7_75t_L g949 ( .A(n_877), .B(n_881), .Y(n_949) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
AOI211xp5_ASAP7_75t_L g945 ( .A1(n_879), .A2(n_946), .B(n_947), .C(n_958), .Y(n_945) );
INVx1_ASAP7_75t_L g1013 ( .A(n_879), .Y(n_1013) );
AND2x2_ASAP7_75t_L g879 ( .A(n_880), .B(n_881), .Y(n_879) );
OR2x2_ASAP7_75t_L g891 ( .A(n_880), .B(n_881), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_880), .B(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g989 ( .A(n_881), .Y(n_989) );
AOI222xp33_ASAP7_75t_L g1037 ( .A1(n_881), .A2(n_905), .B1(n_1038), .B2(n_1039), .C1(n_1041), .C2(n_1042), .Y(n_1037) );
AND2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_888), .Y(n_884) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_885), .B(n_932), .Y(n_931) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g942 ( .A(n_886), .B(n_943), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_886), .B(n_949), .Y(n_948) );
A2O1A1Ixp33_ASAP7_75t_L g1045 ( .A1(n_886), .A2(n_1046), .B(n_1047), .C(n_1049), .Y(n_1045) );
NOR2xp67_ASAP7_75t_SL g1047 ( .A(n_886), .B(n_1048), .Y(n_1047) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_887), .B(n_930), .Y(n_1000) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx3_ASAP7_75t_SL g894 ( .A(n_891), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_894), .B(n_960), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1029 ( .A1(n_894), .A2(n_946), .B1(n_1030), .B2(n_1031), .C(n_1032), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_896), .B(n_924), .Y(n_923) );
INVx2_ASAP7_75t_SL g943 ( .A(n_896), .Y(n_943) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_896), .B(n_925), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_897), .B(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_898), .B(n_979), .Y(n_985) );
AND2x2_ASAP7_75t_L g946 ( .A(n_899), .B(n_929), .Y(n_946) );
AOI321xp33_ASAP7_75t_L g992 ( .A1(n_899), .A2(n_993), .A3(n_994), .B1(n_995), .B2(n_997), .C(n_999), .Y(n_992) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .Y(n_902) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_903), .B(n_998), .Y(n_1021) );
INVx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
OAI221xp5_ASAP7_75t_L g965 ( .A1(n_904), .A2(n_966), .B1(n_971), .B2(n_972), .C(n_973), .Y(n_965) );
OAI321xp33_ASAP7_75t_L g983 ( .A1(n_904), .A2(n_972), .A3(n_984), .B1(n_986), .B2(n_990), .C(n_992), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_904), .B(n_905), .Y(n_1043) );
AND2x2_ASAP7_75t_L g997 ( .A(n_905), .B(n_998), .Y(n_997) );
INVxp67_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_908), .B(n_914), .Y(n_907) );
OAI31xp33_ASAP7_75t_L g921 ( .A1(n_908), .A2(n_922), .A3(n_931), .B(n_934), .Y(n_921) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
AOI211xp5_ASAP7_75t_L g964 ( .A1(n_909), .A2(n_965), .B(n_983), .C(n_1002), .Y(n_964) );
AOI222xp33_ASAP7_75t_L g1009 ( .A1(n_909), .A2(n_953), .B1(n_1010), .B2(n_1011), .C1(n_1014), .C2(n_1019), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g996 ( .A(n_910), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_910), .B(n_929), .Y(n_1044) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g930 ( .A(n_917), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
NAND4xp25_ASAP7_75t_L g920 ( .A(n_921), .B(n_964), .C(n_1009), .D(n_1020), .Y(n_920) );
AOI21xp33_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_926), .B(n_927), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_924), .B(n_936), .Y(n_1006) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_925), .B(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g1046 ( .A(n_926), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
INVx2_ASAP7_75t_L g991 ( .A(n_928), .Y(n_991) );
OAI322xp33_ASAP7_75t_L g1032 ( .A1(n_928), .A2(n_979), .A3(n_989), .B1(n_1012), .B2(n_1033), .C1(n_1034), .C2(n_1036), .Y(n_1032) );
INVx1_ASAP7_75t_L g1019 ( .A(n_929), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_929), .B(n_1016), .Y(n_1036) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
BUFx3_ASAP7_75t_L g968 ( .A(n_930), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g1031 ( .A(n_930), .B(n_970), .Y(n_1031) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_933), .B(n_936), .Y(n_935) );
AOI321xp33_ASAP7_75t_L g1020 ( .A1(n_933), .A2(n_996), .A3(n_1004), .B1(n_1021), .B2(n_1022), .C(n_1023), .Y(n_1020) );
OAI221xp5_ASAP7_75t_SL g934 ( .A1(n_935), .A2(n_938), .B1(n_941), .B2(n_944), .C(n_945), .Y(n_934) );
INVx1_ASAP7_75t_L g971 ( .A(n_936), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_937), .B(n_960), .Y(n_959) );
INVx1_ASAP7_75t_L g979 ( .A(n_937), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g1027 ( .A(n_939), .B(n_970), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_940), .B(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g1040 ( .A(n_940), .Y(n_1040) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
O2A1O1Ixp33_ASAP7_75t_L g999 ( .A1(n_944), .A2(n_996), .B(n_1000), .C(n_1001), .Y(n_999) );
A2O1A1Ixp33_ASAP7_75t_L g947 ( .A1(n_948), .A2(n_950), .B(n_952), .C(n_954), .Y(n_947) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_953), .B(n_991), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g955 ( .A(n_956), .B(n_957), .Y(n_955) );
INVx1_ASAP7_75t_L g994 ( .A(n_956), .Y(n_994) );
AOI21xp33_ASAP7_75t_SL g958 ( .A1(n_959), .A2(n_962), .B(n_963), .Y(n_958) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
OR2x2_ASAP7_75t_L g1012 ( .A(n_961), .B(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1007 ( .A(n_967), .Y(n_1007) );
AND2x2_ASAP7_75t_L g967 ( .A(n_968), .B(n_969), .Y(n_967) );
INVx2_ASAP7_75t_L g982 ( .A(n_968), .Y(n_982) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
AOI21xp33_ASAP7_75t_L g1023 ( .A1(n_971), .A2(n_1024), .B(n_1026), .Y(n_1023) );
AOI21xp5_ASAP7_75t_L g973 ( .A1(n_974), .A2(n_977), .B(n_978), .Y(n_973) );
INVxp67_ASAP7_75t_SL g974 ( .A(n_975), .Y(n_974) );
NOR3xp33_ASAP7_75t_L g978 ( .A(n_979), .B(n_980), .C(n_982), .Y(n_978) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
NOR2xp33_ASAP7_75t_L g1010 ( .A(n_991), .B(n_1006), .Y(n_1010) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_991), .B(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1033 ( .A(n_993), .Y(n_1033) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1005 ( .A(n_996), .Y(n_1005) );
OAI221xp5_ASAP7_75t_SL g1028 ( .A1(n_996), .A2(n_1029), .B1(n_1037), .B2(n_1044), .C(n_1045), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_1003), .A2(n_1006), .B1(n_1007), .B2(n_1008), .Y(n_1002) );
INVxp67_ASAP7_75t_L g1049 ( .A(n_1003), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1005), .Y(n_1003) );
CKINVDCx14_ASAP7_75t_R g1035 ( .A(n_1004), .Y(n_1035) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1008), .Y(n_1038) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1017), .Y(n_1015) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
CKINVDCx14_ASAP7_75t_R g1034 ( .A(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
INVxp67_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
BUFx2_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
BUFx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
XNOR2x1_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1073), .Y(n_1053) );
NOR4xp75_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1059), .C(n_1063), .D(n_1068), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1058), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1062), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1066), .Y(n_1063) );
NAND2xp5_ASAP7_75t_SL g1068 ( .A(n_1069), .B(n_1070), .Y(n_1068) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1081), .Y(n_1098) );
INVxp33_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
NOR2xp33_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1093), .Y(n_1082) );
NAND4xp25_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1086), .C(n_1088), .D(n_1091), .Y(n_1083) );
NAND4xp25_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1095), .C(n_1096), .D(n_1097), .Y(n_1093) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
endmodule