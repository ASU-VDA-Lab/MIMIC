module real_jpeg_24520_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_0),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_0),
.A2(n_33),
.B1(n_38),
.B2(n_40),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_0),
.A2(n_33),
.B1(n_64),
.B2(n_69),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_0),
.A2(n_33),
.B1(n_58),
.B2(n_59),
.Y(n_353)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_2),
.A2(n_55),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_2),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_2),
.A2(n_64),
.B1(n_69),
.B2(n_73),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_2),
.A2(n_38),
.B1(n_40),
.B2(n_73),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_73),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_3),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_3),
.A2(n_64),
.B1(n_69),
.B2(n_108),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_3),
.A2(n_38),
.B1(n_40),
.B2(n_108),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_3),
.A2(n_26),
.B1(n_32),
.B2(n_108),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_4),
.A2(n_38),
.B1(n_40),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_4),
.A2(n_26),
.B1(n_32),
.B2(n_48),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_4),
.A2(n_48),
.B1(n_64),
.B2(n_69),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_4),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_344)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_7),
.A2(n_55),
.B1(n_143),
.B2(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_7),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_7),
.A2(n_64),
.B1(n_69),
.B2(n_159),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_7),
.A2(n_38),
.B1(n_40),
.B2(n_159),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_7),
.A2(n_26),
.B1(n_32),
.B2(n_159),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_9),
.B(n_63),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_9),
.B(n_38),
.C(n_82),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_9),
.A2(n_64),
.B1(n_69),
.B2(n_183),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_9),
.B(n_123),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_9),
.A2(n_38),
.B1(n_40),
.B2(n_183),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_9),
.B(n_26),
.C(n_43),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_9),
.A2(n_25),
.B(n_275),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_10),
.A2(n_64),
.B1(n_69),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_10),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_10),
.A2(n_38),
.B1(n_40),
.B2(n_86),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_86),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_10),
.A2(n_26),
.B1(n_32),
.B2(n_86),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_11),
.A2(n_37),
.B1(n_64),
.B2(n_69),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_11),
.A2(n_37),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_11),
.A2(n_26),
.B1(n_32),
.B2(n_37),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_14),
.A2(n_55),
.B1(n_58),
.B2(n_61),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_14),
.A2(n_61),
.B1(n_64),
.B2(n_69),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_14),
.A2(n_38),
.B1(n_40),
.B2(n_61),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_14),
.A2(n_26),
.B1(n_32),
.B2(n_61),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_16),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_16),
.A2(n_186),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_349),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_336),
.B(n_348),
.Y(n_18)
);

OAI31xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_133),
.A3(n_149),
.B(n_333),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_21),
.B(n_112),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_77),
.C(n_93),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_22),
.A2(n_77),
.B1(n_78),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_22),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_23),
.A2(n_24),
.B(n_52),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_24),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_31),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_25),
.A2(n_28),
.B1(n_31),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_25),
.A2(n_28),
.B1(n_98),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_25),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_25),
.A2(n_188),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_25),
.B(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_25),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_32),
.B1(n_43),
.B2(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_27),
.B(n_183),
.Y(n_300)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_30),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_32),
.B(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_36),
.A2(n_41),
.B1(n_49),
.B2(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_40),
.B1(n_43),
.B2(n_45),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_38),
.A2(n_40),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_38),
.B(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_41),
.A2(n_49),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_41),
.B(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_41),
.A2(n_49),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_46),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_46),
.A2(n_89),
.B1(n_102),
.B2(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_46),
.A2(n_169),
.B(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_46),
.A2(n_209),
.B(n_248),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_46),
.B(n_183),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_47),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_49),
.B(n_210),
.Y(n_263)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_62),
.B(n_70),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_54),
.A2(n_62),
.B1(n_109),
.B2(n_131),
.Y(n_130)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_57),
.B1(n_67),
.B2(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_56),
.B(n_183),
.Y(n_182)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_SL g184 ( 
.A(n_58),
.B(n_67),
.C(n_69),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_58),
.A2(n_182),
.B(n_183),
.Y(n_212)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_72),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_62),
.A2(n_109),
.B1(n_131),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_62),
.A2(n_70),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_63),
.A2(n_75),
.B1(n_107),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_63),
.A2(n_75),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_63),
.A2(n_75),
.B1(n_344),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_63)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_69),
.B1(n_82),
.B2(n_83),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_64),
.A2(n_68),
.B(n_182),
.C(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_64),
.B(n_238),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_75),
.A2(n_111),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_88),
.B(n_92),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_88),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_87),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_80),
.A2(n_81),
.B1(n_125),
.B2(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_80),
.A2(n_176),
.B(n_178),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_80),
.A2(n_178),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_81),
.A2(n_104),
.B(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_81),
.A2(n_162),
.B(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_89),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_89),
.A2(n_263),
.B(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_93),
.A2(n_94),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.C(n_105),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_95),
.A2(n_96),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_97),
.Y(n_171)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_103),
.B(n_105),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_110),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_115),
.C(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_130),
.B2(n_132),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_127),
.C(n_130),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_122),
.A2(n_123),
.B1(n_177),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_122),
.A2(n_123),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_123),
.B(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_127),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_127),
.B(n_140),
.C(n_146),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_130),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_132),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_130),
.B(n_136),
.C(n_139),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_134),
.A2(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_148),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_135),
.B(n_148),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_141),
.Y(n_343)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_147),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_326),
.B(n_332),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_198),
.B(n_325),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_191),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_152),
.B(n_191),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_170),
.C(n_172),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_153),
.A2(n_154),
.B1(n_170),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_160),
.C(n_164),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_165),
.B(n_168),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_185)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_170),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_172),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_179),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_173),
.B(n_175),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_179),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_181),
.B1(n_185),
.B2(n_215),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_193),
.B(n_194),
.C(n_197),
.Y(n_331)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_230),
.B(n_319),
.C(n_324),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_224),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_224),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_213),
.C(n_216),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_201),
.A2(n_202),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_211),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_207),
.C(n_211),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_216),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.C(n_221),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_223),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_312),
.B(n_318),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_264),
.B(n_311),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_253),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_235),
.B(n_253),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_246),
.C(n_250),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_236),
.B(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_239),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B(n_244),
.Y(n_239)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_245),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_246),
.A2(n_250),
.B1(n_251),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_249),
.Y(n_262)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_259),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_254),
.B(n_260),
.C(n_261),
.Y(n_317)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_305),
.B(n_310),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_284),
.B(n_304),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_278),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_278),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_273),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_272),
.C(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_282),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_292),
.B(n_303),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_290),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_290),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_298),
.B(n_302),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_295),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_309),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_317),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_317),
.Y(n_318)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_321),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_331),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_331),
.Y(n_332)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_328),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_338),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_347),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_342),
.B1(n_345),
.B2(n_346),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_340),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_342),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_345),
.C(n_347),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_355),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_352),
.B(n_354),
.Y(n_355)
);


endmodule