module fake_jpeg_868_n_54 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_54);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_15;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_14),
.Y(n_25)
);

NOR2x1_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_19),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_16),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_31),
.C(n_16),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_20),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_36),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_15),
.C(n_12),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_0),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_31),
.B1(n_15),
.B2(n_21),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_30),
.B1(n_17),
.B2(n_21),
.Y(n_41)
);

AOI221xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_17),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_45),
.C(n_4),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_46),
.B1(n_1),
.B2(n_3),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_1),
.Y(n_46)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_45),
.B(n_6),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_48),
.C(n_6),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_51),
.C(n_9),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_8),
.B(n_10),
.Y(n_54)
);


endmodule