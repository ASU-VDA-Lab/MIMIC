module fake_jpeg_26661_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_3),
.B(n_2),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_16),
.B(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_21),
.Y(n_27)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.C(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_13),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_29),
.C(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_10),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_11),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_34),
.B1(n_16),
.B2(n_23),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_29),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_9),
.C(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_8),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_19),
.B1(n_20),
.B2(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_38),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_7),
.B1(n_9),
.B2(n_4),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_31),
.B1(n_6),
.B2(n_35),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_6),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_43),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_45),
.C(n_40),
.Y(n_46)
);

NOR4xp25_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_36),
.C(n_37),
.D(n_45),
.Y(n_47)
);


endmodule