module real_jpeg_24349_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_244;
wire n_202;
wire n_167;
wire n_213;
wire n_179;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_1),
.A2(n_20),
.B1(n_24),
.B2(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_34),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_1),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_1),
.A2(n_34),
.B1(n_54),
.B2(n_55),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_20),
.B1(n_24),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_5),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_6),
.A2(n_20),
.B1(n_24),
.B2(n_30),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_6),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_6),
.A2(n_30),
.B1(n_54),
.B2(n_55),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_6),
.B(n_20),
.C(n_23),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_6),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_6),
.B(n_38),
.C(n_40),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_6),
.B(n_52),
.C(n_55),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_44),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_6),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_6),
.B(n_115),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_85),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_83),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_72),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_14),
.B(n_72),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_16),
.B1(n_60),
.B2(n_61),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_31),
.C(n_47),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_17),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_17),
.A2(n_76),
.B1(n_94),
.B2(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_17),
.B(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_17),
.A2(n_76),
.B1(n_110),
.B2(n_111),
.Y(n_133)
);

AOI211xp5_ASAP7_75t_L g155 ( 
.A1(n_17),
.A2(n_124),
.B(n_127),
.C(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_17),
.A2(n_76),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_17),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_17),
.A2(n_76),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_17),
.A2(n_92),
.B(n_95),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_29),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_19),
.A2(n_25),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_19),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_20),
.A2(n_24),
.B1(n_38),
.B2(n_42),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_20),
.B(n_187),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_27),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_31),
.A2(n_32),
.B1(n_47),
.B2(n_48),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_44),
.B2(n_45),
.Y(n_32)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_37),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_36),
.A2(n_37),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_40),
.B1(n_52),
.B2(n_53),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_40),
.B(n_198),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_47),
.A2(n_48),
.B1(n_79),
.B2(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_76),
.C(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_59),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_50),
.B(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_51),
.A2(n_57),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_55),
.B(n_208),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_70),
.Y(n_61)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_71),
.B(n_81),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.C(n_78),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_110),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_78),
.B(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_79),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI31xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_245),
.A3(n_256),
.B(n_261),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_146),
.B(n_244),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_129),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_88),
.B(n_129),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_118),
.B1(n_119),
.B2(n_128),
.Y(n_88)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_108),
.B2(n_109),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_91),
.B(n_108),
.C(n_118),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_106),
.B2(n_107),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_95),
.B1(n_102),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_99),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_98),
.B(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_122),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_101),
.Y(n_209)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_112),
.B(n_117),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_112),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_154),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_110),
.A2(n_111),
.B1(n_124),
.B2(n_154),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_110),
.A2(n_111),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_159),
.C(n_174),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_111),
.A2(n_124),
.B(n_156),
.C(n_219),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_117),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_117),
.A2(n_250),
.B1(n_254),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_125),
.B(n_126),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_120),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_121),
.A2(n_124),
.B1(n_154),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_121),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_140),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_124),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_124),
.A2(n_154),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_124),
.A2(n_154),
.B1(n_196),
.B2(n_197),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_124),
.A2(n_154),
.B1(n_184),
.B2(n_225),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_125),
.A2(n_126),
.B(n_158),
.Y(n_236)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_138),
.B(n_145),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.C(n_137),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_130),
.A2(n_131),
.B1(n_135),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_133),
.B1(n_158),
.B2(n_165),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_132),
.A2(n_133),
.B1(n_138),
.B2(n_139),
.Y(n_233)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_135),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_137),
.B(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_238),
.B(n_243),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_177),
.B(n_229),
.C(n_237),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_167),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_149),
.B(n_167),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_157),
.B2(n_166),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_152),
.B(n_155),
.C(n_166),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_181),
.C(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_154),
.B(n_160),
.C(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_160),
.B1(n_174),
.B2(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_160),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_159),
.B(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_159),
.A2(n_160),
.B1(n_185),
.B2(n_186),
.Y(n_219)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_160),
.B(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_160),
.B(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.C(n_172),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_169),
.A2(n_170),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_190),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_228),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_191),
.B(n_227),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_188),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_180),
.B(n_188),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_221),
.B(n_226),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_215),
.B(n_220),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_204),
.B(n_214),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_199),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_223),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_231),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_234),
.C(n_236),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_242),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_249),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.C(n_255),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_258),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_260),
.Y(n_262)
);


endmodule