module fake_jpeg_12040_n_433 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_433);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_433;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_46),
.Y(n_138)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_48),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_13),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_57),
.B(n_65),
.Y(n_120)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx11_ASAP7_75t_SL g71 ( 
.A(n_26),
.Y(n_71)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_78),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_15),
.B(n_12),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_12),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_88),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_45),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_18),
.B(n_0),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_54),
.B(n_44),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_116),
.B(n_21),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_47),
.A2(n_35),
.B(n_36),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_66),
.Y(n_145)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_64),
.B(n_34),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_66),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_50),
.A2(n_70),
.B1(n_51),
.B2(n_55),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_45),
.B1(n_84),
.B2(n_20),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_145),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_59),
.B1(n_62),
.B2(n_46),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_148),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_69),
.B1(n_44),
.B2(n_85),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_149),
.A2(n_136),
.B1(n_133),
.B2(n_132),
.Y(n_206)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_36),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_151),
.B(n_168),
.Y(n_204)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_153),
.A2(n_155),
.B1(n_171),
.B2(n_183),
.Y(n_227)
);

BUFx2_ASAP7_75t_SL g154 ( 
.A(n_97),
.Y(n_154)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_45),
.B1(n_39),
.B2(n_35),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_89),
.B1(n_87),
.B2(n_71),
.Y(n_156)
);

AO22x1_ASAP7_75t_SL g207 ( 
.A1(n_156),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_207)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_33),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_158),
.B(n_164),
.Y(n_210)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

CKINVDCx12_ASAP7_75t_R g160 ( 
.A(n_92),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_160),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_33),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_174),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_28),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_103),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_175),
.Y(n_193)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_103),
.A2(n_20),
.B1(n_19),
.B2(n_30),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_128),
.Y(n_173)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_111),
.B(n_41),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_177),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_181),
.Y(n_228)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_182),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_116),
.A2(n_20),
.B1(n_30),
.B2(n_42),
.Y(n_183)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_108),
.A2(n_62),
.B1(n_56),
.B2(n_63),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_49),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_124),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_43),
.Y(n_208)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_29),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_217),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_145),
.A2(n_98),
.B1(n_132),
.B2(n_136),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_201),
.A2(n_231),
.B1(n_152),
.B2(n_173),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_206),
.A2(n_181),
.B1(n_144),
.B2(n_166),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_207),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_208),
.B(n_212),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_156),
.A2(n_143),
.B1(n_105),
.B2(n_101),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_209),
.A2(n_211),
.B1(n_161),
.B2(n_150),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_156),
.A2(n_100),
.B1(n_93),
.B2(n_129),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_28),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_113),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_215),
.B(n_218),
.Y(n_247)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_179),
.A2(n_133),
.A3(n_127),
.B1(n_119),
.B2(n_94),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_107),
.Y(n_218)
);

FAx1_ASAP7_75t_L g220 ( 
.A(n_148),
.B(n_90),
.CI(n_80),
.CON(n_220),
.SN(n_220)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_157),
.B(n_161),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_134),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_229),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_149),
.A2(n_130),
.B1(n_185),
.B2(n_167),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_232),
.Y(n_278)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_228),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_257),
.Y(n_273)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_238),
.Y(n_295)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_187),
.B1(n_174),
.B2(n_146),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_241),
.A2(n_242),
.B1(n_214),
.B2(n_195),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_227),
.A2(n_162),
.B1(n_188),
.B2(n_147),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_243),
.A2(n_252),
.B1(n_260),
.B2(n_262),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_244),
.Y(n_292)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_245),
.Y(n_283)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_172),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_248),
.B(n_249),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_193),
.B(n_186),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_163),
.B1(n_159),
.B2(n_30),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_220),
.B1(n_226),
.B2(n_194),
.Y(n_270)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_251),
.Y(n_294)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_176),
.B1(n_72),
.B2(n_49),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_255),
.A2(n_220),
.B1(n_195),
.B2(n_214),
.Y(n_277)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

OR2x4_ASAP7_75t_L g257 ( 
.A(n_198),
.B(n_1),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_192),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_266),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_193),
.B(n_29),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_261),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_199),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_208),
.B(n_29),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_200),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_212),
.B(n_29),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_263),
.B(n_264),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_225),
.Y(n_264)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_265),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_29),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_196),
.A2(n_63),
.B(n_21),
.C(n_4),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_267),
.A2(n_203),
.B(n_200),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_268),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_270),
.A2(n_281),
.B1(n_285),
.B2(n_286),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_229),
.C(n_197),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_288),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_277),
.A2(n_250),
.B1(n_239),
.B2(n_243),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_235),
.A2(n_207),
.B1(n_217),
.B2(n_221),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_282),
.A2(n_297),
.B1(n_299),
.B2(n_236),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_244),
.A2(n_207),
.B(n_221),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_290),
.B(n_259),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_234),
.A2(n_205),
.B1(n_199),
.B2(n_213),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_234),
.A2(n_205),
.B1(n_213),
.B2(n_194),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_240),
.B(n_222),
.C(n_3),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_237),
.A2(n_222),
.B1(n_3),
.B2(n_4),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_1),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_293),
.B(n_255),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_235),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_11),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_298),
.B(n_238),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_233),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_279),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_315),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_302),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_264),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_303),
.B(n_308),
.Y(n_334)
);

AND2x6_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_267),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_309),
.Y(n_328)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_307),
.A2(n_325),
.B1(n_285),
.B2(n_286),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_248),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_292),
.A2(n_247),
.B1(n_236),
.B2(n_245),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_310),
.Y(n_331)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_266),
.Y(n_313)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_268),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_282),
.A2(n_257),
.B1(n_247),
.B2(n_267),
.Y(n_316)
);

XNOR2x1_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_297),
.Y(n_333)
);

AO22x1_ASAP7_75t_L g337 ( 
.A1(n_317),
.A2(n_290),
.B1(n_271),
.B2(n_270),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_274),
.Y(n_319)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_274),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_323),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_281),
.A2(n_261),
.B1(n_263),
.B2(n_251),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_321),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_273),
.B(n_293),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_322),
.B(n_265),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_R g323 ( 
.A(n_276),
.B(n_253),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_284),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_277),
.A2(n_254),
.B1(n_260),
.B2(n_238),
.Y(n_325)
);

INVx4_ASAP7_75t_SL g326 ( 
.A(n_295),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_326),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_272),
.B(n_296),
.Y(n_327)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_327),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_310),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_329),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_335),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_336),
.A2(n_306),
.B1(n_307),
.B2(n_325),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_337),
.A2(n_304),
.B(n_302),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_340),
.A2(n_344),
.B1(n_318),
.B2(n_309),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_319),
.Y(n_343)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_343),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_316),
.A2(n_289),
.B1(n_283),
.B2(n_288),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_345),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_272),
.Y(n_349)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_349),
.Y(n_358)
);

BUFx12f_ASAP7_75t_L g352 ( 
.A(n_332),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_332),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_301),
.C(n_323),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_360),
.C(n_364),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_355),
.A2(n_340),
.B1(n_331),
.B2(n_350),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_351),
.A2(n_317),
.B(n_306),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_356),
.A2(n_359),
.B1(n_370),
.B2(n_337),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_301),
.C(n_324),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_314),
.Y(n_361)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_361),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_363),
.A2(n_336),
.B(n_328),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_342),
.B(n_280),
.C(n_311),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_349),
.Y(n_365)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_368),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_295),
.C(n_278),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_343),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_371),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_344),
.A2(n_283),
.B1(n_299),
.B2(n_326),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_373),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_374),
.A2(n_384),
.B1(n_352),
.B2(n_260),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_328),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_379),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_333),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_SL g391 ( 
.A(n_378),
.B(n_383),
.Y(n_391)
);

A2O1A1O1Ixp25_ASAP7_75t_L g379 ( 
.A1(n_363),
.A2(n_350),
.B(n_331),
.C(n_337),
.D(n_334),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_380),
.A2(n_382),
.B1(n_354),
.B2(n_352),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_359),
.A2(n_339),
.B1(n_330),
.B2(n_348),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_339),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_355),
.A2(n_341),
.B1(n_330),
.B2(n_348),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_265),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_368),
.C(n_364),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_389),
.B(n_385),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_377),
.B(n_366),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_390),
.B(n_393),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_375),
.A2(n_367),
.B1(n_357),
.B2(n_358),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_392),
.A2(n_398),
.B1(n_399),
.B2(n_232),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_370),
.C(n_361),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_354),
.C(n_341),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_384),
.C(n_383),
.Y(n_403)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_396),
.Y(n_402)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_397),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_386),
.A2(n_373),
.B1(n_381),
.B2(n_378),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_379),
.A2(n_262),
.B1(n_256),
.B2(n_246),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_374),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_400),
.A2(n_408),
.B(n_7),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_401),
.B(n_403),
.Y(n_414)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_406),
.B(n_399),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_376),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_407),
.B(n_409),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_395),
.A2(n_262),
.B(n_232),
.Y(n_408)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_410),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_400),
.Y(n_412)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_412),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_393),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_417),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_404),
.B(n_394),
.C(n_391),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_415),
.B(n_416),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_5),
.C(n_6),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_413),
.B(n_402),
.C(n_405),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_411),
.Y(n_425)
);

AOI31xp67_ASAP7_75t_L g423 ( 
.A1(n_420),
.A2(n_412),
.A3(n_414),
.B(n_408),
.Y(n_423)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_423),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_422),
.B(n_401),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_424),
.B(n_425),
.Y(n_426)
);

AOI21xp33_ASAP7_75t_L g428 ( 
.A1(n_427),
.A2(n_419),
.B(n_421),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_428),
.A2(n_426),
.B(n_416),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_421),
.B(n_411),
.Y(n_430)
);

NAND3xp33_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_8),
.C(n_9),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_8),
.C(n_9),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_9),
.C(n_11),
.Y(n_433)
);


endmodule