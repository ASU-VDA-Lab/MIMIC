module fake_jpeg_13243_n_198 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_198);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_15),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_22),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_8),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_14),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_33),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_89),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_92),
.Y(n_104)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_84),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_106),
.Y(n_120)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_95),
.A2(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_64),
.B(n_63),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_76),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_83),
.B1(n_80),
.B2(n_84),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_75),
.B1(n_77),
.B2(n_85),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_108),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_76),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_94),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_94),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_115),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_126),
.B1(n_1),
.B2(n_2),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_66),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_117),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_81),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_121),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_74),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_70),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_124),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_123),
.B(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_73),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_72),
.B1(n_67),
.B2(n_65),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_100),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_60),
.B(n_2),
.Y(n_130)
);

AOI32xp33_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_7),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

OR2x4_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_25),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_141),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_111),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_11),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_145),
.B(n_39),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_149),
.Y(n_165)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_152),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_12),
.Y(n_159)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_132),
.C(n_34),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_162),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_166),
.C(n_169),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_140),
.Y(n_160)
);

BUFx4f_ASAP7_75t_SL g161 ( 
.A(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_163),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_13),
.B1(n_20),
.B2(n_21),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_26),
.C(n_27),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_56),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_37),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_172),
.B(n_50),
.Y(n_180)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_181),
.Y(n_185)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_146),
.B(n_149),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_165),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_158),
.C(n_167),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_187),
.C(n_159),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_167),
.C(n_169),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_186),
.Y(n_192)
);

OAI311xp33_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_176),
.A3(n_185),
.B1(n_181),
.C1(n_175),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_173),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_51),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_55),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_176),
.Y(n_198)
);


endmodule