module fake_jpeg_25650_n_306 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_306);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_27),
.B1(n_33),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_36),
.B1(n_26),
.B2(n_27),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_59),
.Y(n_71)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_57),
.Y(n_79)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_29),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_28),
.B1(n_27),
.B2(n_18),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_29),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_69),
.B1(n_73),
.B2(n_42),
.Y(n_89)
);

NAND2xp67_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_63),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_74),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_36),
.B1(n_28),
.B2(n_32),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_70),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_36),
.B1(n_42),
.B2(n_32),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_41),
.C(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_81),
.Y(n_83)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_43),
.C(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_47),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_84),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_87),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_42),
.B1(n_54),
.B2(n_56),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_69),
.B1(n_65),
.B2(n_70),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_11),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_92),
.B1(n_75),
.B2(n_81),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_46),
.B1(n_38),
.B2(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_101),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_46),
.B1(n_53),
.B2(n_34),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_11),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_99),
.Y(n_131)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_7),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_92),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_108),
.A2(n_123),
.B1(n_124),
.B2(n_38),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_109),
.A2(n_133),
.B1(n_136),
.B2(n_103),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_137),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_25),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_132),
.B(n_67),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_11),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_23),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_82),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_11),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_64),
.B1(n_77),
.B2(n_37),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_23),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_91),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_135),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_25),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_18),
.B1(n_14),
.B2(n_17),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_80),
.C(n_67),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_109),
.C(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_18),
.B1(n_14),
.B2(n_17),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_126),
.B(n_127),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_139),
.A2(n_140),
.B(n_154),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_152),
.Y(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_146),
.Y(n_197)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_148),
.Y(n_175)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_84),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_114),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_20),
.C(n_13),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_84),
.C(n_105),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_45),
.C(n_21),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_166),
.B1(n_80),
.B2(n_18),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_165),
.Y(n_186)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_6),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_163),
.A2(n_167),
.B(n_169),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_172),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_117),
.B1(n_107),
.B2(n_108),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_110),
.A2(n_103),
.B1(n_99),
.B2(n_97),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_23),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_22),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_23),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_80),
.B1(n_17),
.B2(n_14),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_22),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_23),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_21),
.B(n_17),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_177),
.A2(n_199),
.B1(n_150),
.B2(n_148),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_149),
.B(n_20),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_190),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_166),
.B1(n_143),
.B2(n_162),
.Y(n_184)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_22),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_201),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_171),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_21),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_194),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g193 ( 
.A(n_152),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_202),
.B(n_16),
.Y(n_225)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_21),
.B1(n_16),
.B2(n_13),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_200),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_210),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_185),
.C(n_196),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_208),
.C(n_212),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_141),
.C(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_164),
.C(n_140),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_218),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_142),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_159),
.B1(n_163),
.B2(n_168),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_180),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_179),
.A2(n_147),
.B(n_1),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_207),
.B(n_187),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_147),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_14),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_209),
.B(n_217),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_201),
.C(n_179),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_241),
.C(n_243),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_182),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_237),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_207),
.A2(n_182),
.B(n_188),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_240),
.A2(n_224),
.B(n_195),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_191),
.C(n_181),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_233),
.B1(n_219),
.B2(n_206),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_178),
.C(n_175),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_229),
.B(n_213),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_250),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_16),
.B1(n_13),
.B2(n_12),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_211),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_249),
.A2(n_228),
.B1(n_241),
.B2(n_239),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_238),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_257),
.C(n_254),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_7),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_240),
.A2(n_223),
.B(n_214),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_253),
.A2(n_230),
.B(n_244),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_203),
.C(n_175),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_257),
.C(n_259),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_199),
.C(n_45),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_45),
.C(n_16),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_272),
.B(n_268),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_248),
.B(n_227),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_266),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_252),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_270),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_231),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_265),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_12),
.C(n_2),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_7),
.B(n_1),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_269),
.A2(n_253),
.B(n_12),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_13),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_275),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_258),
.B1(n_259),
.B2(n_245),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_279),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_281),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_6),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_2),
.Y(n_291)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_267),
.B(n_262),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_285),
.A2(n_289),
.B(n_284),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_288),
.B(n_280),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_5),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_7),
.B(n_2),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_292),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_3),
.C(n_4),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_293),
.A2(n_294),
.B(n_295),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_281),
.C(n_3),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_296),
.A2(n_298),
.B(n_3),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_284),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_297),
.C(n_3),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_299),
.C(n_4),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_8),
.B(n_9),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_8),
.B(n_9),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_0),
.B(n_8),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_0),
.Y(n_306)
);


endmodule