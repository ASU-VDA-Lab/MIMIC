module real_jpeg_9856_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_23),
.B1(n_49),
.B2(n_62),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_1),
.A2(n_36),
.B1(n_39),
.B2(n_49),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_3),
.A2(n_36),
.B1(n_39),
.B2(n_56),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_4),
.A2(n_36),
.B1(n_39),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_10),
.A2(n_36),
.B1(n_39),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_10),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_11),
.A2(n_23),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_61),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_11),
.A2(n_36),
.B1(n_39),
.B2(n_61),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_12),
.B(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_12),
.A2(n_27),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_12),
.B(n_27),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_12),
.A2(n_40),
.B1(n_74),
.B2(n_120),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_13),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_96),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_95),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_63),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_18),
.B(n_63),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.C(n_57),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_19),
.A2(n_20),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_33),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_28),
.B2(n_32),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_22),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

HAxp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_25),
.CON(n_22),
.SN(n_22)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_30),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_23),
.A2(n_30),
.B(n_32),
.C(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_23),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_23),
.A2(n_62),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_25),
.B(n_53),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_25),
.B(n_74),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_25),
.B(n_70),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_SL g50 ( 
.A1(n_27),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_51),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_59)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_40),
.B(n_43),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_35),
.B(n_42),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_36),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_39),
.B1(n_51),
.B2(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_36),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_39),
.B(n_54),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_39),
.B(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_40),
.A2(n_74),
.B1(n_102),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_40),
.A2(n_104),
.B(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_41),
.B(n_44),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_41),
.A2(n_42),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_46),
.A2(n_47),
.B1(n_57),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_53),
.B2(n_55),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_48),
.A2(n_50),
.B1(n_53),
.B2(n_110),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_55),
.B(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_50),
.A2(n_53),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_57),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_86),
.B2(n_87),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_72),
.B2(n_85),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_136),
.B(n_141),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_127),
.B(n_135),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_116),
.B(n_126),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_105),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_111),
.B2(n_115),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_115),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_121),
.B(n_125),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_118),
.B(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_129),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_130),
.B(n_137),
.Y(n_141)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.CI(n_133),
.CON(n_130),
.SN(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);


endmodule