module fake_jpeg_16885_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_11),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_5),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_53),
.Y(n_75)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_27),
.B1(n_31),
.B2(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_2),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_60),
.Y(n_87)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_15),
.B(n_29),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_37),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_20),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_30),
.B1(n_34),
.B2(n_19),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_15),
.B(n_6),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_33),
.C(n_26),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_32),
.C(n_35),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_71),
.Y(n_108)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_66),
.B(n_76),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_67),
.A2(n_23),
.B1(n_68),
.B2(n_92),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_48),
.Y(n_76)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_37),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_33),
.C(n_25),
.Y(n_104)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_34),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_28),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_94),
.Y(n_116)
);

BUFx16f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_97),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_87),
.B(n_79),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_30),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_100),
.Y(n_126)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_63),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_109),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_33),
.C(n_25),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_119),
.C(n_79),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_54),
.B1(n_31),
.B2(n_27),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_107),
.B(n_121),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_44),
.B1(n_25),
.B2(n_10),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_109),
.A2(n_115),
.B(n_110),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_8),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_117),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_16),
.B1(n_35),
.B2(n_23),
.Y(n_114)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_120),
.B(n_116),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_12),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_16),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_16),
.B1(n_23),
.B2(n_14),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_67),
.A2(n_14),
.B1(n_23),
.B2(n_92),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_94),
.Y(n_122)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_125),
.A3(n_130),
.B1(n_124),
.B2(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_124),
.B(n_91),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_69),
.Y(n_125)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_123),
.B(n_103),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_84),
.A2(n_78),
.B1(n_65),
.B2(n_64),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_96),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_110),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_119),
.B(n_70),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_137),
.C(n_146),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_142),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_70),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_147),
.B1(n_154),
.B2(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_152),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_145),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_84),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_151),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_126),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_106),
.C(n_129),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_131),
.B1(n_134),
.B2(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_117),
.B(n_111),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_149),
.B(n_155),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_111),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_157),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_133),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_164),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_137),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_172),
.Y(n_191)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_159),
.B1(n_154),
.B2(n_139),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_181),
.B1(n_160),
.B2(n_138),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_134),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_136),
.Y(n_195)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_183),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_134),
.A2(n_148),
.B1(n_159),
.B2(n_156),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_196),
.B1(n_163),
.B2(n_173),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_189),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_135),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_152),
.B(n_155),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_195),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_136),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_177),
.B(n_167),
.C(n_165),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_147),
.B1(n_151),
.B2(n_145),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_169),
.B(n_149),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_200),
.B(n_191),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_147),
.B(n_171),
.C(n_164),
.D(n_181),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_170),
.B(n_161),
.C(n_168),
.D(n_178),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_147),
.C(n_174),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_197),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_207),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_209),
.B(n_212),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_168),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_205),
.C(n_193),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

BUFx12_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_196),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_213),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_192),
.C(n_184),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_218),
.C(n_222),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_SL g215 ( 
.A1(n_206),
.A2(n_199),
.B(n_190),
.C(n_189),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_215),
.A2(n_219),
.B1(n_216),
.B2(n_208),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_194),
.C(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_217),
.B(n_212),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_226),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_233)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_207),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_218),
.C(n_204),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_224),
.C(n_202),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_215),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g236 ( 
.A1(n_231),
.A2(n_232),
.A3(n_210),
.B1(n_213),
.B2(n_233),
.C1(n_234),
.C2(n_230),
.Y(n_236)
);

NOR2x1_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_211),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_237),
.B(n_231),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_232),
.C(n_210),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_238),
.Y(n_241)
);


endmodule