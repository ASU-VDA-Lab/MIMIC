module real_aes_8111_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g104 ( .A(n_0), .Y(n_104) );
INVx1_ASAP7_75t_L g434 ( .A(n_1), .Y(n_434) );
INVx1_ASAP7_75t_L g237 ( .A(n_2), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_3), .A2(n_36), .B1(n_187), .B2(n_473), .Y(n_509) );
AOI21xp33_ASAP7_75t_L g198 ( .A1(n_4), .A2(n_120), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_5), .B(n_142), .Y(n_459) );
AND2x6_ASAP7_75t_L g125 ( .A(n_6), .B(n_126), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_7), .A2(n_119), .B(n_127), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_8), .B(n_37), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_9), .B(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g204 ( .A(n_10), .Y(n_204) );
INVx1_ASAP7_75t_L g117 ( .A(n_11), .Y(n_117) );
INVx1_ASAP7_75t_L g428 ( .A(n_12), .Y(n_428) );
INVx1_ASAP7_75t_L g137 ( .A(n_13), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_14), .B(n_211), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_15), .B(n_143), .Y(n_461) );
AO32x2_ASAP7_75t_L g507 ( .A1(n_16), .A2(n_142), .A3(n_158), .B1(n_447), .B2(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_17), .B(n_187), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_18), .B(n_154), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_19), .B(n_143), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_20), .A2(n_48), .B1(n_187), .B2(n_473), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_21), .B(n_120), .Y(n_147) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_22), .A2(n_73), .B1(n_187), .B2(n_211), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_23), .B(n_187), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_24), .B(n_197), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g133 ( .A1(n_25), .A2(n_134), .B(n_136), .C(n_138), .Y(n_133) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_26), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_27), .B(n_113), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_28), .B(n_169), .Y(n_238) );
AOI222xp33_ASAP7_75t_SL g100 ( .A1(n_29), .A2(n_87), .B1(n_101), .B2(n_693), .C1(n_694), .C2(n_697), .Y(n_100) );
INVx1_ASAP7_75t_L g693 ( .A(n_29), .Y(n_693) );
INVx1_ASAP7_75t_L g216 ( .A(n_30), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_31), .B(n_113), .Y(n_485) );
INVx2_ASAP7_75t_L g123 ( .A(n_32), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_33), .B(n_187), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_34), .B(n_113), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_35), .A2(n_125), .B(n_130), .C(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g214 ( .A(n_38), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_39), .B(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_40), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_41), .B(n_187), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_42), .A2(n_83), .B1(n_139), .B2(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_43), .B(n_187), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_44), .B(n_187), .Y(n_429) );
CKINVDCx16_ASAP7_75t_R g217 ( .A(n_45), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_46), .B(n_433), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_47), .B(n_120), .Y(n_188) );
AOI22xp33_ASAP7_75t_SL g465 ( .A1(n_49), .A2(n_58), .B1(n_187), .B2(n_211), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_50), .A2(n_130), .B1(n_211), .B2(n_213), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_51), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_52), .B(n_187), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_53), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_54), .B(n_187), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_55), .A2(n_202), .B(n_203), .C(n_205), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_56), .Y(n_173) );
INVx1_ASAP7_75t_L g200 ( .A(n_57), .Y(n_200) );
INVx1_ASAP7_75t_L g126 ( .A(n_59), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_60), .B(n_187), .Y(n_435) );
INVx1_ASAP7_75t_L g116 ( .A(n_61), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_62), .Y(n_706) );
AO32x2_ASAP7_75t_L g470 ( .A1(n_63), .A2(n_142), .A3(n_179), .B1(n_447), .B2(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g445 ( .A(n_64), .Y(n_445) );
INVx1_ASAP7_75t_L g480 ( .A(n_65), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_SL g224 ( .A1(n_66), .A2(n_154), .B(n_205), .C(n_225), .Y(n_224) );
INVxp67_ASAP7_75t_L g226 ( .A(n_67), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_68), .B(n_211), .Y(n_481) );
INVx1_ASAP7_75t_L g705 ( .A(n_69), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_70), .Y(n_219) );
INVx1_ASAP7_75t_L g164 ( .A(n_71), .Y(n_164) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_72), .A2(n_99), .B1(n_701), .B2(n_710), .C1(n_719), .C2(n_725), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_72), .A2(n_106), .B1(n_695), .B2(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_72), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_74), .A2(n_125), .B(n_130), .C(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_75), .B(n_473), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_76), .B(n_211), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_77), .B(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g114 ( .A(n_78), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_79), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_80), .B(n_211), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_81), .A2(n_125), .B(n_130), .C(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g102 ( .A(n_82), .B(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g417 ( .A(n_82), .Y(n_417) );
OR2x2_ASAP7_75t_L g709 ( .A(n_82), .B(n_700), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_84), .A2(n_97), .B1(n_211), .B2(n_212), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_85), .B(n_113), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_86), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_88), .A2(n_125), .B(n_130), .C(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_89), .Y(n_190) );
INVx1_ASAP7_75t_L g223 ( .A(n_90), .Y(n_223) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_91), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_92), .B(n_151), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_93), .B(n_211), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_94), .B(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_95), .A2(n_120), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_96), .B(n_705), .Y(n_704) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_106), .B1(n_414), .B2(n_418), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g694 ( .A1(n_102), .A2(n_416), .B1(n_695), .B2(n_696), .Y(n_694) );
OR2x2_ASAP7_75t_L g416 ( .A(n_103), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g700 ( .A(n_103), .Y(n_700) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx2_ASAP7_75t_SL g695 ( .A(n_106), .Y(n_695) );
OR4x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_310), .C(n_369), .D(n_396), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_252), .C(n_277), .Y(n_107) );
O2A1O1Ixp33_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_175), .B(n_195), .C(n_228), .Y(n_108) );
AOI211xp5_ASAP7_75t_SL g400 ( .A1(n_109), .A2(n_401), .B(n_403), .C(n_406), .Y(n_400) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_144), .Y(n_109) );
INVx1_ASAP7_75t_L g275 ( .A(n_110), .Y(n_275) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g250 ( .A(n_111), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g282 ( .A(n_111), .Y(n_282) );
AND2x2_ASAP7_75t_L g337 ( .A(n_111), .B(n_306), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_111), .B(n_193), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_111), .B(n_194), .Y(n_395) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g256 ( .A(n_112), .Y(n_256) );
AND2x2_ASAP7_75t_L g299 ( .A(n_112), .B(n_162), .Y(n_299) );
AND2x2_ASAP7_75t_L g317 ( .A(n_112), .B(n_194), .Y(n_317) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_118), .B(n_141), .Y(n_112) );
INVx1_ASAP7_75t_L g174 ( .A(n_113), .Y(n_174) );
INVx2_ASAP7_75t_L g179 ( .A(n_113), .Y(n_179) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_113), .A2(n_478), .B(n_485), .Y(n_477) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_113), .A2(n_487), .B(n_495), .Y(n_486) );
AND2x2_ASAP7_75t_SL g113 ( .A(n_114), .B(n_115), .Y(n_113) );
AND2x2_ASAP7_75t_L g143 ( .A(n_114), .B(n_115), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_125), .Y(n_120) );
NAND2x1p5_ASAP7_75t_L g165 ( .A(n_121), .B(n_125), .Y(n_165) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
INVx1_ASAP7_75t_L g433 ( .A(n_122), .Y(n_433) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g131 ( .A(n_123), .Y(n_131) );
INVx1_ASAP7_75t_L g212 ( .A(n_123), .Y(n_212) );
INVx1_ASAP7_75t_L g132 ( .A(n_124), .Y(n_132) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_124), .Y(n_135) );
INVx3_ASAP7_75t_L g152 ( .A(n_124), .Y(n_152) );
INVx1_ASAP7_75t_L g154 ( .A(n_124), .Y(n_154) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
INVx4_ASAP7_75t_SL g140 ( .A(n_125), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g426 ( .A1(n_125), .A2(n_427), .B(n_431), .Y(n_426) );
BUFx3_ASAP7_75t_L g447 ( .A(n_125), .Y(n_447) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_125), .A2(n_453), .B(n_456), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_125), .A2(n_479), .B(n_482), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_125), .A2(n_488), .B(n_492), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B(n_133), .C(n_140), .Y(n_127) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_129), .A2(n_140), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_129), .A2(n_140), .B(n_223), .C(n_224), .Y(n_222) );
INVx5_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
BUFx3_ASAP7_75t_L g139 ( .A(n_131), .Y(n_139) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
INVx1_ASAP7_75t_L g473 ( .A(n_131), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_134), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g430 ( .A(n_134), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_134), .A2(n_483), .B(n_484), .Y(n_482) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g213 ( .A1(n_135), .A2(n_214), .B1(n_215), .B2(n_216), .Y(n_213) );
INVx2_ASAP7_75t_L g215 ( .A(n_135), .Y(n_215) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g156 ( .A(n_139), .Y(n_156) );
OAI22xp33_ASAP7_75t_L g209 ( .A1(n_140), .A2(n_165), .B1(n_210), .B2(n_217), .Y(n_209) );
INVx4_ASAP7_75t_L g161 ( .A(n_142), .Y(n_161) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_142), .A2(n_221), .B(n_227), .Y(n_220) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_142), .A2(n_452), .B(n_459), .Y(n_451) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g158 ( .A(n_143), .Y(n_158) );
INVx4_ASAP7_75t_L g249 ( .A(n_144), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_144), .A2(n_305), .B(n_307), .Y(n_304) );
AND2x2_ASAP7_75t_L g385 ( .A(n_144), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_162), .Y(n_144) );
INVx1_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
AND2x2_ASAP7_75t_L g254 ( .A(n_145), .B(n_194), .Y(n_254) );
OR2x2_ASAP7_75t_L g283 ( .A(n_145), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g297 ( .A(n_145), .Y(n_297) );
INVx3_ASAP7_75t_L g306 ( .A(n_145), .Y(n_306) );
AND2x2_ASAP7_75t_L g316 ( .A(n_145), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g349 ( .A(n_145), .B(n_255), .Y(n_349) );
AND2x2_ASAP7_75t_L g373 ( .A(n_145), .B(n_329), .Y(n_373) );
OR2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_159), .Y(n_145) );
AOI21xp5_ASAP7_75t_SL g146 ( .A1(n_147), .A2(n_148), .B(n_157), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B(n_155), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_151), .A2(n_237), .B(n_238), .C(n_239), .Y(n_236) );
INVx2_ASAP7_75t_L g436 ( .A(n_151), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_151), .A2(n_442), .B(n_443), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_151), .A2(n_454), .B(n_455), .Y(n_453) );
O2A1O1Ixp5_ASAP7_75t_SL g479 ( .A1(n_151), .A2(n_205), .B(n_480), .C(n_481), .Y(n_479) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_152), .B(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_152), .B(n_226), .Y(n_225) );
OAI22xp5_ASAP7_75t_SL g471 ( .A1(n_152), .A2(n_169), .B1(n_472), .B2(n_474), .Y(n_471) );
INVx1_ASAP7_75t_L g491 ( .A(n_154), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_155), .A2(n_168), .B(n_170), .Y(n_167) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g171 ( .A(n_157), .Y(n_171) );
OA21x2_ASAP7_75t_L g425 ( .A1(n_157), .A2(n_426), .B(n_437), .Y(n_425) );
OA21x2_ASAP7_75t_L g439 ( .A1(n_157), .A2(n_440), .B(n_448), .Y(n_439) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_158), .A2(n_209), .B(n_218), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_158), .B(n_219), .Y(n_218) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_158), .A2(n_233), .B(n_240), .Y(n_232) );
NOR2xp33_ASAP7_75t_SL g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx3_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_161), .B(n_447), .C(n_463), .Y(n_462) );
AO21x1_ASAP7_75t_L g541 ( .A1(n_161), .A2(n_463), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g194 ( .A(n_162), .Y(n_194) );
AND2x2_ASAP7_75t_L g409 ( .A(n_162), .B(n_251), .Y(n_409) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_171), .B(n_172), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_166), .Y(n_163) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_165), .A2(n_234), .B(n_235), .Y(n_233) );
INVx4_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
INVx2_ASAP7_75t_L g202 ( .A(n_169), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_169), .A2(n_436), .B1(n_464), .B2(n_465), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_169), .A2(n_436), .B1(n_509), .B2(n_510), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_174), .B(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_174), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_191), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_177), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g329 ( .A(n_177), .B(n_317), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_177), .B(n_306), .Y(n_391) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g251 ( .A(n_178), .Y(n_251) );
AND2x2_ASAP7_75t_L g255 ( .A(n_178), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g296 ( .A(n_178), .B(n_297), .Y(n_296) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_189), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_188), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_186), .Y(n_182) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx3_ASAP7_75t_L g205 ( .A(n_187), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_191), .B(n_292), .Y(n_314) );
INVx1_ASAP7_75t_L g353 ( .A(n_191), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_191), .B(n_280), .Y(n_397) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
AND2x2_ASAP7_75t_L g260 ( .A(n_192), .B(n_255), .Y(n_260) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_194), .B(n_251), .Y(n_284) );
INVx1_ASAP7_75t_L g363 ( .A(n_194), .Y(n_363) );
AOI322xp5_ASAP7_75t_L g387 ( .A1(n_195), .A2(n_302), .A3(n_362), .B1(n_388), .B2(n_390), .C1(n_392), .C2(n_394), .Y(n_387) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_196), .B(n_207), .Y(n_195) );
AND2x2_ASAP7_75t_L g242 ( .A(n_196), .B(n_220), .Y(n_242) );
INVx1_ASAP7_75t_SL g245 ( .A(n_196), .Y(n_245) );
AND2x2_ASAP7_75t_L g247 ( .A(n_196), .B(n_208), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_196), .B(n_264), .Y(n_270) );
INVx2_ASAP7_75t_L g289 ( .A(n_196), .Y(n_289) );
AND2x2_ASAP7_75t_L g302 ( .A(n_196), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g340 ( .A(n_196), .B(n_264), .Y(n_340) );
BUFx2_ASAP7_75t_L g357 ( .A(n_196), .Y(n_357) );
AND2x2_ASAP7_75t_L g371 ( .A(n_196), .B(n_231), .Y(n_371) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_206), .Y(n_196) );
O2A1O1Ixp5_ASAP7_75t_L g444 ( .A1(n_202), .A2(n_432), .B(n_445), .C(n_446), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_202), .A2(n_493), .B(n_494), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_207), .B(n_259), .Y(n_286) );
AND2x2_ASAP7_75t_L g413 ( .A(n_207), .B(n_289), .Y(n_413) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_220), .Y(n_207) );
OR2x2_ASAP7_75t_L g258 ( .A(n_208), .B(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g264 ( .A(n_208), .Y(n_264) );
AND2x2_ASAP7_75t_L g309 ( .A(n_208), .B(n_232), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_208), .B(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_208), .Y(n_393) );
INVx2_ASAP7_75t_L g239 ( .A(n_211), .Y(n_239) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g244 ( .A(n_220), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g266 ( .A(n_220), .Y(n_266) );
BUFx2_ASAP7_75t_L g272 ( .A(n_220), .Y(n_272) );
AND2x2_ASAP7_75t_L g291 ( .A(n_220), .B(n_264), .Y(n_291) );
INVx3_ASAP7_75t_L g303 ( .A(n_220), .Y(n_303) );
OR2x2_ASAP7_75t_L g313 ( .A(n_220), .B(n_264), .Y(n_313) );
AOI31xp33_ASAP7_75t_SL g228 ( .A1(n_229), .A2(n_243), .A3(n_246), .B(n_248), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_242), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_230), .B(n_265), .Y(n_276) );
OR2x2_ASAP7_75t_L g300 ( .A(n_230), .B(n_270), .Y(n_300) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_231), .B(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g321 ( .A(n_231), .B(n_313), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_231), .B(n_303), .Y(n_331) );
AND2x2_ASAP7_75t_L g338 ( .A(n_231), .B(n_339), .Y(n_338) );
NAND2x1_ASAP7_75t_L g366 ( .A(n_231), .B(n_302), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_231), .B(n_357), .Y(n_367) );
AND2x2_ASAP7_75t_L g379 ( .A(n_231), .B(n_264), .Y(n_379) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx3_ASAP7_75t_L g259 ( .A(n_232), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g427 ( .A1(n_239), .A2(n_428), .B(n_429), .C(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g325 ( .A(n_242), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_242), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_244), .B(n_320), .Y(n_354) );
AND2x4_ASAP7_75t_L g265 ( .A(n_245), .B(n_266), .Y(n_265) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g344 ( .A(n_250), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_250), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g292 ( .A(n_251), .B(n_282), .Y(n_292) );
AND2x2_ASAP7_75t_L g386 ( .A(n_251), .B(n_256), .Y(n_386) );
INVx1_ASAP7_75t_L g411 ( .A(n_251), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_257), .B1(n_260), .B2(n_261), .C(n_267), .Y(n_252) );
CKINVDCx14_ASAP7_75t_R g273 ( .A(n_253), .Y(n_273) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_254), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_257), .B(n_308), .Y(n_327) );
INVx3_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g376 ( .A(n_258), .B(n_272), .Y(n_376) );
AND2x2_ASAP7_75t_L g290 ( .A(n_259), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g320 ( .A(n_259), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_259), .B(n_303), .Y(n_348) );
NOR3xp33_ASAP7_75t_L g390 ( .A(n_259), .B(n_360), .C(n_391), .Y(n_390) );
AOI211xp5_ASAP7_75t_SL g323 ( .A1(n_260), .A2(n_324), .B(n_326), .C(n_334), .Y(n_323) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI22xp33_ASAP7_75t_L g312 ( .A1(n_262), .A2(n_313), .B1(n_314), .B2(n_315), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_263), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_263), .B(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g405 ( .A(n_265), .B(n_379), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_273), .B1(n_274), .B2(n_276), .Y(n_267) );
NOR2xp33_ASAP7_75t_SL g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_271), .B(n_320), .Y(n_351) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_274), .A2(n_366), .B1(n_397), .B2(n_404), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_285), .B1(n_287), .B2(n_292), .C(n_293), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVxp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI221xp5_ASAP7_75t_L g293 ( .A1(n_283), .A2(n_294), .B1(n_300), .B2(n_301), .C(n_304), .Y(n_293) );
INVx1_ASAP7_75t_L g336 ( .A(n_284), .Y(n_336) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_SL g308 ( .A(n_289), .Y(n_308) );
OR2x2_ASAP7_75t_L g381 ( .A(n_289), .B(n_313), .Y(n_381) );
AND2x2_ASAP7_75t_L g383 ( .A(n_289), .B(n_291), .Y(n_383) );
INVx1_ASAP7_75t_L g322 ( .A(n_292), .Y(n_322) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
AOI21xp33_ASAP7_75t_SL g352 ( .A1(n_295), .A2(n_353), .B(n_354), .Y(n_352) );
OR2x2_ASAP7_75t_L g359 ( .A(n_295), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g333 ( .A(n_296), .B(n_317), .Y(n_333) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp33_ASAP7_75t_SL g350 ( .A(n_301), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_302), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_303), .B(n_339), .Y(n_402) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_306), .A2(n_319), .B(n_321), .C(n_322), .Y(n_318) );
NAND2x1_ASAP7_75t_SL g343 ( .A(n_306), .B(n_344), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_307), .A2(n_356), .B1(n_358), .B2(n_361), .Y(n_355) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_309), .B(n_399), .Y(n_398) );
NAND5xp2_ASAP7_75t_L g310 ( .A(n_311), .B(n_323), .C(n_341), .D(n_355), .E(n_364), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_318), .Y(n_311) );
INVx1_ASAP7_75t_L g368 ( .A(n_314), .Y(n_368) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_316), .A2(n_335), .B1(n_375), .B2(n_377), .C(n_380), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_317), .B(n_411), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_320), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_320), .B(n_386), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B1(n_330), .B2(n_332), .Y(n_326) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_338), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
AND2x2_ASAP7_75t_L g408 ( .A(n_337), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_345), .B1(n_349), .B2(n_350), .C(n_352), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g392 ( .A(n_347), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g399 ( .A(n_357), .Y(n_399) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI21xp5_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_367), .B(n_368), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI211xp5_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_372), .B(n_374), .C(n_387), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
A2O1A1Ixp33_ASAP7_75t_L g396 ( .A1(n_372), .A2(n_397), .B(n_398), .C(n_400), .Y(n_396) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_376), .B(n_378), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_384), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI21xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_410), .B(n_412), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NOR2x2_ASAP7_75t_L g699 ( .A(n_417), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g696 ( .A(n_418), .Y(n_696) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OR5x1_ASAP7_75t_L g420 ( .A(n_421), .B(n_584), .C(n_642), .D(n_678), .E(n_685), .Y(n_420) );
NAND3xp33_ASAP7_75t_SL g421 ( .A(n_422), .B(n_530), .C(n_554), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_466), .B1(n_496), .B2(n_501), .C(n_511), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_423), .A2(n_665), .B(n_667), .Y(n_664) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_449), .Y(n_423) );
NAND2x1p5_ASAP7_75t_L g654 ( .A(n_424), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_438), .Y(n_424) );
INVx2_ASAP7_75t_L g500 ( .A(n_425), .Y(n_500) );
AND2x2_ASAP7_75t_L g513 ( .A(n_425), .B(n_451), .Y(n_513) );
AND2x2_ASAP7_75t_L g567 ( .A(n_425), .B(n_450), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_425), .B(n_439), .Y(n_582) );
O2A1O1Ixp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B(n_435), .C(n_436), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_436), .A2(n_457), .B(n_458), .Y(n_456) );
AND2x2_ASAP7_75t_L g600 ( .A(n_438), .B(n_541), .Y(n_600) );
AND2x2_ASAP7_75t_L g633 ( .A(n_438), .B(n_451), .Y(n_633) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g540 ( .A(n_439), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g553 ( .A(n_439), .B(n_451), .Y(n_553) );
AND2x2_ASAP7_75t_L g560 ( .A(n_439), .B(n_541), .Y(n_560) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_439), .Y(n_569) );
AND2x2_ASAP7_75t_L g576 ( .A(n_439), .B(n_450), .Y(n_576) );
INVx1_ASAP7_75t_L g607 ( .A(n_439), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_444), .B(n_447), .Y(n_440) );
INVx1_ASAP7_75t_L g583 ( .A(n_449), .Y(n_583) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_460), .Y(n_449) );
INVx2_ASAP7_75t_L g539 ( .A(n_450), .Y(n_539) );
AND2x2_ASAP7_75t_L g561 ( .A(n_450), .B(n_500), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_450), .B(n_607), .Y(n_612) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_451), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g684 ( .A(n_451), .B(n_648), .Y(n_684) );
INVx2_ASAP7_75t_L g498 ( .A(n_460), .Y(n_498) );
INVx3_ASAP7_75t_L g599 ( .A(n_460), .Y(n_599) );
OR2x2_ASAP7_75t_L g629 ( .A(n_460), .B(n_630), .Y(n_629) );
NOR2x1_ASAP7_75t_L g655 ( .A(n_460), .B(n_539), .Y(n_655) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g542 ( .A(n_461), .Y(n_542) );
AOI33xp33_ASAP7_75t_L g675 ( .A1(n_466), .A2(n_513), .A3(n_527), .B1(n_599), .B2(n_676), .B3(n_677), .Y(n_675) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_475), .Y(n_467) );
OR2x2_ASAP7_75t_L g528 ( .A(n_468), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_468), .B(n_525), .Y(n_587) );
OR2x2_ASAP7_75t_L g640 ( .A(n_468), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g566 ( .A(n_469), .B(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g591 ( .A(n_469), .B(n_475), .Y(n_591) );
AND2x2_ASAP7_75t_L g658 ( .A(n_469), .B(n_503), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_469), .A2(n_558), .B(n_684), .Y(n_683) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g505 ( .A(n_470), .Y(n_505) );
INVx1_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
AND2x2_ASAP7_75t_L g537 ( .A(n_470), .B(n_507), .Y(n_537) );
AND2x2_ASAP7_75t_L g586 ( .A(n_470), .B(n_506), .Y(n_586) );
INVx2_ASAP7_75t_SL g628 ( .A(n_475), .Y(n_628) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
INVx2_ASAP7_75t_L g548 ( .A(n_476), .Y(n_548) );
INVx1_ASAP7_75t_L g679 ( .A(n_476), .Y(n_679) );
AND2x2_ASAP7_75t_L g692 ( .A(n_476), .B(n_573), .Y(n_692) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g519 ( .A(n_477), .Y(n_519) );
OR2x2_ASAP7_75t_L g525 ( .A(n_477), .B(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_477), .Y(n_536) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_486), .Y(n_503) );
AND2x2_ASAP7_75t_L g520 ( .A(n_486), .B(n_506), .Y(n_520) );
INVx1_ASAP7_75t_L g526 ( .A(n_486), .Y(n_526) );
INVx1_ASAP7_75t_L g533 ( .A(n_486), .Y(n_533) );
AND2x2_ASAP7_75t_L g558 ( .A(n_486), .B(n_507), .Y(n_558) );
INVx2_ASAP7_75t_L g574 ( .A(n_486), .Y(n_574) );
AND2x2_ASAP7_75t_L g667 ( .A(n_486), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_486), .B(n_548), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_491), .Y(n_488) );
INVx1_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g522 ( .A(n_498), .Y(n_522) );
INVx1_ASAP7_75t_L g551 ( .A(n_498), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_498), .B(n_582), .Y(n_648) );
INVx1_ASAP7_75t_SL g608 ( .A(n_499), .Y(n_608) );
INVx2_ASAP7_75t_L g529 ( .A(n_500), .Y(n_529) );
AND2x2_ASAP7_75t_L g598 ( .A(n_500), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g614 ( .A(n_500), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
INVx1_ASAP7_75t_L g676 ( .A(n_502), .Y(n_676) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g531 ( .A(n_504), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g634 ( .A(n_504), .B(n_624), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_504), .A2(n_645), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_L g547 ( .A(n_505), .B(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g572 ( .A(n_505), .Y(n_572) );
INVx1_ASAP7_75t_L g596 ( .A(n_505), .Y(n_596) );
OR2x2_ASAP7_75t_L g660 ( .A(n_506), .B(n_519), .Y(n_660) );
NOR2xp67_ASAP7_75t_L g668 ( .A(n_506), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g573 ( .A(n_507), .B(n_574), .Y(n_573) );
BUFx2_ASAP7_75t_L g580 ( .A(n_507), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_514), .B1(n_521), .B2(n_523), .Y(n_511) );
OR2x2_ASAP7_75t_L g590 ( .A(n_512), .B(n_540), .Y(n_590) );
INVx1_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
AOI222xp33_ASAP7_75t_L g631 ( .A1(n_513), .A2(n_632), .B1(n_634), .B2(n_635), .C1(n_636), .C2(n_639), .Y(n_631) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_520), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g578 ( .A(n_517), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
AND2x2_ASAP7_75t_SL g532 ( .A(n_519), .B(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_519), .Y(n_603) );
AND2x2_ASAP7_75t_L g651 ( .A(n_519), .B(n_520), .Y(n_651) );
INVx1_ASAP7_75t_L g669 ( .A(n_519), .Y(n_669) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g635 ( .A(n_522), .B(n_561), .Y(n_635) );
AND2x2_ASAP7_75t_L g677 ( .A(n_522), .B(n_553), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_524), .B(n_572), .Y(n_659) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_525), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g552 ( .A(n_529), .B(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g620 ( .A(n_529), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_534), .B(n_538), .C(n_543), .Y(n_530) );
INVxp67_ASAP7_75t_L g544 ( .A(n_531), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_532), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_532), .B(n_579), .Y(n_674) );
BUFx3_ASAP7_75t_L g638 ( .A(n_533), .Y(n_638) );
INVx1_ASAP7_75t_L g545 ( .A(n_534), .Y(n_545) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g564 ( .A(n_536), .B(n_558), .Y(n_564) );
INVx1_ASAP7_75t_SL g604 ( .A(n_537), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g594 ( .A(n_539), .Y(n_594) );
AND2x2_ASAP7_75t_L g617 ( .A(n_539), .B(n_600), .Y(n_617) );
INVx1_ASAP7_75t_SL g588 ( .A(n_540), .Y(n_588) );
INVx1_ASAP7_75t_L g615 ( .A(n_541), .Y(n_615) );
AOI31xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .A3(n_546), .B(n_549), .Y(n_543) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g636 ( .A(n_547), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g610 ( .A(n_548), .Y(n_610) );
BUFx2_ASAP7_75t_L g624 ( .A(n_548), .Y(n_624) );
AND2x2_ASAP7_75t_L g652 ( .A(n_548), .B(n_573), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_SL g625 ( .A(n_552), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_553), .B(n_620), .Y(n_666) );
AND2x2_ASAP7_75t_L g673 ( .A(n_553), .B(n_599), .Y(n_673) );
AOI211xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_559), .B(n_562), .C(n_577), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_559), .A2(n_586), .B1(n_587), .B2(n_588), .C(n_589), .Y(n_585) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g593 ( .A(n_560), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g630 ( .A(n_561), .Y(n_630) );
OAI32xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .A3(n_568), .B1(n_570), .B2(n_575), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_564), .A2(n_617), .B(n_618), .C(n_621), .Y(n_616) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OAI21xp5_ASAP7_75t_SL g680 ( .A1(n_572), .A2(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g641 ( .A(n_573), .Y(n_641) );
INVxp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_579), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g627 ( .A(n_579), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g644 ( .A(n_581), .Y(n_644) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NAND4xp25_ASAP7_75t_SL g584 ( .A(n_585), .B(n_597), .C(n_616), .D(n_631), .Y(n_584) );
AND2x2_ASAP7_75t_L g623 ( .A(n_586), .B(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g645 ( .A(n_586), .B(n_638), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_588), .B(n_620), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_592), .B2(n_595), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_590), .A2(n_641), .B1(n_672), .B2(n_674), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g678 ( .A1(n_590), .A2(n_679), .B(n_680), .C(n_683), .Y(n_678) );
INVx2_ASAP7_75t_L g649 ( .A(n_591), .Y(n_649) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI222xp33_ASAP7_75t_L g643 ( .A1(n_593), .A2(n_627), .B1(n_644), .B2(n_645), .C1(n_646), .C2(n_649), .Y(n_643) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .B(n_601), .C(n_605), .Y(n_597) );
INVx1_ASAP7_75t_L g663 ( .A(n_598), .Y(n_663) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_602), .A2(n_606), .B1(n_609), .B2(n_611), .Y(n_605) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g632 ( .A(n_614), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g690 ( .A(n_617), .Y(n_690) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_625), .B1(n_626), .B2(n_629), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_624), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g681 ( .A(n_629), .Y(n_681) );
INVx1_ASAP7_75t_L g662 ( .A(n_633), .Y(n_662) );
CKINVDCx16_ASAP7_75t_R g689 ( .A(n_635), .Y(n_689) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND5xp2_ASAP7_75t_L g642 ( .A(n_643), .B(n_650), .C(n_664), .D(n_670), .E(n_675), .Y(n_642) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B(n_653), .C(n_656), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI31xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .A3(n_660), .B(n_661), .Y(n_656) );
INVx1_ASAP7_75t_L g682 ( .A(n_658), .Y(n_682) );
OR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI222xp33_ASAP7_75t_L g685 ( .A1(n_672), .A2(n_674), .B1(n_686), .B2(n_689), .C1(n_690), .C2(n_691), .Y(n_685) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_707), .Y(n_702) );
NOR2xp33_ASAP7_75t_SL g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVx1_ASAP7_75t_SL g724 ( .A(n_704), .Y(n_724) );
INVx1_ASAP7_75t_L g723 ( .A(n_706), .Y(n_723) );
OA21x2_ASAP7_75t_L g726 ( .A1(n_706), .A2(n_724), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g715 ( .A(n_709), .Y(n_715) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_709), .Y(n_717) );
BUFx2_ASAP7_75t_L g727 ( .A(n_709), .Y(n_727) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B(n_716), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NOR2xp33_ASAP7_75t_SL g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
CKINVDCx6p67_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
endmodule