module real_jpeg_10412_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_11;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_2),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_2),
.A2(n_7),
.B(n_28),
.C(n_32),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_2),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_2),
.A2(n_26),
.B1(n_30),
.B2(n_40),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_2),
.A2(n_6),
.B(n_22),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_2),
.B(n_38),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_3),
.A2(n_30),
.B1(n_40),
.B2(n_42),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_22),
.B1(n_25),
.B2(n_42),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_22),
.B1(n_25),
.B2(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_6),
.A2(n_30),
.B(n_52),
.C(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_6),
.B(n_30),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_7),
.A2(n_32),
.B(n_39),
.C(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_7),
.B(n_32),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_9),
.A2(n_30),
.B1(n_40),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_56),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_9),
.A2(n_22),
.B1(n_25),
.B2(n_56),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_91),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_90),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_59),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_14),
.B(n_59),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_35),
.C(n_48),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_15),
.A2(n_16),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_27),
.B2(n_34),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_27),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B(n_24),
.Y(n_18)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_19),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_20),
.B(n_26),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_21),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_21),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_21),
.B(n_77),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_25),
.B(n_117),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_29),
.B(n_30),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_26),
.A2(n_40),
.B(n_53),
.C(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_26),
.B(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_32),
.A2(n_33),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_35),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_52),
.B(n_55),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_85),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_81),
.B2(n_82),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_113),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_87),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_132),
.B(n_137),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_120),
.B(n_131),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_108),
.B(n_119),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_114),
.B(n_118),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_112),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_122),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_127),
.C(n_129),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_134),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);


endmodule