module real_jpeg_26583_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx11_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_1),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_1),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_2),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_SL g87 ( 
.A1(n_2),
.A2(n_60),
.B(n_64),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_2),
.A2(n_56),
.B1(n_58),
.B2(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_2),
.B(n_62),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_2),
.A2(n_44),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_44),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_2),
.B(n_79),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_2),
.A2(n_26),
.B1(n_36),
.B2(n_199),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_2),
.A2(n_63),
.B(n_215),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_4),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_4),
.A2(n_56),
.B1(n_58),
.B2(n_70),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_70),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_4),
.A2(n_28),
.B1(n_34),
.B2(n_70),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_6),
.A2(n_28),
.B1(n_34),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_6),
.Y(n_99)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_77),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_9),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_9),
.A2(n_28),
.B1(n_34),
.B2(n_42),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_28),
.B1(n_34),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_11),
.A2(n_55),
.B1(n_63),
.B2(n_64),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_11),
.A2(n_28),
.B1(n_34),
.B2(n_55),
.Y(n_192)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_13),
.A2(n_56),
.B1(n_58),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_13),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_93),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_93),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_13),
.A2(n_28),
.B1(n_34),
.B2(n_93),
.Y(n_199)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_15),
.A2(n_56),
.B1(n_58),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_15),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_15),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_15),
.A2(n_28),
.B1(n_34),
.B2(n_67),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_15),
.A2(n_43),
.B1(n_44),
.B2(n_67),
.Y(n_219)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_17),
.A2(n_43),
.B1(n_44),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_17),
.A2(n_28),
.B1(n_34),
.B2(n_51),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_17),
.A2(n_51),
.B1(n_63),
.B2(n_64),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_122),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_102),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_22),
.B(n_102),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_80),
.C(n_96),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_23),
.B(n_96),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_52),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_53),
.C(n_68),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_25),
.B(n_39),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_26),
.A2(n_36),
.B1(n_37),
.B2(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_26),
.A2(n_36),
.B(n_98),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_26),
.A2(n_36),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_26),
.A2(n_192),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_26),
.A2(n_36),
.B1(n_187),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_27),
.A2(n_30),
.B1(n_89),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_27),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_28),
.B(n_48),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_28),
.B(n_205),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g200 ( 
.A(n_30),
.Y(n_200)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_34),
.A2(n_44),
.A3(n_47),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_36),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_36),
.B(n_86),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_41),
.A2(n_108),
.B1(n_111),
.B2(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_43),
.A2(n_63),
.A3(n_73),
.B1(n_216),
.B2(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_44),
.B(n_77),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_45),
.A2(n_46),
.B1(n_50),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_45),
.A2(n_46),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_45),
.A2(n_46),
.B1(n_173),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_45),
.A2(n_46),
.B1(n_140),
.B2(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_46),
.B(n_86),
.Y(n_201)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_68),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_59),
.B1(n_62),
.B2(n_66),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_65),
.B(n_86),
.C(n_87),
.Y(n_85)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_58),
.B(n_60),
.Y(n_61)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_59),
.A2(n_62),
.B1(n_66),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_59),
.A2(n_62),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_62),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_73),
.B(n_75),
.C(n_76),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_73),
.Y(n_75)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_64),
.B(n_86),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B1(n_78),
.B2(n_79),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_78),
.B1(n_79),
.B2(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_71),
.A2(n_79),
.B1(n_134),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_76),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_72),
.A2(n_76),
.B1(n_82),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_72),
.A2(n_76),
.B1(n_155),
.B2(n_214),
.Y(n_213)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.C(n_90),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_90),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_84),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_85),
.B(n_88),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_92),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_100),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_120),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_112),
.B2(n_113),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_108),
.A2(n_111),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_114),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_117),
.CI(n_119),
.CON(n_114),
.SN(n_114)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_160),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_143),
.B(n_159),
.Y(n_124)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_141),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_141),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.C(n_130),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_130),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.C(n_138),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_132),
.B1(n_138),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_146),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_151),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_147),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_248),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_150),
.Y(n_248)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_153),
.B(n_235),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_156),
.B(n_158),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_157),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_244),
.B(n_249),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_230),
.B(n_243),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_209),
.B(n_229),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_188),
.B(n_208),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_178),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_168),
.B(n_178),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_183),
.C(n_185),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_184),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_196),
.B(n_207),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_195),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_202),
.B(n_206),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_198),
.B(n_201),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_211),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_222),
.B1(n_227),
.B2(n_228),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_221),
.C(n_228),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_225),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_232),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_239),
.C(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);


endmodule