module real_aes_2015_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_0), .B(n_129), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_1), .A2(n_138), .B(n_143), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_2), .B(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_3), .B(n_145), .Y(n_183) );
INVx1_ASAP7_75t_L g136 ( .A(n_4), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_5), .B(n_145), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_6), .B(n_155), .Y(n_539) );
INVx1_ASAP7_75t_L g519 ( .A(n_7), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g787 ( .A(n_8), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_9), .Y(n_485) );
NAND2xp33_ASAP7_75t_L g172 ( .A(n_10), .B(n_147), .Y(n_172) );
INVx2_ASAP7_75t_L g126 ( .A(n_11), .Y(n_126) );
AOI221x1_ASAP7_75t_L g218 ( .A1(n_12), .A2(n_24), .B1(n_129), .B2(n_138), .C(n_219), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_13), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_14), .B(n_129), .Y(n_168) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_15), .A2(n_166), .B(n_167), .Y(n_165) );
INVx1_ASAP7_75t_L g547 ( .A(n_16), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_17), .B(n_149), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_18), .B(n_145), .Y(n_159) );
AO21x1_ASAP7_75t_L g178 ( .A1(n_19), .A2(n_129), .B(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
INVx1_ASAP7_75t_L g545 ( .A(n_21), .Y(n_545) );
INVx1_ASAP7_75t_SL g467 ( .A(n_22), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_23), .B(n_130), .Y(n_535) );
NAND2x1_ASAP7_75t_L g191 ( .A(n_25), .B(n_145), .Y(n_191) );
AOI33xp33_ASAP7_75t_L g505 ( .A1(n_26), .A2(n_54), .A3(n_450), .B1(n_455), .B2(n_506), .B3(n_507), .Y(n_505) );
NAND2x1_ASAP7_75t_L g210 ( .A(n_27), .B(n_147), .Y(n_210) );
INVx1_ASAP7_75t_L g478 ( .A(n_28), .Y(n_478) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_29), .A2(n_88), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g151 ( .A(n_29), .B(n_88), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_30), .B(n_458), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_31), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_32), .B(n_145), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_33), .B(n_147), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_34), .A2(n_138), .B(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g135 ( .A(n_35), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g139 ( .A(n_35), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g449 ( .A(n_35), .Y(n_449) );
OR2x6_ASAP7_75t_L g109 ( .A(n_36), .B(n_110), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_37), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_38), .B(n_129), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_39), .B(n_458), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_40), .A2(n_124), .B1(n_155), .B2(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_41), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_42), .B(n_130), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_43), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_44), .B(n_147), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_45), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_46), .Y(n_809) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_47), .B(n_166), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_48), .B(n_130), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_49), .A2(n_138), .B(n_209), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_50), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_51), .A2(n_85), .B1(n_800), .B2(n_801), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_51), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_52), .A2(n_80), .B1(n_770), .B2(n_771), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_52), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_53), .B(n_147), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_55), .B(n_130), .Y(n_496) );
INVx1_ASAP7_75t_L g132 ( .A(n_56), .Y(n_132) );
INVx1_ASAP7_75t_L g142 ( .A(n_56), .Y(n_142) );
AND2x2_ASAP7_75t_L g497 ( .A(n_57), .B(n_149), .Y(n_497) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_58), .A2(n_74), .B1(n_447), .B2(n_458), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_59), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_60), .B(n_145), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_61), .B(n_124), .Y(n_487) );
AOI21xp5_ASAP7_75t_SL g446 ( .A1(n_62), .A2(n_447), .B(n_452), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_63), .A2(n_138), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g542 ( .A(n_64), .Y(n_542) );
AO21x1_ASAP7_75t_L g180 ( .A1(n_65), .A2(n_138), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_66), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g495 ( .A(n_67), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_68), .B(n_129), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_69), .A2(n_447), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g203 ( .A(n_70), .B(n_150), .Y(n_203) );
INVx1_ASAP7_75t_L g134 ( .A(n_71), .Y(n_134) );
INVx1_ASAP7_75t_L g140 ( .A(n_71), .Y(n_140) );
AND2x2_ASAP7_75t_L g214 ( .A(n_72), .B(n_123), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_73), .B(n_458), .Y(n_508) );
AND2x2_ASAP7_75t_L g469 ( .A(n_75), .B(n_123), .Y(n_469) );
INVx1_ASAP7_75t_L g543 ( .A(n_76), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_77), .A2(n_447), .B(n_466), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_78), .A2(n_103), .B1(n_780), .B2(n_791), .C1(n_810), .C2(n_814), .Y(n_102) );
OAI22xp5_ASAP7_75t_SL g797 ( .A1(n_78), .A2(n_798), .B1(n_799), .B2(n_802), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_78), .Y(n_802) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_79), .A2(n_447), .B(n_500), .C(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_80), .Y(n_770) );
INVx1_ASAP7_75t_L g112 ( .A(n_81), .Y(n_112) );
AND2x2_ASAP7_75t_L g122 ( .A(n_82), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_83), .B(n_129), .Y(n_161) );
AND2x2_ASAP7_75t_SL g444 ( .A(n_84), .B(n_123), .Y(n_444) );
INVx1_ASAP7_75t_L g800 ( .A(n_85), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_86), .A2(n_447), .B1(n_503), .B2(n_504), .Y(n_502) );
AND2x2_ASAP7_75t_L g179 ( .A(n_87), .B(n_155), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_89), .B(n_147), .Y(n_160) );
AND2x2_ASAP7_75t_L g195 ( .A(n_90), .B(n_123), .Y(n_195) );
INVx1_ASAP7_75t_L g453 ( .A(n_91), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_92), .B(n_145), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_93), .A2(n_768), .B1(n_769), .B2(n_772), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_93), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_94), .A2(n_138), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_95), .B(n_147), .Y(n_220) );
AND2x2_ASAP7_75t_L g509 ( .A(n_96), .B(n_123), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_97), .B(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_98), .A2(n_476), .B(n_477), .C(n_480), .Y(n_475) );
BUFx2_ASAP7_75t_L g788 ( .A(n_99), .Y(n_788) );
BUFx2_ASAP7_75t_SL g818 ( .A(n_99), .Y(n_818) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_100), .A2(n_138), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_101), .B(n_130), .Y(n_456) );
OAI222xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_766), .B1(n_767), .B2(n_773), .C1(n_778), .C2(n_779), .Y(n_103) );
AOI22x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_113), .B1(n_431), .B2(n_434), .Y(n_104) );
INVx3_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx11_ASAP7_75t_R g777 ( .A(n_107), .Y(n_777) );
AND2x6_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .Y(n_107) );
OR2x6_ASAP7_75t_SL g432 ( .A(n_108), .B(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g778 ( .A(n_108), .B(n_109), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_108), .B(n_433), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_109), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_113), .A2(n_114), .B1(n_797), .B2(n_803), .Y(n_796) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx3_ASAP7_75t_L g776 ( .A(n_114), .Y(n_776) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_340), .Y(n_114) );
NOR4xp25_ASAP7_75t_L g115 ( .A(n_116), .B(n_258), .C(n_284), .D(n_324), .Y(n_115) );
OAI211xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_173), .B(n_204), .C(n_244), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_152), .Y(n_118) );
AND2x2_ASAP7_75t_L g411 ( .A(n_119), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_120), .B(n_152), .Y(n_278) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g205 ( .A(n_121), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_121), .B(n_231), .Y(n_230) );
INVx5_ASAP7_75t_L g264 ( .A(n_121), .Y(n_264) );
NOR2x1_ASAP7_75t_SL g306 ( .A(n_121), .B(n_153), .Y(n_306) );
AND2x2_ASAP7_75t_L g362 ( .A(n_121), .B(n_165), .Y(n_362) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_127), .Y(n_121) );
INVx3_ASAP7_75t_L g194 ( .A(n_123), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_123), .A2(n_194), .B1(n_475), .B2(n_481), .Y(n_474) );
INVx4_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_124), .B(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx4f_ASAP7_75t_L g166 ( .A(n_125), .Y(n_166) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_126), .B(n_151), .Y(n_150) );
AND2x4_ASAP7_75t_L g155 ( .A(n_126), .B(n_151), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_137), .B(n_149), .Y(n_127) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_135), .Y(n_129) );
INVx1_ASAP7_75t_L g479 ( .A(n_130), .Y(n_479) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
AND2x6_ASAP7_75t_L g147 ( .A(n_131), .B(n_140), .Y(n_147) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g145 ( .A(n_133), .B(n_142), .Y(n_145) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx5_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_135), .Y(n_480) );
AND2x2_ASAP7_75t_L g141 ( .A(n_136), .B(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_136), .Y(n_460) );
AND2x6_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
BUFx3_ASAP7_75t_L g461 ( .A(n_139), .Y(n_461) );
INVx2_ASAP7_75t_L g451 ( .A(n_140), .Y(n_451) );
AND2x4_ASAP7_75t_L g447 ( .A(n_141), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g455 ( .A(n_142), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_146), .B(n_148), .Y(n_143) );
INVxp67_ASAP7_75t_L g548 ( .A(n_145), .Y(n_548) );
INVxp67_ASAP7_75t_L g546 ( .A(n_147), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_148), .A2(n_159), .B(n_160), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_148), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_148), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_148), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_148), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_148), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_148), .A2(n_220), .B(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_148), .A2(n_453), .B(n_454), .C(n_456), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_SL g466 ( .A1(n_148), .A2(n_454), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_148), .A2(n_454), .B(n_495), .C(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g503 ( .A(n_148), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_148), .A2(n_454), .B(n_519), .C(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_148), .A2(n_535), .B(n_536), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_148), .B(n_155), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_149), .Y(n_213) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_149), .A2(n_218), .B(n_222), .Y(n_217) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_149), .A2(n_218), .B(n_222), .Y(n_257) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_164), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_153), .B(n_165), .Y(n_234) );
AND2x2_ASAP7_75t_L g295 ( .A(n_153), .B(n_264), .Y(n_295) );
AO21x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_162), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_154), .B(n_163), .Y(n_162) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_154), .A2(n_156), .B(n_162), .Y(n_248) );
INVx1_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_155), .A2(n_168), .B(n_169), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_155), .B(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_155), .A2(n_446), .B(n_457), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_161), .Y(n_156) );
AND2x2_ASAP7_75t_L g307 ( .A(n_164), .B(n_231), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_164), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g351 ( .A(n_164), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g384 ( .A(n_164), .B(n_205), .Y(n_384) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g228 ( .A(n_165), .Y(n_228) );
AND2x2_ASAP7_75t_L g261 ( .A(n_165), .B(n_262), .Y(n_261) );
BUFx3_ASAP7_75t_L g296 ( .A(n_165), .Y(n_296) );
OR2x2_ASAP7_75t_L g372 ( .A(n_165), .B(n_231), .Y(n_372) );
INVx2_ASAP7_75t_SL g500 ( .A(n_166), .Y(n_500) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_166), .A2(n_517), .B(n_521), .Y(n_516) );
INVx1_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_186), .Y(n_174) );
AOI211x1_ASAP7_75t_SL g301 ( .A1(n_175), .A2(n_293), .B(n_302), .C(n_304), .Y(n_301) );
AND2x2_ASAP7_75t_SL g346 ( .A(n_175), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_175), .B(n_344), .Y(n_391) );
BUFx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g241 ( .A(n_176), .Y(n_241) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g216 ( .A(n_177), .Y(n_216) );
OAI21x1_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_180), .B(n_184), .Y(n_177) );
INVx1_ASAP7_75t_L g185 ( .A(n_179), .Y(n_185) );
AOI322xp5_ASAP7_75t_L g204 ( .A1(n_186), .A2(n_205), .A3(n_215), .B1(n_223), .B2(n_226), .C1(n_232), .C2(n_235), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_186), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_196), .Y(n_186) );
INVx2_ASAP7_75t_L g239 ( .A(n_187), .Y(n_239) );
INVxp67_ASAP7_75t_L g281 ( .A(n_187), .Y(n_281) );
BUFx3_ASAP7_75t_L g345 ( .A(n_187), .Y(n_345) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_194), .B(n_195), .Y(n_187) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_188), .A2(n_194), .B(n_195), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_193), .Y(n_188) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_194), .A2(n_197), .B(n_203), .Y(n_196) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_194), .A2(n_197), .B(n_203), .Y(n_243) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_194), .A2(n_491), .B(n_497), .Y(n_490) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_194), .A2(n_491), .B(n_497), .Y(n_513) );
INVx2_ASAP7_75t_L g254 ( .A(n_196), .Y(n_254) );
AND2x2_ASAP7_75t_L g303 ( .A(n_196), .B(n_217), .Y(n_303) );
AND2x2_ASAP7_75t_L g347 ( .A(n_196), .B(n_256), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_198), .B(n_202), .Y(n_197) );
AND2x2_ASAP7_75t_L g232 ( .A(n_205), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_205), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_SL g426 ( .A(n_205), .B(n_261), .Y(n_426) );
INVx4_ASAP7_75t_L g231 ( .A(n_206), .Y(n_231) );
AND2x2_ASAP7_75t_L g263 ( .A(n_206), .B(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_206), .Y(n_316) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_213), .B(n_214), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_212), .Y(n_207) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_213), .A2(n_463), .B(n_469), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_215), .B(n_300), .Y(n_325) );
INVx1_ASAP7_75t_SL g364 ( .A(n_215), .Y(n_364) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
AND2x4_ASAP7_75t_L g255 ( .A(n_216), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_216), .B(n_254), .Y(n_323) );
AND2x2_ASAP7_75t_L g375 ( .A(n_216), .B(n_225), .Y(n_375) );
OR2x2_ASAP7_75t_L g399 ( .A(n_216), .B(n_217), .Y(n_399) );
AND2x2_ASAP7_75t_L g223 ( .A(n_217), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g273 ( .A(n_217), .B(n_254), .Y(n_273) );
AND2x2_ASAP7_75t_SL g329 ( .A(n_217), .B(n_241), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_223), .B(n_336), .Y(n_353) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
BUFx2_ASAP7_75t_L g288 ( .A(n_225), .Y(n_288) );
AND2x4_ASAP7_75t_SL g328 ( .A(n_225), .B(n_242), .Y(n_328) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
OR2x2_ASAP7_75t_L g276 ( .A(n_227), .B(n_230), .Y(n_276) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g245 ( .A(n_228), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g393 ( .A(n_228), .B(n_306), .Y(n_393) );
AND2x2_ASAP7_75t_L g409 ( .A(n_228), .B(n_263), .Y(n_409) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AOI311xp33_ASAP7_75t_L g379 ( .A1(n_230), .A2(n_318), .A3(n_380), .B(n_382), .C(n_389), .Y(n_379) );
AND2x4_ASAP7_75t_L g246 ( .A(n_231), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g250 ( .A(n_231), .Y(n_250) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_231), .B(n_264), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_231), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g363 ( .A(n_231), .B(n_350), .Y(n_363) );
AND2x2_ASAP7_75t_L g249 ( .A(n_233), .B(n_250), .Y(n_249) );
INVxp67_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
INVxp67_ASAP7_75t_SL g267 ( .A(n_234), .Y(n_267) );
OR2x2_ASAP7_75t_L g356 ( .A(n_234), .B(n_320), .Y(n_356) );
INVx1_ASAP7_75t_L g412 ( .A(n_234), .Y(n_412) );
INVx1_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_240), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g321 ( .A(n_238), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g335 ( .A(n_238), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g410 ( .A(n_238), .B(n_283), .Y(n_410) );
BUFx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g253 ( .A(n_239), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g272 ( .A(n_239), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g334 ( .A(n_240), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_240), .A2(n_390), .B1(n_391), .B2(n_392), .Y(n_389) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
AND2x2_ASAP7_75t_L g283 ( .A(n_241), .B(n_254), .Y(n_283) );
AND2x4_ASAP7_75t_L g336 ( .A(n_241), .B(n_243), .Y(n_336) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OAI21xp33_ASAP7_75t_SL g244 ( .A1(n_245), .A2(n_249), .B(n_251), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_245), .A2(n_331), .B1(n_335), .B2(n_337), .Y(n_330) );
AND2x2_ASAP7_75t_SL g290 ( .A(n_246), .B(n_264), .Y(n_290) );
INVx2_ASAP7_75t_L g352 ( .A(n_246), .Y(n_352) );
AND2x2_ASAP7_75t_L g366 ( .A(n_246), .B(n_362), .Y(n_366) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g262 ( .A(n_248), .Y(n_262) );
INVx1_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
INVx1_ASAP7_75t_L g266 ( .A(n_250), .Y(n_266) );
AND3x2_ASAP7_75t_L g294 ( .A(n_250), .B(n_295), .C(n_296), .Y(n_294) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx1_ASAP7_75t_L g358 ( .A(n_253), .Y(n_358) );
AND2x2_ASAP7_75t_L g286 ( .A(n_255), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g357 ( .A(n_255), .B(n_358), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_255), .A2(n_369), .B1(n_373), .B2(n_376), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_255), .B(n_403), .Y(n_407) );
BUFx2_ASAP7_75t_L g298 ( .A(n_256), .Y(n_298) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g269 ( .A(n_257), .Y(n_269) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_257), .Y(n_388) );
OAI221xp5_ASAP7_75t_SL g258 ( .A1(n_259), .A2(n_268), .B1(n_270), .B2(n_271), .C(n_274), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_265), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g350 ( .A(n_262), .Y(n_350) );
INVx2_ASAP7_75t_SL g339 ( .A(n_263), .Y(n_339) );
AND2x2_ASAP7_75t_L g421 ( .A(n_263), .B(n_288), .Y(n_421) );
INVx4_ASAP7_75t_L g312 ( .A(n_264), .Y(n_312) );
INVx1_ASAP7_75t_L g270 ( .A(n_265), .Y(n_270) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AND2x4_ASAP7_75t_L g381 ( .A(n_269), .B(n_336), .Y(n_381) );
INVx1_ASAP7_75t_SL g420 ( .A(n_269), .Y(n_420) );
AND2x2_ASAP7_75t_L g425 ( .A(n_269), .B(n_328), .Y(n_425) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g367 ( .A(n_273), .Y(n_367) );
OAI21xp5_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_277), .B(n_279), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g300 ( .A(n_281), .Y(n_300) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g297 ( .A(n_283), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g387 ( .A(n_283), .B(n_388), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_289), .B(n_291), .C(n_308), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g380 ( .A(n_287), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_288), .B(n_303), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_288), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g413 ( .A(n_288), .B(n_336), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g324 ( .A1(n_289), .A2(n_313), .B1(n_325), .B2(n_326), .C(n_330), .Y(n_324) );
INVx3_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g395 ( .A(n_290), .B(n_296), .Y(n_395) );
OAI32xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_297), .A3(n_299), .B1(n_301), .B2(n_305), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_295), .Y(n_385) );
INVx2_ASAP7_75t_L g318 ( .A(n_296), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g427 ( .A1(n_296), .A2(n_348), .B(n_428), .C(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
OR2x2_ASAP7_75t_L g429 ( .A(n_298), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_302), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g390 ( .A(n_305), .Y(n_390) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g371 ( .A(n_306), .Y(n_371) );
OAI21xp33_ASAP7_75t_SL g308 ( .A1(n_309), .A2(n_317), .B(n_321), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
OR2x2_ASAP7_75t_L g348 ( .A(n_311), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_312), .B(n_315), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_314), .A2(n_346), .B1(n_415), .B2(n_418), .C(n_422), .Y(n_414) );
INVx2_ASAP7_75t_L g417 ( .A(n_314), .Y(n_417) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
OR2x2_ASAP7_75t_L g338 ( .A(n_318), .B(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g405 ( .A(n_318), .B(n_363), .Y(n_405) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVxp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g403 ( .A(n_328), .Y(n_403) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_336), .B(n_366), .Y(n_423) );
INVx2_ASAP7_75t_L g430 ( .A(n_336), .Y(n_430) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_338), .A2(n_401), .B1(n_404), .B2(n_406), .C(n_408), .Y(n_400) );
AND5x1_ASAP7_75t_L g340 ( .A(n_341), .B(n_379), .C(n_394), .D(n_414), .E(n_424), .Y(n_340) );
NOR2xp33_ASAP7_75t_SL g341 ( .A(n_342), .B(n_359), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_348), .B1(n_351), .B2(n_353), .C(n_354), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI221xp5_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_364), .B1(n_365), .B2(n_367), .C(n_368), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_364), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
OR2x2_ASAP7_75t_L g377 ( .A(n_372), .B(n_378), .Y(n_377) );
CKINVDCx16_ASAP7_75t_R g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B(n_386), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_400), .Y(n_394) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_411), .B2(n_413), .Y(n_408) );
O2A1O1Ixp33_ASAP7_75t_L g424 ( .A1(n_410), .A2(n_425), .B(n_426), .C(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g428 ( .A(n_421), .Y(n_428) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g775 ( .A(n_431), .Y(n_775) );
CKINVDCx11_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
OAI22x1_ASAP7_75t_L g774 ( .A1(n_434), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_774) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
AND3x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_656), .C(n_719), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_620), .Y(n_437) );
NOR3xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_561), .C(n_590), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_440), .B(n_550), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_470), .B1(n_510), .B2(n_522), .Y(n_440) );
NAND2x1_ASAP7_75t_L g705 ( .A(n_441), .B(n_551), .Y(n_705) );
INVx2_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_462), .Y(n_442) );
INVx2_ASAP7_75t_L g524 ( .A(n_443), .Y(n_524) );
INVx4_ASAP7_75t_L g566 ( .A(n_443), .Y(n_566) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_443), .Y(n_586) );
AND2x4_ASAP7_75t_L g597 ( .A(n_443), .B(n_565), .Y(n_597) );
AND2x2_ASAP7_75t_L g603 ( .A(n_443), .B(n_527), .Y(n_603) );
NOR2x1_ASAP7_75t_SL g733 ( .A(n_443), .B(n_538), .Y(n_733) );
OR2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVxp67_ASAP7_75t_L g486 ( .A(n_447), .Y(n_486) );
NOR2x1p5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x6_ASAP7_75t_L g454 ( .A(n_451), .B(n_455), .Y(n_454) );
INVxp67_ASAP7_75t_L g476 ( .A(n_454), .Y(n_476) );
INVx2_ASAP7_75t_L g537 ( .A(n_454), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_454), .A2(n_479), .B1(n_542), .B2(n_543), .Y(n_541) );
AND2x2_ASAP7_75t_L g459 ( .A(n_455), .B(n_460), .Y(n_459) );
INVxp33_ASAP7_75t_L g506 ( .A(n_455), .Y(n_506) );
INVx1_ASAP7_75t_L g488 ( .A(n_458), .Y(n_488) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g530 ( .A(n_459), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_461), .Y(n_531) );
INVx2_ASAP7_75t_L g569 ( .A(n_462), .Y(n_569) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_462), .Y(n_583) );
INVx1_ASAP7_75t_L g594 ( .A(n_462), .Y(n_594) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_462), .Y(n_606) );
AND2x2_ASAP7_75t_L g638 ( .A(n_462), .B(n_538), .Y(n_638) );
AND2x2_ASAP7_75t_L g670 ( .A(n_462), .B(n_554), .Y(n_670) );
INVx1_ASAP7_75t_L g677 ( .A(n_462), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_489), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g619 ( .A(n_472), .B(n_558), .Y(n_619) );
INVx2_ASAP7_75t_L g693 ( .A(n_472), .Y(n_693) );
AND2x2_ASAP7_75t_L g716 ( .A(n_472), .B(n_489), .Y(n_716) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_473), .B(n_513), .Y(n_557) );
INVx2_ASAP7_75t_L g578 ( .A(n_473), .Y(n_578) );
AND2x4_ASAP7_75t_L g600 ( .A(n_473), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g635 ( .A(n_473), .Y(n_635) );
AND2x2_ASAP7_75t_L g712 ( .A(n_473), .B(n_516), .Y(n_712) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g683 ( .A(n_489), .Y(n_683) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_498), .Y(n_489) );
NOR2xp67_ASAP7_75t_L g608 ( .A(n_490), .B(n_578), .Y(n_608) );
AND2x2_ASAP7_75t_L g613 ( .A(n_490), .B(n_578), .Y(n_613) );
INVx2_ASAP7_75t_L g626 ( .A(n_490), .Y(n_626) );
NOR2x1_ASAP7_75t_L g674 ( .A(n_490), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
AND2x4_ASAP7_75t_L g599 ( .A(n_498), .B(n_512), .Y(n_599) );
AND2x2_ASAP7_75t_L g614 ( .A(n_498), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g667 ( .A(n_498), .Y(n_667) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_499), .B(n_516), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_499), .B(n_513), .Y(n_671) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B(n_509), .Y(n_499) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_500), .A2(n_501), .B(n_509), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_502), .B(n_508), .Y(n_501) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVxp33_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .Y(n_511) );
INVx3_ASAP7_75t_L g575 ( .A(n_512), .Y(n_575) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_513), .Y(n_573) );
AND2x2_ASAP7_75t_L g742 ( .A(n_513), .B(n_743), .Y(n_742) );
INVx3_ASAP7_75t_L g630 ( .A(n_514), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_514), .B(n_667), .Y(n_762) );
BUFx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g577 ( .A(n_515), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x4_ASAP7_75t_L g558 ( .A(n_516), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g601 ( .A(n_516), .Y(n_601) );
INVxp67_ASAP7_75t_L g615 ( .A(n_516), .Y(n_615) );
INVx1_ASAP7_75t_L g675 ( .A(n_516), .Y(n_675) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_516), .Y(n_743) );
INVx1_ASAP7_75t_L g727 ( .A(n_522), .Y(n_727) );
NOR2x1_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_523), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g681 ( .A(n_524), .B(n_553), .Y(n_681) );
OR2x2_ASAP7_75t_L g717 ( .A(n_525), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g699 ( .A(n_526), .B(n_677), .Y(n_699) );
AND2x2_ASAP7_75t_L g751 ( .A(n_526), .B(n_586), .Y(n_751) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_538), .Y(n_526) );
AND2x4_ASAP7_75t_L g553 ( .A(n_527), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g565 ( .A(n_527), .Y(n_565) );
INVx2_ASAP7_75t_L g582 ( .A(n_527), .Y(n_582) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_527), .Y(n_760) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
NOR3xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .C(n_532), .Y(n_529) );
INVx3_ASAP7_75t_L g554 ( .A(n_538), .Y(n_554) );
INVx2_ASAP7_75t_L g648 ( .A(n_538), .Y(n_648) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_544), .B(n_549), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B1(n_547), .B2(n_548), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_555), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_552), .B(n_628), .Y(n_645) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_552), .B(n_566), .Y(n_687) );
INVx4_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_553), .B(n_628), .Y(n_765) );
AND2x2_ASAP7_75t_L g581 ( .A(n_554), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g595 ( .A(n_554), .Y(n_595) );
AOI22xp5_ASAP7_75t_SL g643 ( .A1(n_555), .A2(n_644), .B1(n_645), .B2(n_646), .Y(n_643) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g640 ( .A(n_556), .B(n_614), .Y(n_640) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g701 ( .A(n_557), .B(n_589), .Y(n_701) );
AND2x2_ASAP7_75t_L g571 ( .A(n_558), .B(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g607 ( .A(n_558), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g703 ( .A(n_558), .B(n_693), .Y(n_703) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g625 ( .A(n_560), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g651 ( .A(n_560), .Y(n_651) );
AND2x2_ASAP7_75t_L g741 ( .A(n_560), .B(n_578), .Y(n_741) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_570), .B1(n_574), .B2(n_579), .C(n_584), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
INVx1_ASAP7_75t_L g642 ( .A(n_564), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_564), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_564), .B(n_638), .Y(n_757) );
AND2x4_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NOR2xp67_ASAP7_75t_SL g610 ( .A(n_566), .B(n_611), .Y(n_610) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_566), .Y(n_623) );
OR2x2_ASAP7_75t_L g707 ( .A(n_566), .B(n_708), .Y(n_707) );
AND2x4_ASAP7_75t_SL g759 ( .A(n_566), .B(n_760), .Y(n_759) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx3_ASAP7_75t_L g628 ( .A(n_568), .Y(n_628) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_569), .Y(n_718) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AOI221x1_ASAP7_75t_L g658 ( .A1(n_571), .A2(n_659), .B1(n_661), .B2(n_664), .C(n_668), .Y(n_658) );
AND2x2_ASAP7_75t_L g644 ( .A(n_572), .B(n_600), .Y(n_644) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AND2x2_ASAP7_75t_L g587 ( .A(n_575), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_575), .B(n_577), .Y(n_714) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
AND2x2_ASAP7_75t_SL g585 ( .A(n_581), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_581), .B(n_594), .Y(n_611) );
INVx2_ASAP7_75t_L g618 ( .A(n_581), .Y(n_618) );
INVx1_ASAP7_75t_L g663 ( .A(n_582), .Y(n_663) );
BUFx2_ASAP7_75t_L g752 ( .A(n_583), .Y(n_752) );
NAND2xp33_ASAP7_75t_SL g584 ( .A(n_585), .B(n_587), .Y(n_584) );
OR2x6_ASAP7_75t_L g617 ( .A(n_586), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g698 ( .A(n_586), .B(n_638), .Y(n_698) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_609), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_598), .B1(n_602), .B2(n_607), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
AND2x2_ASAP7_75t_SL g655 ( .A(n_593), .B(n_597), .Y(n_655) );
AND2x4_ASAP7_75t_L g661 ( .A(n_593), .B(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_SL g593 ( .A(n_594), .B(n_595), .Y(n_593) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_594), .Y(n_686) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_597), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_597), .B(n_628), .Y(n_660) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_597), .Y(n_744) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g691 ( .A(n_599), .B(n_692), .Y(n_691) );
INVx3_ASAP7_75t_L g652 ( .A(n_600), .Y(n_652) );
NAND2x1_ASAP7_75t_SL g696 ( .A(n_600), .B(n_651), .Y(n_696) );
AND2x2_ASAP7_75t_L g730 ( .A(n_600), .B(n_625), .Y(n_730) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B1(n_616), .B2(n_619), .Y(n_609) );
BUFx2_ASAP7_75t_L g725 ( .A(n_611), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_612), .A2(n_681), .B1(n_755), .B2(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_613), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g633 ( .A(n_614), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g749 ( .A(n_618), .B(n_750), .C(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g653 ( .A(n_619), .Y(n_653) );
AOI211x1_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_629), .B(n_631), .C(n_649), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_624), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
AND2x2_ASAP7_75t_L g711 ( .A(n_625), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_625), .B(n_692), .Y(n_723) );
AND2x2_ASAP7_75t_L g755 ( .A(n_625), .B(n_693), .Y(n_755) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g736 ( .A(n_628), .Y(n_736) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g665 ( .A(n_630), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_643), .Y(n_631) );
AOI22xp5_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_636), .B1(n_639), .B2(n_641), .Y(n_632) );
BUFx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g673 ( .A(n_635), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g688 ( .A(n_635), .Y(n_688) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_SL g758 ( .A(n_638), .B(n_759), .Y(n_758) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g694 ( .A(n_647), .B(n_677), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B(n_654), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_651), .B(n_673), .Y(n_748) );
OR2x2_ASAP7_75t_L g726 ( .A(n_652), .B(n_671), .Y(n_726) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND3x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_678), .C(n_702), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_661), .A2(n_691), .B1(n_694), .B2(n_695), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_662), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_SL g735 ( .A(n_662), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_662), .B(n_736), .Y(n_739) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI222xp33_ASAP7_75t_L g722 ( .A1(n_666), .A2(n_723), .B1(n_724), .B2(n_725), .C1(n_726), .C2(n_727), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B1(n_672), .B2(n_676), .Y(n_668) );
INVx1_ASAP7_75t_SL g708 ( .A(n_670), .Y(n_708) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g745 ( .A(n_674), .B(n_741), .Y(n_745) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_689), .Y(n_678) );
AOI21xp5_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_682), .B(n_688), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_697), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_696), .B(n_710), .Y(n_709) );
OAI21xp5_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_699), .B(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g724 ( .A(n_699), .Y(n_724) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_706), .B2(n_709), .C(n_713), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
NAND3x1_ASAP7_75t_L g720 ( .A(n_721), .B(n_746), .C(n_753), .Y(n_720) );
NOR2x1_ASAP7_75t_L g721 ( .A(n_722), .B(n_728), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_737), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_730), .B(n_731), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_732), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_740), .B1(n_744), .B2(n_745), .Y(n_737) );
AND2x4_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_747), .B(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_763), .Y(n_753) );
AOI22xp5_ASAP7_75t_SL g754 ( .A1(n_755), .A2(n_756), .B1(n_758), .B2(n_761), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVxp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g772 ( .A(n_769), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_789), .Y(n_782) );
INVxp67_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_SL g784 ( .A(n_785), .B(n_788), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_SL g813 ( .A(n_786), .B(n_788), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g815 ( .A1(n_786), .A2(n_816), .B(n_819), .Y(n_815) );
INVx1_ASAP7_75t_SL g794 ( .A(n_789), .Y(n_794) );
BUFx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
BUFx3_ASAP7_75t_L g808 ( .A(n_790), .Y(n_808) );
BUFx2_ASAP7_75t_L g820 ( .A(n_790), .Y(n_820) );
INVxp67_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .B(n_804), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g803 ( .A(n_797), .Y(n_803) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NOR2xp33_ASAP7_75t_SL g804 ( .A(n_805), .B(n_809), .Y(n_804) );
INVx1_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
BUFx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
CKINVDCx9p33_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
CKINVDCx11_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
CKINVDCx8_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
endmodule