module real_jpeg_24563_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_1),
.A2(n_41),
.B1(n_45),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_1),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_2),
.A2(n_41),
.B1(n_45),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_6),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_6),
.A2(n_27),
.B1(n_37),
.B2(n_97),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_6),
.A2(n_41),
.B1(n_45),
.B2(n_97),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_7),
.A2(n_41),
.B1(n_45),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_46),
.B1(n_55),
.B2(n_56),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_11),
.A2(n_27),
.B1(n_37),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_11),
.A2(n_31),
.B1(n_66),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_66),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_11),
.A2(n_41),
.B1(n_45),
.B2(n_66),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_13),
.A2(n_32),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_13),
.A2(n_27),
.B1(n_37),
.B2(n_71),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_71),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_13),
.A2(n_41),
.B1(n_45),
.B2(n_71),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_14),
.A2(n_27),
.B1(n_37),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_14),
.A2(n_32),
.B1(n_36),
.B2(n_63),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_14),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_14),
.A2(n_41),
.B1(n_45),
.B2(n_63),
.Y(n_197)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_15),
.B(n_74),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_15),
.B(n_56),
.C(n_58),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_15),
.A2(n_27),
.B1(n_33),
.B2(n_37),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_15),
.B(n_67),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_15),
.A2(n_33),
.B1(n_55),
.B2(n_56),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_15),
.B(n_41),
.C(n_93),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_15),
.A2(n_40),
.B(n_198),
.Y(n_228)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_16),
.Y(n_117)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_16),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_135),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_109),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_21),
.B(n_109),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_82),
.C(n_99),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_22),
.B(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_23),
.B(n_52),
.C(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_30),
.C(n_34),
.Y(n_25)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_26),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_26),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_81)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_27),
.A2(n_37),
.B1(n_58),
.B2(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_27),
.B(n_163),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_30),
.A2(n_80),
.B(n_108),
.Y(n_107)
);

HAxp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_33),
.CON(n_30),
.SN(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_33),
.B(n_95),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_33),
.B(n_226),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_36),
.C(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_38),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_39),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_40),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_40),
.A2(n_85),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_40),
.A2(n_44),
.B1(n_48),
.B2(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_40),
.B(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_40),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_41),
.A2(n_45),
.B1(n_93),
.B2(n_94),
.Y(n_95)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_45),
.B(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_48),
.Y(n_166)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_48),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_68),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_61),
.B(n_64),
.Y(n_52)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_53),
.A2(n_64),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_54),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_54),
.A2(n_133),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_56),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_56),
.B(n_207),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_67),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_65),
.B(n_106),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B(n_75),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_70),
.A2(n_74),
.B1(n_80),
.B2(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_99),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_89),
.Y(n_134)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_90),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_90),
.A2(n_186),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_91),
.A2(n_121),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_96),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_95),
.A2(n_102),
.B(n_171),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.C(n_107),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_101),
.B1(n_104),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_103),
.B(n_121),
.Y(n_186)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_105),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_124),
.B2(n_125),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_118),
.B1(n_122),
.B2(n_123),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_114),
.Y(n_122)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_134),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_246),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_157),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_155),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_140),
.B(n_155),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.C(n_148),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_141),
.A2(n_142),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_148),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_180),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_239),
.B(n_245),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_187),
.B(n_238),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_176),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_160),
.B(n_176),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_169),
.C(n_173),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_161),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_164),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B(n_167),
.Y(n_164)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_168),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_169),
.A2(n_173),
.B1(n_174),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_169),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_183),
.C(n_184),
.Y(n_244)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_232),
.B(n_237),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_208),
.B(n_231),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_202),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_202),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_217),
.B(n_230),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_215),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_223),
.B(n_229),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_220),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_236),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_244),
.Y(n_245)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);


endmodule