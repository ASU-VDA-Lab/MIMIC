module fake_jpeg_21497_n_260 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_34),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_26),
.B(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_19),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_17),
.B1(n_27),
.B2(n_24),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_63),
.Y(n_93)
);

AO22x2_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_17),
.B1(n_27),
.B2(n_34),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_40),
.B1(n_39),
.B2(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_34),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_42),
.B1(n_17),
.B2(n_27),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_66),
.B1(n_57),
.B2(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_67),
.B(n_78),
.Y(n_119)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_70),
.Y(n_105)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_76),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_94),
.B1(n_57),
.B2(n_55),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_18),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_90),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_39),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_85),
.Y(n_111)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_86),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_23),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_63),
.B(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_37),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_37),
.B1(n_24),
.B2(n_21),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_72),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_62),
.C(n_55),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_117),
.C(n_77),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_56),
.Y(n_100)
);

AND2x4_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_53),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_109),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_30),
.B(n_22),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_103),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_110),
.B1(n_118),
.B2(n_88),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_32),
.C(n_21),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_29),
.B1(n_22),
.B2(n_31),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_32),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_81),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_31),
.B(n_30),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_28),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_135),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_84),
.B1(n_85),
.B2(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_125),
.B(n_127),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_98),
.CI(n_120),
.CON(n_154),
.SN(n_154)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_139),
.B1(n_114),
.B2(n_104),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_96),
.A2(n_94),
.B1(n_95),
.B2(n_65),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_141),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_78),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_132),
.B(n_134),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_91),
.B1(n_89),
.B2(n_74),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_28),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_65),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_137),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_20),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_74),
.B1(n_70),
.B2(n_69),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_111),
.C(n_100),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_98),
.C(n_104),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_32),
.Y(n_141)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_20),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_146),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_86),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_83),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_114),
.B(n_111),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_130),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_169),
.C(n_174),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_103),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_162),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_101),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_165),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_152),
.B1(n_155),
.B2(n_123),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_109),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_109),
.Y(n_167)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_120),
.C(n_116),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_150),
.B(n_141),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_83),
.C(n_33),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_0),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_143),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_178),
.B(n_136),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

AOI211xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_170),
.B(n_163),
.C(n_155),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_196),
.B(n_172),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_165),
.B1(n_156),
.B2(n_169),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_171),
.B1(n_174),
.B2(n_148),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_130),
.C(n_129),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_194),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_193),
.B(n_160),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_198),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_164),
.B1(n_158),
.B2(n_156),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_210),
.B1(n_215),
.B2(n_216),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_206),
.Y(n_218)
);

AOI221xp5_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_153),
.B1(n_167),
.B2(n_157),
.C(n_154),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_192),
.B(n_194),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_176),
.B(n_168),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_212),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_161),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_211),
.C(n_186),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_189),
.A2(n_176),
.B1(n_154),
.B2(n_162),
.Y(n_210)
);

OAI321xp33_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_33),
.A3(n_16),
.B1(n_15),
.B2(n_3),
.C(n_4),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_217),
.Y(n_221)
);

OAI22x1_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_216)
);

BUFx12_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

AOI31xp33_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_227),
.A3(n_226),
.B(n_223),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_220),
.B(n_224),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_190),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_226),
.C(n_228),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_187),
.B(n_185),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_183),
.C(n_188),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_183),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_188),
.C(n_195),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_211),
.C(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_228),
.C(n_210),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_203),
.B1(n_202),
.B2(n_217),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_218),
.B1(n_221),
.B2(n_225),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_242)
);

INVx11_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_240),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_214),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_215),
.B(n_206),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_249),
.Y(n_253)
);

NAND5xp2_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_233),
.C(n_232),
.D(n_235),
.E(n_240),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_248),
.B1(n_10),
.B2(n_11),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_SL g248 ( 
.A1(n_241),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_9),
.C(n_10),
.Y(n_249)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_238),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_SL g254 ( 
.A(n_250),
.B(n_244),
.C(n_248),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_244),
.C(n_246),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_256),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_253),
.A2(n_248),
.B(n_13),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_250),
.B1(n_251),
.B2(n_14),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_257),
.B(n_14),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_258),
.Y(n_260)
);


endmodule