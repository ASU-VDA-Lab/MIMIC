module fake_jpeg_26126_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_57),
.Y(n_61)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_48),
.B1(n_51),
.B2(n_50),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_5),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_51),
.B1(n_52),
.B2(n_49),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_45),
.B1(n_47),
.B2(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_6),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_82),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_1),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_40),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g98 ( 
.A(n_79),
.Y(n_98)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_87),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_40),
.C(n_4),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_84)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_82),
.B1(n_88),
.B2(n_78),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_89),
.B1(n_19),
.B2(n_20),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_27),
.B1(n_36),
.B2(n_35),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_7),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_91),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_84),
.B(n_22),
.C(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_99),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_105),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_21),
.B(n_24),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_29),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_114),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_95),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_106),
.B1(n_104),
.B2(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_98),
.C(n_83),
.Y(n_119)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_120),
.B1(n_116),
.B2(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_121),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_121),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_31),
.C(n_32),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_127),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_33),
.Y(n_129)
);


endmodule