module fake_netlist_1_6306_n_33 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_6), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_0), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_4), .Y(n_12) );
OAI22xp33_ASAP7_75t_SL g13 ( .A1(n_4), .A2(n_7), .B1(n_2), .B2(n_3), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
A2O1A1Ixp33_ASAP7_75t_L g15 ( .A1(n_9), .A2(n_1), .B(n_2), .C(n_3), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
AND2x2_ASAP7_75t_SL g17 ( .A(n_13), .B(n_1), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_14), .B(n_10), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
CKINVDCx16_ASAP7_75t_R g21 ( .A(n_14), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_16), .Y(n_22) );
INVx5_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
NOR2xp67_ASAP7_75t_L g24 ( .A(n_19), .B(n_5), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_20), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
AOI211xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_24), .B(n_18), .C(n_15), .Y(n_28) );
OAI221xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_23), .B1(n_22), .B2(n_20), .C(n_12), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g30 ( .A(n_29), .B(n_23), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_28), .B(n_23), .Y(n_31) );
XNOR2xp5_ASAP7_75t_L g32 ( .A(n_31), .B(n_17), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_30), .B1(n_5), .B2(n_8), .Y(n_33) );
endmodule