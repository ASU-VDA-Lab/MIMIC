module fake_jpeg_14347_n_58 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_4),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_27),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_9),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_26),
.B(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_16),
.B1(n_10),
.B2(n_11),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_11),
.B1(n_16),
.B2(n_10),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_13),
.B1(n_20),
.B2(n_19),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_26),
.B(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_27),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_40),
.C(n_32),
.Y(n_41)
);

AO22x1_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_25),
.B1(n_19),
.B2(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_39),
.B2(n_34),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_40),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_47),
.C(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_48),
.B1(n_38),
.B2(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_23),
.B1(n_15),
.B2(n_29),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_51),
.B(n_30),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_37),
.C(n_28),
.Y(n_55)
);

OAI321xp33_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_14),
.A3(n_17),
.B1(n_8),
.B2(n_7),
.C(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_55),
.C(n_29),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_29),
.Y(n_58)
);


endmodule