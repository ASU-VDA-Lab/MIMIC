module fake_jpeg_25344_n_168 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_40),
.B1(n_38),
.B2(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_53),
.Y(n_64)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_25),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_30),
.B1(n_15),
.B2(n_23),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_15),
.B1(n_41),
.B2(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_17),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_76),
.B1(n_56),
.B2(n_73),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_75),
.B1(n_44),
.B2(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_72),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_27),
.B(n_26),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_27),
.B(n_26),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_70),
.B(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_44),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_65),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_34),
.B1(n_32),
.B2(n_40),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_34),
.B1(n_18),
.B2(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_80),
.B1(n_85),
.B2(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_90),
.Y(n_97)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_64),
.B1(n_62),
.B2(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_96),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_101),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_108),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_61),
.B1(n_66),
.B2(n_32),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_107),
.A2(n_94),
.B1(n_91),
.B2(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_72),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_48),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_18),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_24),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_79),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_113),
.B(n_31),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_92),
.B(n_77),
.C(n_18),
.D(n_24),
.Y(n_116)
);

AOI221xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_102),
.B1(n_96),
.B2(n_95),
.C(n_108),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_86),
.C(n_93),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_124),
.C(n_106),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_110),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_91),
.B1(n_45),
.B2(n_58),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_123),
.B(n_31),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_29),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_100),
.B(n_31),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_130),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_135),
.B1(n_119),
.B2(n_117),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_129),
.C(n_134),
.Y(n_137)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_132),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_139),
.C(n_143),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_121),
.C(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_142),
.B(n_140),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_115),
.C(n_111),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_SL g144 ( 
.A(n_135),
.B(n_116),
.C(n_11),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_10),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_16),
.B(n_8),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_136),
.B1(n_133),
.B2(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_148),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_130),
.C(n_58),
.Y(n_148)
);

AOI321xp33_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_9),
.A3(n_10),
.B1(n_12),
.B2(n_6),
.C(n_7),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g155 ( 
.A(n_149),
.B(n_151),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_150),
.A2(n_152),
.B(n_8),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_141),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_157),
.Y(n_161)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_156),
.Y(n_159)
);

NOR2xp67_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_16),
.Y(n_158)
);

OAI21x1_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_16),
.B(n_45),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_11),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_160),
.B(n_12),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_156),
.B1(n_155),
.B2(n_7),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_159),
.C(n_2),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_0),
.B(n_2),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_165),
.Y(n_168)
);


endmodule