module fake_jpeg_31459_n_526 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_56),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_9),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_59),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_18),
.B(n_9),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_18),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_72),
.Y(n_105)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_21),
.B(n_8),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_75),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_88),
.Y(n_161)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_37),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_89),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_21),
.B(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_97),
.B(n_101),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_27),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_25),
.B(n_44),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_25),
.Y(n_118)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_38),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_48),
.B1(n_46),
.B2(n_43),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_110),
.A2(n_87),
.B1(n_70),
.B2(n_69),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_78),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_123),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_118),
.B(n_120),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_57),
.B(n_39),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_61),
.B(n_39),
.Y(n_123)
);

BUFx4f_ASAP7_75t_SL g129 ( 
.A(n_56),
.Y(n_129)
);

BUFx16f_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_56),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_143),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_55),
.B(n_28),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_134),
.B(n_160),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_135),
.Y(n_215)
);

NAND2x1_ASAP7_75t_SL g138 ( 
.A(n_82),
.B(n_23),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_138),
.A2(n_164),
.B(n_12),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_74),
.B(n_28),
.Y(n_160)
);

HAxp5_ASAP7_75t_SL g164 ( 
.A(n_81),
.B(n_23),
.CON(n_164),
.SN(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_68),
.B(n_38),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_49),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_109),
.A2(n_100),
.B1(n_91),
.B2(n_90),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_166),
.A2(n_169),
.B1(n_196),
.B2(n_200),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_164),
.A2(n_99),
.B1(n_35),
.B2(n_27),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_105),
.A2(n_63),
.B1(n_83),
.B2(n_76),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_138),
.A2(n_35),
.B1(n_46),
.B2(n_48),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_171),
.A2(n_198),
.B1(n_199),
.B2(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_175),
.B(n_217),
.Y(n_251)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_176),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_31),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_179),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_31),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_151),
.B1(n_124),
.B2(n_111),
.Y(n_224)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx5_ASAP7_75t_SL g238 ( 
.A(n_182),
.Y(n_238)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_130),
.Y(n_185)
);

BUFx2_ASAP7_75t_SL g230 ( 
.A(n_185),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_189),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_115),
.B(n_153),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_195),
.B(n_201),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_115),
.A2(n_64),
.B1(n_62),
.B2(n_58),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_149),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_133),
.A2(n_43),
.B1(n_152),
.B2(n_141),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_131),
.A2(n_29),
.B1(n_51),
.B2(n_40),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_51),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_203),
.A2(n_126),
.B(n_121),
.Y(n_234)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_113),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_206),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_119),
.B(n_31),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_106),
.B(n_49),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_207),
.B(n_211),
.Y(n_236)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_31),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_212),
.Y(n_219)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_137),
.B(n_49),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_159),
.A2(n_29),
.B1(n_40),
.B2(n_49),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_126),
.B1(n_162),
.B2(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_136),
.B(n_49),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_144),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_218),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_181),
.A2(n_111),
.B1(n_151),
.B2(n_124),
.Y(n_220)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_220),
.A2(n_234),
.B(n_240),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_224),
.B(n_243),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_177),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_241),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_181),
.B(n_201),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_187),
.B(n_161),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_150),
.C(n_148),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_172),
.B(n_129),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_257),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_175),
.B(n_159),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_211),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_173),
.A2(n_110),
.B1(n_150),
.B2(n_40),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_255),
.A2(n_218),
.B1(n_185),
.B2(n_212),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_186),
.B(n_29),
.Y(n_257)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_264),
.Y(n_299)
);

INVx6_ASAP7_75t_SL g263 ( 
.A(n_230),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_283),
.Y(n_297)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_205),
.B(n_180),
.C(n_207),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_265),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_266),
.A2(n_274),
.B1(n_238),
.B2(n_248),
.Y(n_314)
);

CKINVDCx12_ASAP7_75t_R g267 ( 
.A(n_231),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_267),
.Y(n_310)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_227),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_270),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_237),
.B(n_195),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_269),
.B(n_281),
.C(n_287),
.Y(n_319)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_271),
.A2(n_280),
.B(n_294),
.Y(n_307)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_273),
.Y(n_303)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_225),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_245),
.A2(n_217),
.B1(n_146),
.B2(n_147),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_278),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_237),
.A2(n_148),
.B1(n_147),
.B2(n_146),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_276),
.A2(n_222),
.B1(n_218),
.B2(n_185),
.Y(n_302)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_186),
.Y(n_279)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_279),
.B(n_40),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_232),
.A2(n_183),
.B(n_170),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_259),
.B(n_194),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_228),
.B(n_202),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_236),
.B(n_208),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_285),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_216),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_286),
.B(n_288),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_167),
.C(n_204),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_210),
.Y(n_288)
);

AND2x6_ASAP7_75t_L g289 ( 
.A(n_240),
.B(n_167),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_289),
.A2(n_248),
.B(n_167),
.Y(n_317)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_291),
.Y(n_311)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_295),
.Y(n_313)
);

CKINVDCx12_ASAP7_75t_R g294 ( 
.A(n_231),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_246),
.B(n_219),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_191),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_248),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_233),
.B(n_232),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_298),
.A2(n_320),
.B(n_327),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_245),
.B1(n_221),
.B2(n_255),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_300),
.A2(n_305),
.B1(n_308),
.B2(n_263),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_317),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_251),
.B1(n_243),
.B2(n_224),
.Y(n_305)
);

OAI32xp33_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_251),
.A3(n_234),
.B1(n_252),
.B2(n_224),
.Y(n_306)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_306),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_224),
.B1(n_222),
.B2(n_239),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_249),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_312),
.C(n_323),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_249),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_314),
.A2(n_315),
.B1(n_318),
.B2(n_326),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_274),
.A2(n_239),
.B1(n_250),
.B2(n_238),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_327),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_266),
.A2(n_238),
.B1(n_125),
.B2(n_190),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_289),
.A2(n_229),
.B(n_256),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_284),
.B(n_247),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_267),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_281),
.B(n_279),
.C(n_269),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_182),
.C(n_192),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_265),
.A2(n_125),
.B1(n_214),
.B2(n_193),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_277),
.B(n_254),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_277),
.A2(n_229),
.B(n_258),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_329),
.A2(n_293),
.B(n_294),
.Y(n_345)
);

OAI32xp33_ASAP7_75t_L g330 ( 
.A1(n_277),
.A2(n_282),
.A3(n_265),
.B1(n_262),
.B2(n_283),
.Y(n_330)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_330),
.Y(n_341)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_317),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_331),
.A2(n_344),
.B(n_345),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_297),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_333),
.B(n_356),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_282),
.Y(n_334)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_334),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_304),
.B(n_270),
.Y(n_335)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_335),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_272),
.Y(n_336)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_336),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_299),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_338),
.Y(n_375)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_301),
.Y(n_342)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_342),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_346),
.A2(n_348),
.B(n_324),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_262),
.Y(n_347)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_329),
.A2(n_273),
.B(n_268),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_349),
.A2(n_363),
.B1(n_324),
.B2(n_306),
.Y(n_376)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_353),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_309),
.B(n_286),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_352),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_316),
.B(n_261),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_303),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_359),
.Y(n_367)
);

OAI22x1_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_275),
.B1(n_242),
.B2(n_292),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_355),
.A2(n_318),
.B1(n_315),
.B2(n_310),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_313),
.B(n_291),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_264),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_357),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_309),
.B(n_292),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_312),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_278),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_308),
.A2(n_253),
.B(n_256),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_362),
.Y(n_382)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_319),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_313),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_321),
.A2(n_326),
.B1(n_314),
.B2(n_300),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_355),
.Y(n_364)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_364),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_337),
.B(n_323),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_379),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_334),
.B(n_310),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_384),
.C(n_356),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_341),
.A2(n_305),
.B1(n_321),
.B2(n_298),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_370),
.A2(n_376),
.B1(n_355),
.B2(n_362),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_371),
.A2(n_385),
.B1(n_343),
.B2(n_346),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_372),
.A2(n_345),
.B(n_332),
.Y(n_404)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_342),
.B(n_323),
.Y(n_377)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_312),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_391),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_307),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_336),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_319),
.C(n_299),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_387),
.C(n_344),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_253),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_383),
.Y(n_406)
);

OAI21xp33_ASAP7_75t_L g384 ( 
.A1(n_333),
.A2(n_322),
.B(n_311),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_341),
.A2(n_311),
.B1(n_322),
.B2(n_302),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_242),
.C(n_188),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_260),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_174),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_395),
.B(n_360),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_417),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_397),
.A2(n_371),
.B1(n_410),
.B2(n_415),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_349),
.C(n_339),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_402),
.C(n_408),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_400),
.B(n_401),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_339),
.C(n_335),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_340),
.B1(n_332),
.B2(n_348),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_403),
.A2(n_412),
.B1(n_385),
.B2(n_394),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_404),
.A2(n_372),
.B(n_367),
.Y(n_432)
);

OAI22x1_ASAP7_75t_SL g405 ( 
.A1(n_364),
.A2(n_363),
.B1(n_331),
.B2(n_346),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_405),
.A2(n_409),
.B1(n_414),
.B2(n_399),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_407),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_338),
.C(n_359),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_389),
.A2(n_357),
.B1(n_343),
.B2(n_353),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_388),
.B(n_235),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_420),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_376),
.A2(n_260),
.B1(n_235),
.B2(n_184),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_415),
.A2(n_422),
.B1(n_394),
.B2(n_390),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_375),
.B(n_260),
.Y(n_416)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_416),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_235),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_176),
.C(n_197),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_379),
.C(n_380),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_382),
.B(n_235),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_215),
.Y(n_421)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_421),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_370),
.A2(n_0),
.B1(n_1),
.B2(n_40),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_393),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_388),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_381),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_398),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_416),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_411),
.Y(n_455)
);

BUFx24_ASAP7_75t_SL g430 ( 
.A(n_414),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_430),
.B(n_418),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_431),
.A2(n_436),
.B1(n_439),
.B2(n_446),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_432),
.B(n_441),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_440),
.C(n_443),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_410),
.Y(n_435)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_435),
.Y(n_449)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_396),
.B(n_369),
.C(n_377),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_398),
.B(n_369),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_378),
.C(n_366),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_401),
.B(n_366),
.C(n_367),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_444),
.B(n_10),
.C(n_3),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_445),
.A2(n_405),
.B1(n_422),
.B2(n_409),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_397),
.A2(n_392),
.B1(n_391),
.B2(n_215),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_448),
.A2(n_431),
.B1(n_436),
.B2(n_427),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_433),
.B(n_437),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_450),
.B(n_452),
.Y(n_467)
);

FAx1_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_402),
.CI(n_411),
.CON(n_451),
.SN(n_451)
);

XNOR2x1_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_454),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_435),
.A2(n_404),
.B(n_392),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_453),
.B(n_457),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_441),
.B(n_417),
.Y(n_454)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_455),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_406),
.Y(n_456)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

NOR3xp33_ASAP7_75t_SL g457 ( 
.A(n_440),
.B(n_418),
.C(n_419),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_460),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_443),
.B(n_8),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_462),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_10),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_426),
.C(n_425),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_465),
.A2(n_458),
.B1(n_449),
.B2(n_448),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_466),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_447),
.B(n_444),
.CI(n_425),
.CON(n_469),
.SN(n_469)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_474),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_470),
.A2(n_471),
.B1(n_464),
.B2(n_454),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_451),
.A2(n_427),
.B1(n_434),
.B2(n_429),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_473),
.B(n_6),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_10),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_0),
.C(n_16),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_7),
.C(n_3),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_457),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_480),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_7),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_7),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_482),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_475),
.B(n_451),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_485),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_478),
.B(n_459),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_479),
.B(n_452),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_490),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_481),
.B(n_447),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_488),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_497),
.C(n_482),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_467),
.B(n_13),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_492),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_482),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_0),
.C(n_6),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_496),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_470),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_466),
.B(n_14),
.C(n_15),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_502),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_477),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_493),
.B(n_468),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_503),
.B(n_506),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_481),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_507),
.B(n_508),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_484),
.A2(n_476),
.B1(n_469),
.B2(n_472),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_499),
.Y(n_510)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_510),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_486),
.C(n_489),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_511),
.A2(n_513),
.B(n_515),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_496),
.C(n_488),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_501),
.B(n_498),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_514),
.A2(n_508),
.B(n_497),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_519),
.C(n_509),
.Y(n_520)
);

AOI211x1_ASAP7_75t_L g519 ( 
.A1(n_512),
.A2(n_469),
.B(n_473),
.C(n_505),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_521),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_490),
.C(n_15),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_522),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_523),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_518),
.B(n_15),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_16),
.B(n_493),
.Y(n_526)
);


endmodule