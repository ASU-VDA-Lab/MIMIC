module fake_jpeg_14513_n_38 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_23),
.B(n_24),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_26),
.C(n_27),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

AND2x6_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_16),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_29),
.C(n_30),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_11),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_35),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_26),
.B1(n_13),
.B2(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_32),
.Y(n_37)
);

AO21x1_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_15),
.B(n_17),
.Y(n_38)
);


endmodule