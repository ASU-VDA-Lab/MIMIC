module fake_ariane_183_n_2192 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2192);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2192;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_967;
wire n_274;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_70),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_120),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_205),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_122),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_147),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_155),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_12),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_40),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_76),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_87),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_202),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_3),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_154),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_66),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_102),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_137),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_158),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_7),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_144),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_124),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_70),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_146),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_157),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_164),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_59),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_177),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_142),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_59),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_208),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_29),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_107),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_203),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_93),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_30),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_159),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_91),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_26),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_4),
.Y(n_265)
);

INVx4_ASAP7_75t_R g266 ( 
.A(n_176),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_163),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_20),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_149),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_76),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_108),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_27),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_152),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_136),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_50),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_24),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_45),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_170),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_63),
.Y(n_280)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_78),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_62),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_212),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_187),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_105),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_186),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_98),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_145),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_150),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_174),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_119),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_130),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_2),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_72),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_16),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_66),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_166),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_9),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_20),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_220),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_78),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_101),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_40),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_195),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_26),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_94),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_85),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_30),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_199),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_71),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_190),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_61),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_189),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_172),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_77),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_36),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_143),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_97),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_109),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_115),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_14),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_167),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_22),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_83),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_52),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_179),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_193),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_96),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_95),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_181),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_71),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_54),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_28),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_15),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_43),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_211),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_52),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_88),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_42),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_180),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_51),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_19),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_183),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_117),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_56),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_173),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_99),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_68),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_13),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_161),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_165),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_12),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_111),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_169),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_139),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_65),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_118),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_50),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_39),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_68),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_75),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_19),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_72),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_16),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_61),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_153),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_42),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_218),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_86),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_191),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_21),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_129),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_45),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_23),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_38),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_135),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_213),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_56),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_18),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_69),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_81),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_92),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_127),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_15),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_38),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_162),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_214),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_33),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_126),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_17),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_182),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_21),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_104),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_160),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_192),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_63),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_0),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_55),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_201),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_106),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_140),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_215),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_128),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_110),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_10),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_133),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_219),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_77),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_49),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_89),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_3),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_206),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_51),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_39),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_17),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_134),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_112),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_82),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_131),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_65),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_25),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_5),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_11),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_67),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_9),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_22),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_185),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_46),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_24),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_13),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_23),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_125),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_32),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_113),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_151),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_216),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_80),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_254),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_281),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_235),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_281),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_243),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_281),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_257),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_279),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_298),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_345),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_281),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_281),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_281),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_281),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_413),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_385),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_418),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_281),
.Y(n_456)
);

INVxp33_ASAP7_75t_SL g457 ( 
.A(n_306),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_385),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_301),
.B(n_321),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_230),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_281),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_242),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_301),
.B(n_0),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_251),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_343),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_221),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_270),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_221),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_303),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_273),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_224),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_224),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_238),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_234),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_276),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_299),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_283),
.B(n_1),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_234),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_372),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_299),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_321),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_278),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_280),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_223),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_239),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_239),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_305),
.Y(n_487)
);

INVxp33_ASAP7_75t_SL g488 ( 
.A(n_296),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_250),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_223),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_236),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_297),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_246),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_265),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_300),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_250),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_309),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_304),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_261),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_261),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_236),
.Y(n_501)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_318),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_283),
.B(n_1),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_353),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_271),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_362),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_256),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_271),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_311),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_275),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_285),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_256),
.Y(n_512)
);

BUFx6f_ASAP7_75t_SL g513 ( 
.A(n_396),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_376),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_263),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_386),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_313),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_263),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_275),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_R g520 ( 
.A(n_222),
.B(n_90),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_286),
.B(n_2),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_285),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_286),
.B(n_5),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_305),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_316),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_288),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_322),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_288),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_324),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_332),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_334),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_335),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_291),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_336),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_338),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_291),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_293),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_340),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_349),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_350),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_359),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_293),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_360),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_231),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_308),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_308),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_312),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_363),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_364),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_303),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_312),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_314),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_314),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_366),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_319),
.Y(n_555)
);

NOR2xp67_ASAP7_75t_L g556 ( 
.A(n_379),
.B(n_6),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_319),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_320),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_440),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_443),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_440),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_454),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_473),
.A2(n_268),
.B1(n_438),
.B2(n_295),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_442),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_442),
.Y(n_565)
);

INVx6_ASAP7_75t_L g566 ( 
.A(n_511),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_459),
.B(n_247),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_445),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_511),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_444),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_511),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_480),
.B(n_264),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_466),
.B(n_231),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_487),
.B(n_320),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_469),
.B(n_396),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_446),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_444),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_449),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_449),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_450),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_450),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_447),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_451),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_511),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_476),
.B(n_232),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_487),
.B(n_327),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_448),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_511),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_453),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_522),
.Y(n_590)
);

OAI21x1_ASAP7_75t_L g591 ( 
.A1(n_461),
.A2(n_352),
.B(n_327),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_522),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_451),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_452),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_452),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_522),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_466),
.B(n_260),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_544),
.B(n_232),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_460),
.B(n_396),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_524),
.B(n_352),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_456),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_522),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_455),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_493),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_524),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_468),
.B(n_260),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_461),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_456),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_441),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_522),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_468),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_471),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_481),
.B(n_355),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_471),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_463),
.B(n_294),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_494),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_472),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_544),
.B(n_232),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_472),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_474),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_462),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_474),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_478),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_458),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_490),
.B(n_232),
.Y(n_625)
);

BUFx8_ASAP7_75t_L g626 ( 
.A(n_513),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_478),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_485),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_485),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_497),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_486),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_486),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_489),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_464),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_489),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_496),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_467),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_496),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_SL g639 ( 
.A(n_550),
.B(n_380),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_499),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_499),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_491),
.B(n_294),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_500),
.B(n_355),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_500),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_470),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_504),
.B(n_506),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_505),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_505),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_475),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_482),
.B(n_396),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_508),
.B(n_356),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_483),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_567),
.A2(n_510),
.B1(n_519),
.B2(n_508),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_SL g654 ( 
.A(n_621),
.B(n_513),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_612),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_611),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_567),
.B(n_502),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_635),
.B(n_510),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_L g659 ( 
.A(n_624),
.B(n_523),
.C(n_521),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_611),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_598),
.B(n_618),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_607),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_612),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_607),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_625),
.B(n_356),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_615),
.A2(n_457),
.B1(n_488),
.B2(n_477),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_615),
.B(n_501),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_635),
.B(n_519),
.Y(n_668)
);

INVx6_ASAP7_75t_L g669 ( 
.A(n_626),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_605),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_612),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_635),
.B(n_644),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_612),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_625),
.B(n_370),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_614),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_634),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_612),
.B(n_492),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_607),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_635),
.B(n_513),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_615),
.A2(n_528),
.B1(n_533),
.B2(n_526),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_604),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_607),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_562),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_614),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_598),
.B(n_495),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_619),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_L g687 ( 
.A(n_637),
.B(n_509),
.C(n_498),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_619),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_645),
.B(n_527),
.C(n_517),
.Y(n_689)
);

INVxp33_ASAP7_75t_L g690 ( 
.A(n_562),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_559),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_560),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_612),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_605),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_615),
.A2(n_530),
.B1(n_531),
.B2(n_529),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_618),
.B(n_370),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_605),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_624),
.B(n_563),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_644),
.B(n_526),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_615),
.A2(n_533),
.B1(n_536),
.B2(n_528),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_585),
.A2(n_599),
.B1(n_650),
.B2(n_575),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_622),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_559),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_627),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_620),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_644),
.B(n_536),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_644),
.B(n_532),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_648),
.B(n_537),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_620),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_620),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_620),
.B(n_534),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_627),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_573),
.A2(n_545),
.B1(n_546),
.B2(n_542),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_572),
.B(n_465),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_620),
.B(n_285),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_561),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_561),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_628),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_620),
.B(n_535),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_585),
.A2(n_539),
.B1(n_540),
.B2(n_538),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_649),
.B(n_541),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_632),
.Y(n_722)
);

OR2x6_ASAP7_75t_L g723 ( 
.A(n_563),
.B(n_439),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_648),
.B(n_542),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_564),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_632),
.B(n_543),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_632),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_628),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_631),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_632),
.Y(n_730)
);

INVx6_ASAP7_75t_L g731 ( 
.A(n_626),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_631),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_616),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_572),
.B(n_479),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_573),
.A2(n_547),
.B1(n_551),
.B2(n_546),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_632),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_652),
.B(n_525),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_633),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_633),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_568),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_640),
.B(n_548),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_573),
.A2(n_551),
.B1(n_552),
.B2(n_547),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_564),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_626),
.Y(n_744)
);

AND2x6_ASAP7_75t_L g745 ( 
.A(n_640),
.B(n_373),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_641),
.B(n_549),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_SL g747 ( 
.A(n_626),
.B(n_554),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_641),
.B(n_552),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_632),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_565),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_636),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_617),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_565),
.B(n_553),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_617),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_636),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_642),
.B(n_507),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_617),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_570),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_636),
.B(n_373),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_576),
.B(n_484),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_570),
.B(n_553),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_646),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_577),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_636),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_613),
.A2(n_503),
.B1(n_426),
.B2(n_556),
.Y(n_765)
);

AND3x2_ASAP7_75t_L g766 ( 
.A(n_642),
.B(n_277),
.C(n_264),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_623),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_623),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_636),
.Y(n_769)
);

NOR2x1p5_ASAP7_75t_L g770 ( 
.A(n_582),
.B(n_512),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_623),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_577),
.B(n_555),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_630),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_578),
.Y(n_774)
);

NOR2x1p5_ASAP7_75t_L g775 ( 
.A(n_587),
.B(n_515),
.Y(n_775)
);

CKINVDCx8_ASAP7_75t_R g776 ( 
.A(n_609),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_578),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_579),
.B(n_555),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_629),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_579),
.Y(n_780)
);

NOR2x1p5_ASAP7_75t_L g781 ( 
.A(n_589),
.B(n_518),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_SL g782 ( 
.A(n_643),
.B(n_557),
.Y(n_782)
);

INVx6_ASAP7_75t_L g783 ( 
.A(n_636),
.Y(n_783)
);

BUFx6f_ASAP7_75t_SL g784 ( 
.A(n_573),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_580),
.B(n_378),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_597),
.B(n_557),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_580),
.B(n_581),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_581),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_629),
.Y(n_789)
);

INVx5_ASAP7_75t_L g790 ( 
.A(n_584),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_574),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_583),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_583),
.B(n_558),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_593),
.B(n_378),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_597),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_584),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_597),
.A2(n_558),
.B1(n_606),
.B2(n_629),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_593),
.B(n_388),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_638),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_638),
.Y(n_800)
);

INVx5_ASAP7_75t_L g801 ( 
.A(n_584),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_594),
.B(n_388),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_594),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_595),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_595),
.B(n_237),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_601),
.Y(n_806)
);

AND2x6_ASAP7_75t_L g807 ( 
.A(n_638),
.B(n_392),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_601),
.B(n_392),
.Y(n_808)
);

OAI221xp5_ASAP7_75t_L g809 ( 
.A1(n_653),
.A2(n_406),
.B1(n_277),
.B2(n_282),
.C(n_302),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_791),
.B(n_647),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_741),
.B(n_603),
.C(n_639),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_707),
.B(n_608),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_758),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_665),
.A2(n_520),
.B1(n_647),
.B2(n_643),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_707),
.B(n_647),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_758),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_679),
.B(n_608),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_691),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_657),
.B(n_514),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_690),
.B(n_516),
.Y(n_820)
);

OAI22xp33_ASAP7_75t_L g821 ( 
.A1(n_701),
.A2(n_651),
.B1(n_326),
.B2(n_374),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_679),
.B(n_651),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_680),
.B(n_591),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_661),
.B(n_597),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_665),
.B(n_606),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_667),
.B(n_606),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_665),
.B(n_606),
.Y(n_827)
);

AND2x6_ASAP7_75t_L g828 ( 
.A(n_744),
.B(n_403),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_669),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_760),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_685),
.B(n_646),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_665),
.B(n_574),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_669),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_721),
.B(n_586),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_690),
.B(n_586),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_740),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_665),
.B(n_600),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_737),
.B(n_600),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_674),
.B(n_358),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_691),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_772),
.A2(n_591),
.B(n_302),
.C(n_317),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_680),
.B(n_591),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_700),
.B(n_403),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_674),
.A2(n_326),
.B1(n_374),
.B2(n_430),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_674),
.B(n_325),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_795),
.B(n_420),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_674),
.B(n_325),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_720),
.B(n_382),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_674),
.A2(n_420),
.B1(n_436),
.B2(n_435),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_741),
.B(n_430),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_700),
.B(n_433),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_746),
.B(n_393),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_746),
.B(n_433),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_734),
.B(n_282),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_669),
.B(n_317),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_696),
.B(n_653),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_788),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_696),
.B(n_435),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_696),
.B(n_436),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_756),
.B(n_333),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_667),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_703),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_788),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_703),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_683),
.B(n_333),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_731),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_695),
.B(n_397),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_716),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_696),
.A2(n_384),
.B1(n_390),
.B2(n_437),
.Y(n_869)
);

INVx8_ASAP7_75t_L g870 ( 
.A(n_745),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_696),
.B(n_342),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_667),
.B(n_772),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_795),
.A2(n_398),
.B1(n_399),
.B2(n_409),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_795),
.A2(n_412),
.B1(n_415),
.B2(n_416),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_655),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_733),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_672),
.B(n_384),
.Y(n_877)
);

NAND2xp33_ASAP7_75t_L g878 ( 
.A(n_745),
.B(n_423),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_745),
.A2(n_797),
.B1(n_723),
.B2(n_659),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_793),
.B(n_342),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_744),
.B(n_346),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_656),
.A2(n_424),
.B1(n_427),
.B2(n_429),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_716),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_786),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_745),
.A2(n_390),
.B1(n_351),
.B2(n_305),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_655),
.Y(n_886)
);

NOR2x1p5_ASAP7_75t_L g887 ( 
.A(n_692),
.B(n_431),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_676),
.B(n_714),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_786),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_666),
.B(n_432),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_672),
.B(n_663),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_L g892 ( 
.A(n_745),
.B(n_285),
.Y(n_892)
);

NAND2x1_ASAP7_75t_L g893 ( 
.A(n_783),
.B(n_566),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_687),
.B(n_346),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_670),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_663),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_782),
.A2(n_249),
.B1(n_252),
.B2(n_253),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_717),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_L g899 ( 
.A(n_689),
.B(n_361),
.C(n_357),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_660),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_793),
.B(n_357),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_675),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_677),
.B(n_361),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_684),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_663),
.B(n_272),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_677),
.B(n_365),
.Y(n_906)
);

NOR3x1_ASAP7_75t_L g907 ( 
.A(n_765),
.B(n_368),
.C(n_365),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_686),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_805),
.B(n_368),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_711),
.B(n_375),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_797),
.B(n_375),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_681),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_663),
.B(n_272),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_723),
.A2(n_351),
.B1(n_408),
.B2(n_244),
.Y(n_914)
);

INVx8_ASAP7_75t_L g915 ( 
.A(n_784),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_713),
.B(n_381),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_713),
.B(n_381),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_717),
.Y(n_918)
);

AND2x6_ASAP7_75t_SL g919 ( 
.A(n_723),
.B(n_698),
.Y(n_919)
);

AND2x6_ASAP7_75t_SL g920 ( 
.A(n_698),
.B(n_389),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_694),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_725),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_694),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_782),
.A2(n_240),
.B1(n_227),
.B2(n_226),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_SL g925 ( 
.A(n_692),
.B(n_244),
.Y(n_925)
);

BUFx12f_ASAP7_75t_L g926 ( 
.A(n_676),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_711),
.B(n_389),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_673),
.B(n_289),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_725),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_698),
.A2(n_408),
.B1(n_351),
.B2(n_391),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_673),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_688),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_719),
.B(n_726),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_743),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_770),
.B(n_775),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_784),
.A2(n_408),
.B1(n_434),
.B2(n_419),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_676),
.B(n_391),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_781),
.B(n_406),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_735),
.B(n_410),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_735),
.B(n_410),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_719),
.B(n_414),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_742),
.B(n_414),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_742),
.B(n_419),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_743),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_702),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_704),
.B(n_421),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_750),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_712),
.B(n_421),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_726),
.A2(n_225),
.B1(n_229),
.B2(n_233),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_718),
.B(n_728),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_654),
.A2(n_347),
.B1(n_241),
.B2(n_245),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_802),
.A2(n_425),
.B(n_422),
.C(n_434),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_750),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_729),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_732),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_738),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_763),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_731),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_673),
.B(n_289),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_673),
.B(n_705),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_705),
.B(n_404),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_655),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_705),
.B(n_404),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_747),
.B(n_731),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_776),
.B(n_422),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_763),
.Y(n_966)
);

OR2x2_ASAP7_75t_SL g967 ( 
.A(n_681),
.B(n_425),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_774),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_697),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_722),
.B(n_285),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_739),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_774),
.A2(n_337),
.B1(n_228),
.B2(n_344),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_777),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_722),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_L g975 ( 
.A(n_722),
.B(n_337),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_787),
.A2(n_348),
.B1(n_255),
.B2(n_258),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_658),
.B(n_248),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_722),
.B(n_337),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_896),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_822),
.A2(n_780),
.B(n_777),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_822),
.A2(n_815),
.B(n_817),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_852),
.A2(n_808),
.B(n_802),
.C(n_699),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_817),
.A2(n_792),
.B(n_780),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_838),
.B(n_748),
.Y(n_984)
);

AO21x1_ASAP7_75t_L g985 ( 
.A1(n_933),
.A2(n_808),
.B(n_794),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_888),
.B(n_762),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_818),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_812),
.A2(n_803),
.B(n_792),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_823),
.A2(n_804),
.B(n_803),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_835),
.B(n_668),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_834),
.B(n_830),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_896),
.Y(n_992)
);

OAI21xp33_ASAP7_75t_L g993 ( 
.A1(n_853),
.A2(n_708),
.B(n_706),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_891),
.A2(n_806),
.B(n_724),
.Y(n_994)
);

O2A1O1Ixp5_ASAP7_75t_L g995 ( 
.A1(n_877),
.A2(n_785),
.B(n_794),
.C(n_798),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_856),
.A2(n_807),
.B1(n_785),
.B2(n_798),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_830),
.B(n_654),
.Y(n_997)
);

NOR3xp33_ASAP7_75t_L g998 ( 
.A(n_819),
.B(n_761),
.C(n_753),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_891),
.A2(n_841),
.B(n_840),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_826),
.Y(n_1000)
);

INVx3_ASAP7_75t_SL g1001 ( 
.A(n_915),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_810),
.A2(n_960),
.B(n_877),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_820),
.B(n_762),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_829),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_912),
.B(n_773),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_872),
.B(n_778),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_850),
.B(n_662),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_841),
.A2(n_754),
.B(n_752),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_950),
.A2(n_730),
.B(n_671),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_848),
.A2(n_800),
.B(n_799),
.C(n_789),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_831),
.B(n_773),
.Y(n_1011)
);

AO21x1_ASAP7_75t_L g1012 ( 
.A1(n_823),
.A2(n_767),
.B(n_757),
.Y(n_1012)
);

O2A1O1Ixp5_ASAP7_75t_L g1013 ( 
.A1(n_880),
.A2(n_901),
.B(n_842),
.C(n_903),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_895),
.A2(n_923),
.B(n_921),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_861),
.B(n_664),
.Y(n_1015)
);

AO21x1_ASAP7_75t_L g1016 ( 
.A1(n_842),
.A2(n_771),
.B(n_768),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_884),
.B(n_671),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_879),
.A2(n_783),
.B1(n_730),
.B2(n_736),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_846),
.A2(n_764),
.B1(n_749),
.B2(n_736),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_895),
.A2(n_749),
.B(n_736),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_846),
.A2(n_764),
.B1(n_749),
.B2(n_727),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_900),
.A2(n_764),
.B1(n_710),
.B2(n_727),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_L g1023 ( 
.A(n_867),
.B(n_779),
.C(n_759),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_840),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_L g1025 ( 
.A(n_890),
.B(n_766),
.C(n_759),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_889),
.B(n_709),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_921),
.A2(n_710),
.B(n_709),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_926),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_813),
.B(n_751),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_923),
.A2(n_769),
.B(n_751),
.Y(n_1030)
);

BUFx4f_ASAP7_75t_L g1031 ( 
.A(n_926),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_854),
.B(n_664),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_826),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_862),
.A2(n_678),
.B(n_682),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_925),
.B(n_755),
.Y(n_1035)
);

CKINVDCx10_ASAP7_75t_R g1036 ( 
.A(n_967),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_816),
.B(n_857),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_826),
.B(n_678),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_824),
.B(n_807),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_906),
.A2(n_755),
.B(n_715),
.C(n_693),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_910),
.A2(n_755),
.B(n_715),
.C(n_693),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_902),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_863),
.B(n_783),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_894),
.A2(n_807),
.B1(n_755),
.B2(n_693),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_927),
.B(n_807),
.Y(n_1045)
);

AO21x1_ASAP7_75t_L g1046 ( 
.A1(n_941),
.A2(n_596),
.B(n_569),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_SL g1047 ( 
.A(n_836),
.B(n_807),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_897),
.A2(n_371),
.B(n_369),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_821),
.B(n_693),
.Y(n_1049)
);

AOI21x1_ASAP7_75t_L g1050 ( 
.A1(n_905),
.A2(n_596),
.B(n_569),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_860),
.B(n_796),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_904),
.A2(n_796),
.B1(n_801),
.B2(n_790),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_969),
.A2(n_796),
.B(n_801),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_875),
.A2(n_801),
.B(n_790),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_952),
.A2(n_610),
.B(n_569),
.C(n_571),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_875),
.A2(n_790),
.B(n_610),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_908),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_864),
.A2(n_883),
.B(n_868),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_932),
.B(n_790),
.Y(n_1059)
);

OAI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_924),
.A2(n_341),
.B(n_262),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_886),
.A2(n_962),
.B(n_977),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_829),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_829),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_886),
.A2(n_602),
.B(n_596),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_849),
.A2(n_367),
.B1(n_267),
.B2(n_269),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_905),
.A2(n_610),
.B(n_602),
.Y(n_1066)
);

NAND2x1_ASAP7_75t_L g1067 ( 
.A(n_962),
.B(n_566),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_945),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_811),
.B(n_6),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_962),
.A2(n_592),
.B(n_571),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_935),
.B(n_259),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_954),
.B(n_955),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_956),
.B(n_274),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_864),
.A2(n_883),
.B(n_868),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_898),
.A2(n_922),
.B(n_918),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_898),
.A2(n_592),
.B(n_588),
.C(n_571),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_915),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_971),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_876),
.B(n_284),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_918),
.A2(n_592),
.B(n_588),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_922),
.A2(n_602),
.B(n_588),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_909),
.B(n_287),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_929),
.A2(n_377),
.B(n_290),
.Y(n_1083)
);

AO21x1_ASAP7_75t_L g1084 ( 
.A1(n_892),
.A2(n_266),
.B(n_337),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_937),
.B(n_292),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_896),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_911),
.B(n_307),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_929),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_934),
.A2(n_387),
.B(n_310),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_814),
.A2(n_383),
.B(n_315),
.C(n_428),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_944),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_952),
.A2(n_7),
.B(n_8),
.C(n_10),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_843),
.B(n_851),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_944),
.A2(n_394),
.B(n_323),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_947),
.A2(n_395),
.B(n_328),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_964),
.B(n_8),
.Y(n_1096)
);

AO21x1_ASAP7_75t_L g1097 ( 
.A1(n_892),
.A2(n_266),
.B(n_337),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_947),
.A2(n_401),
.B(n_330),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_825),
.B(n_11),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_843),
.B(n_329),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_809),
.A2(n_882),
.B(n_948),
.C(n_946),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_915),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_953),
.A2(n_402),
.B(n_331),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_827),
.B(n_881),
.Y(n_1104)
);

BUFx8_ASAP7_75t_SL g1105 ( 
.A(n_935),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_865),
.B(n_339),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_965),
.B(n_354),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_953),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_855),
.B(n_881),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_957),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_869),
.A2(n_407),
.B(n_400),
.C(n_417),
.Y(n_1111)
);

AOI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_839),
.A2(n_411),
.B(n_405),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_881),
.B(n_935),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_832),
.B(n_14),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_896),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_870),
.B(n_590),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_957),
.A2(n_566),
.B(n_584),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_855),
.B(n_18),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_966),
.A2(n_973),
.B(n_968),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_878),
.A2(n_566),
.B1(n_337),
.B2(n_590),
.Y(n_1120)
);

OA21x2_ASAP7_75t_L g1121 ( 
.A1(n_966),
.A2(n_590),
.B(n_584),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_968),
.A2(n_590),
.B(n_584),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_938),
.B(n_25),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_837),
.A2(n_590),
.B(n_28),
.C(n_29),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_870),
.B(n_590),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_973),
.A2(n_566),
.B(n_217),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_914),
.B(n_27),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_916),
.B(n_31),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_855),
.B(n_31),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_917),
.B(n_939),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_870),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_871),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_1132)
);

NAND2x1_ASAP7_75t_L g1133 ( 
.A(n_931),
.B(n_210),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_974),
.A2(n_207),
.B(n_200),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_855),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_878),
.A2(n_198),
.B(n_188),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_833),
.B(n_35),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_873),
.A2(n_37),
.B(n_41),
.C(n_43),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_940),
.B(n_942),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_845),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_870),
.B(n_41),
.Y(n_1141)
);

BUFx12f_ASAP7_75t_L g1142 ( 
.A(n_920),
.Y(n_1142)
);

NOR3xp33_ASAP7_75t_L g1143 ( 
.A(n_899),
.B(n_44),
.C(n_46),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_SL g1144 ( 
.A(n_915),
.B(n_44),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_943),
.B(n_47),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_874),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_833),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_930),
.B(n_48),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_847),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_893),
.A2(n_961),
.B(n_928),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_976),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_844),
.B(n_53),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_828),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_828),
.B(n_57),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_913),
.A2(n_100),
.B(n_171),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_858),
.B(n_58),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_828),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_984),
.A2(n_859),
.B(n_975),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1004),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_981),
.A2(n_975),
.B(n_961),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1013),
.A2(n_963),
.B(n_913),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1005),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1006),
.B(n_828),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1139),
.B(n_828),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1061),
.A2(n_959),
.B(n_928),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_989),
.A2(n_963),
.B(n_959),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_991),
.B(n_866),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1042),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1013),
.A2(n_978),
.B(n_970),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1096),
.A2(n_951),
.B(n_885),
.C(n_936),
.Y(n_1170)
);

AOI221xp5_ASAP7_75t_L g1171 ( 
.A1(n_991),
.A2(n_972),
.B1(n_949),
.B2(n_907),
.C(n_919),
.Y(n_1171)
);

OAI22x1_ASAP7_75t_L g1172 ( 
.A1(n_1129),
.A2(n_887),
.B1(n_828),
.B2(n_866),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1003),
.B(n_958),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1004),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1057),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_987),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1139),
.B(n_958),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_990),
.A2(n_103),
.B(n_168),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_982),
.A2(n_1072),
.B1(n_1099),
.B2(n_1096),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_995),
.A2(n_60),
.B(n_62),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1062),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1031),
.Y(n_1182)
);

AOI221x1_ASAP7_75t_L g1183 ( 
.A1(n_1069),
.A2(n_64),
.B1(n_67),
.B2(n_69),
.C(n_73),
.Y(n_1183)
);

AOI21xp33_ASAP7_75t_L g1184 ( 
.A1(n_1156),
.A2(n_1069),
.B(n_1099),
.Y(n_1184)
);

AO21x1_ASAP7_75t_L g1185 ( 
.A1(n_1126),
.A2(n_116),
.B(n_156),
.Y(n_1185)
);

INVxp67_ASAP7_75t_L g1186 ( 
.A(n_1011),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1072),
.B(n_64),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_980),
.A2(n_114),
.B(n_148),
.Y(n_1188)
);

AO21x1_ASAP7_75t_L g1189 ( 
.A1(n_1156),
.A2(n_175),
.B(n_141),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1076),
.A2(n_983),
.B(n_999),
.Y(n_1190)
);

AOI21xp33_ASAP7_75t_L g1191 ( 
.A1(n_985),
.A2(n_73),
.B(n_74),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1002),
.A2(n_138),
.B(n_132),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1068),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1104),
.B(n_74),
.Y(n_1194)
);

OA21x2_ASAP7_75t_L g1195 ( 
.A1(n_1012),
.A2(n_123),
.B(n_121),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1074),
.A2(n_84),
.B(n_79),
.Y(n_1196)
);

AOI211x1_ASAP7_75t_L g1197 ( 
.A1(n_1078),
.A2(n_75),
.B(n_79),
.C(n_80),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_994),
.A2(n_81),
.B(n_82),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_L g1199 ( 
.A1(n_1016),
.A2(n_83),
.B(n_84),
.C(n_1046),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1028),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1101),
.A2(n_998),
.B(n_995),
.C(n_997),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1009),
.A2(n_988),
.B(n_1014),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1088),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1091),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1075),
.A2(n_1119),
.B(n_1058),
.Y(n_1205)
);

AOI21x1_ASAP7_75t_SL g1206 ( 
.A1(n_1154),
.A2(n_1114),
.B(n_1128),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1008),
.A2(n_1034),
.B(n_1122),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_998),
.A2(n_997),
.B(n_1129),
.C(n_1118),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1104),
.A2(n_1010),
.B(n_1085),
.C(n_1023),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1020),
.A2(n_993),
.B(n_1027),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_1031),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1030),
.A2(n_1007),
.B(n_1056),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1150),
.A2(n_1081),
.B(n_1070),
.Y(n_1213)
);

AOI211x1_ASAP7_75t_L g1214 ( 
.A1(n_1131),
.A2(n_1148),
.B(n_1127),
.C(n_1123),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1045),
.A2(n_1157),
.B(n_1041),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1090),
.A2(n_1039),
.B(n_1055),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1064),
.A2(n_1117),
.B(n_1080),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1051),
.A2(n_1054),
.B(n_1019),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1067),
.A2(n_1059),
.B(n_1021),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1032),
.B(n_1107),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1024),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1153),
.A2(n_1145),
.B1(n_996),
.B2(n_1093),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1109),
.B(n_1000),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_996),
.A2(n_1018),
.B(n_1124),
.Y(n_1224)
);

AOI221xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1138),
.A2(n_1146),
.B1(n_1151),
.B2(n_1092),
.C(n_1132),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1130),
.B(n_1140),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_986),
.B(n_1113),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1037),
.A2(n_1136),
.B(n_1111),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1001),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1053),
.A2(n_1022),
.B(n_1029),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1077),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1029),
.A2(n_1082),
.B(n_1116),
.Y(n_1232)
);

NOR3xp33_ASAP7_75t_L g1233 ( 
.A(n_1143),
.B(n_1071),
.C(n_1113),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1108),
.B(n_1110),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1037),
.A2(n_1023),
.B(n_1094),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1121),
.A2(n_1134),
.B(n_1052),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1125),
.A2(n_1049),
.B(n_1017),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1033),
.B(n_1149),
.Y(n_1238)
);

OAI22x1_ASAP7_75t_L g1239 ( 
.A1(n_1025),
.A2(n_1135),
.B1(n_1137),
.B2(n_1079),
.Y(n_1239)
);

AOI222xp33_ASAP7_75t_L g1240 ( 
.A1(n_1142),
.A2(n_1144),
.B1(n_1036),
.B2(n_1135),
.C1(n_1152),
.C2(n_1106),
.Y(n_1240)
);

INVx8_ASAP7_75t_L g1241 ( 
.A(n_1105),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1017),
.A2(n_1073),
.B(n_1089),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1137),
.A2(n_1141),
.B1(n_1143),
.B2(n_1038),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1035),
.A2(n_1098),
.B(n_1026),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1149),
.B(n_1026),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1062),
.B(n_1063),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1084),
.A2(n_1097),
.A3(n_1040),
.B(n_1087),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1063),
.B(n_1086),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1015),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1043),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1121),
.A2(n_1133),
.B(n_1155),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1083),
.A2(n_1095),
.B(n_1103),
.Y(n_1252)
);

OAI22x1_ASAP7_75t_L g1253 ( 
.A1(n_1001),
.A2(n_1044),
.B1(n_1065),
.B2(n_1100),
.Y(n_1253)
);

OAI21xp33_ASAP7_75t_L g1254 ( 
.A1(n_1048),
.A2(n_1060),
.B(n_1047),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1115),
.B(n_979),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1120),
.A2(n_1043),
.B(n_992),
.Y(n_1256)
);

OR2x6_ASAP7_75t_L g1257 ( 
.A(n_1147),
.B(n_979),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1112),
.A2(n_979),
.B(n_992),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_979),
.A2(n_992),
.B(n_1147),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1013),
.A2(n_981),
.B(n_995),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_984),
.B(n_1006),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_984),
.B(n_1006),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1012),
.A2(n_1016),
.A3(n_1046),
.B(n_985),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1137),
.B(n_915),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1042),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1042),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1001),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1031),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_991),
.B(n_838),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1013),
.A2(n_981),
.B(n_995),
.Y(n_1270)
);

OA22x2_ASAP7_75t_L g1271 ( 
.A1(n_986),
.A2(n_698),
.B1(n_723),
.B2(n_831),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_989),
.A2(n_1066),
.B(n_1050),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_989),
.A2(n_1066),
.B(n_1050),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_989),
.A2(n_1066),
.B(n_1050),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_984),
.B(n_1006),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1012),
.A2(n_1016),
.B(n_1046),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_984),
.A2(n_981),
.B(n_1061),
.Y(n_1277)
);

OA22x2_ASAP7_75t_L g1278 ( 
.A1(n_986),
.A2(n_698),
.B1(n_723),
.B2(n_831),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_989),
.A2(n_1066),
.B(n_1050),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1077),
.B(n_1102),
.Y(n_1280)
);

NAND2x1_ASAP7_75t_L g1281 ( 
.A(n_1004),
.B(n_1062),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1003),
.B(n_443),
.Y(n_1282)
);

AOI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1050),
.A2(n_1066),
.B(n_1046),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_984),
.A2(n_981),
.B(n_1061),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_984),
.A2(n_981),
.B(n_1061),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1042),
.Y(n_1286)
);

OA22x2_ASAP7_75t_L g1287 ( 
.A1(n_986),
.A2(n_698),
.B1(n_723),
.B2(n_831),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_989),
.A2(n_1066),
.B(n_1050),
.Y(n_1288)
);

AOI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1050),
.A2(n_1066),
.B(n_1046),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1013),
.A2(n_981),
.B(n_995),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1147),
.B(n_861),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_1028),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1013),
.A2(n_981),
.B(n_995),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_984),
.A2(n_981),
.B(n_1061),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_984),
.A2(n_981),
.B(n_1061),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_984),
.B(n_1006),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1012),
.A2(n_1016),
.A3(n_1046),
.B(n_985),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_989),
.A2(n_1066),
.B(n_1050),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_991),
.B(n_838),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_991),
.B(n_838),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1001),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_984),
.B(n_1006),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1012),
.A2(n_1016),
.A3(n_1046),
.B(n_985),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_984),
.A2(n_981),
.B(n_1061),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_984),
.B(n_838),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_984),
.B(n_838),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1011),
.B(n_733),
.Y(n_1307)
);

NAND2x1_ASAP7_75t_L g1308 ( 
.A(n_1004),
.B(n_1062),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_989),
.A2(n_1066),
.B(n_1050),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1269),
.B(n_1299),
.Y(n_1310)
);

AOI21xp33_ASAP7_75t_L g1311 ( 
.A1(n_1184),
.A2(n_1179),
.B(n_1282),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1179),
.A2(n_1305),
.B1(n_1306),
.B2(n_1296),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1229),
.Y(n_1313)
);

NAND2xp33_ASAP7_75t_L g1314 ( 
.A(n_1261),
.B(n_1262),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1229),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1300),
.B(n_1261),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1257),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1221),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1262),
.B(n_1275),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1245),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1175),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1277),
.A2(n_1285),
.B(n_1284),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1271),
.A2(n_1287),
.B1(n_1278),
.B2(n_1187),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1203),
.Y(n_1324)
);

BUFx12f_ASAP7_75t_L g1325 ( 
.A(n_1200),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1257),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1264),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1294),
.A2(n_1304),
.B(n_1295),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1275),
.B(n_1296),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1184),
.A2(n_1208),
.B(n_1302),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1209),
.A2(n_1235),
.B(n_1201),
.C(n_1224),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1302),
.A2(n_1187),
.B1(n_1220),
.B2(n_1194),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1164),
.A2(n_1163),
.B(n_1222),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1193),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1264),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1307),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1257),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1227),
.B(n_1226),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1186),
.B(n_1162),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1265),
.Y(n_1340)
);

BUFx12f_ASAP7_75t_L g1341 ( 
.A(n_1229),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1271),
.B(n_1278),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1204),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1226),
.B(n_1223),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1266),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1267),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1238),
.B(n_1173),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1286),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1234),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1267),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1238),
.B(n_1171),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1267),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1234),
.Y(n_1353)
);

INVx3_ASAP7_75t_SL g1354 ( 
.A(n_1241),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1212),
.A2(n_1202),
.B(n_1228),
.Y(n_1355)
);

INVx3_ASAP7_75t_SL g1356 ( 
.A(n_1241),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1301),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1233),
.B(n_1245),
.Y(n_1358)
);

INVxp67_ASAP7_75t_SL g1359 ( 
.A(n_1260),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1249),
.B(n_1250),
.Y(n_1360)
);

O2A1O1Ixp5_ASAP7_75t_L g1361 ( 
.A1(n_1228),
.A2(n_1185),
.B(n_1180),
.C(n_1235),
.Y(n_1361)
);

INVx3_ASAP7_75t_SL g1362 ( 
.A(n_1241),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1287),
.A2(n_1222),
.B1(n_1224),
.B2(n_1243),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1301),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1240),
.B(n_1239),
.Y(n_1365)
);

NAND2xp33_ASAP7_75t_L g1366 ( 
.A(n_1180),
.B(n_1260),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1291),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1280),
.B(n_1182),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1164),
.B(n_1177),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1183),
.A2(n_1194),
.B1(n_1243),
.B2(n_1177),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1167),
.B(n_1211),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1301),
.B(n_1268),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1231),
.B(n_1259),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1210),
.A2(n_1230),
.B(n_1218),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1259),
.B(n_1159),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1291),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1170),
.A2(n_1214),
.B1(n_1163),
.B2(n_1246),
.Y(n_1377)
);

OAI21xp33_ASAP7_75t_L g1378 ( 
.A1(n_1191),
.A2(n_1198),
.B(n_1254),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1292),
.A2(n_1172),
.B1(n_1225),
.B2(n_1253),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1196),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1255),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1159),
.B(n_1181),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1215),
.B(n_1258),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1270),
.A2(n_1293),
.B(n_1290),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1174),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1174),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1181),
.B(n_1248),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1248),
.B(n_1246),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1258),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1256),
.B(n_1281),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1270),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1290),
.A2(n_1293),
.B(n_1158),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1191),
.B(n_1263),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1232),
.A2(n_1242),
.B1(n_1216),
.B2(n_1197),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1308),
.Y(n_1395)
);

CKINVDCx6p67_ASAP7_75t_R g1396 ( 
.A(n_1206),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1244),
.B(n_1237),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1189),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1216),
.B(n_1263),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1199),
.A2(n_1161),
.B(n_1169),
.C(n_1178),
.Y(n_1400)
);

O2A1O1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1161),
.A2(n_1169),
.B(n_1252),
.C(n_1219),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1297),
.B(n_1303),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1297),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1297),
.B(n_1303),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1207),
.B(n_1236),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1276),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1195),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1205),
.B(n_1251),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1192),
.Y(n_1409)
);

INVx3_ASAP7_75t_SL g1410 ( 
.A(n_1195),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1247),
.B(n_1190),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1166),
.Y(n_1412)
);

CKINVDCx11_ASAP7_75t_R g1413 ( 
.A(n_1188),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1272),
.A2(n_1273),
.B(n_1298),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1213),
.B(n_1217),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1247),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1309),
.Y(n_1417)
);

INVx5_ASAP7_75t_L g1418 ( 
.A(n_1160),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1165),
.B(n_1289),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1274),
.B(n_1279),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1288),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1305),
.B(n_1306),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1168),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1179),
.A2(n_1284),
.B(n_1277),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1264),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1305),
.B(n_1306),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1264),
.B(n_915),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1257),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1184),
.A2(n_1179),
.B(n_1208),
.C(n_1209),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1229),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1264),
.B(n_1000),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1307),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1269),
.B(n_1299),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1168),
.Y(n_1434)
);

INVx6_ASAP7_75t_SL g1435 ( 
.A(n_1264),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1264),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1162),
.B(n_1269),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1257),
.Y(n_1438)
);

NOR2xp67_ASAP7_75t_L g1439 ( 
.A(n_1211),
.B(n_926),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1179),
.A2(n_1306),
.B1(n_1305),
.B2(n_852),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1257),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1168),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1305),
.B(n_1306),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1168),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1282),
.A2(n_852),
.B1(n_819),
.B2(n_1003),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1168),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1176),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1264),
.B(n_1000),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1269),
.B(n_1299),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1179),
.A2(n_1284),
.B(n_1277),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1179),
.A2(n_1284),
.B(n_1277),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1229),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1179),
.A2(n_1306),
.B1(n_1305),
.B2(n_852),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1184),
.B(n_1179),
.Y(n_1454)
);

BUFx2_ASAP7_75t_SL g1455 ( 
.A(n_1292),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1282),
.A2(n_852),
.B1(n_819),
.B2(n_1003),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1179),
.A2(n_1284),
.B(n_1277),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1307),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1264),
.B(n_1000),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_1292),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1257),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1269),
.B(n_1299),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1176),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1264),
.B(n_915),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1264),
.Y(n_1465)
);

INVx5_ASAP7_75t_L g1466 ( 
.A(n_1257),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1168),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1345),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1383),
.B(n_1333),
.Y(n_1469)
);

BUFx8_ASAP7_75t_L g1470 ( 
.A(n_1325),
.Y(n_1470)
);

BUFx2_ASAP7_75t_R g1471 ( 
.A(n_1354),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1460),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1348),
.Y(n_1473)
);

CKINVDCx16_ASAP7_75t_R g1474 ( 
.A(n_1460),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1365),
.A2(n_1398),
.B1(n_1342),
.B2(n_1351),
.Y(n_1475)
);

BUFx2_ASAP7_75t_SL g1476 ( 
.A(n_1439),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1320),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1398),
.A2(n_1440),
.B1(n_1453),
.B2(n_1332),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1310),
.B(n_1433),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1321),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1334),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1340),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1363),
.A2(n_1323),
.B1(n_1311),
.B2(n_1454),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1317),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1423),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1363),
.A2(n_1323),
.B1(n_1454),
.B2(n_1445),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1312),
.A2(n_1330),
.B1(n_1358),
.B2(n_1416),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1434),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1442),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1456),
.A2(n_1314),
.B1(n_1370),
.B2(n_1426),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1314),
.A2(n_1370),
.B1(n_1443),
.B2(n_1422),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1381),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1444),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1422),
.A2(n_1426),
.B1(n_1443),
.B2(n_1379),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1354),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1331),
.A2(n_1429),
.B(n_1361),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1446),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1466),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1429),
.A2(n_1331),
.B1(n_1316),
.B2(n_1319),
.Y(n_1499)
);

NOR2x1_ASAP7_75t_R g1500 ( 
.A(n_1455),
.B(n_1341),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1467),
.Y(n_1501)
);

BUFx2_ASAP7_75t_R g1502 ( 
.A(n_1356),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1324),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1343),
.Y(n_1504)
);

CKINVDCx11_ASAP7_75t_R g1505 ( 
.A(n_1356),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1329),
.A2(n_1338),
.B1(n_1320),
.B2(n_1344),
.Y(n_1506)
);

AOI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1355),
.A2(n_1450),
.B(n_1457),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1360),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1435),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1449),
.B(n_1462),
.Y(n_1510)
);

AOI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1355),
.A2(n_1457),
.B(n_1424),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1368),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1402),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1424),
.A2(n_1450),
.B(n_1451),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1404),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1366),
.A2(n_1409),
.B1(n_1407),
.B2(n_1383),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1378),
.A2(n_1458),
.B1(n_1413),
.B2(n_1366),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_SL g1518 ( 
.A1(n_1383),
.A2(n_1403),
.B1(n_1377),
.B2(n_1432),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1315),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1322),
.A2(n_1328),
.B(n_1361),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1318),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1458),
.A2(n_1413),
.B1(n_1393),
.B2(n_1353),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1392),
.A2(n_1384),
.B(n_1397),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1380),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_1362),
.Y(n_1525)
);

OR2x6_ASAP7_75t_L g1526 ( 
.A(n_1427),
.B(n_1464),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1391),
.A2(n_1339),
.B1(n_1359),
.B2(n_1396),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1384),
.A2(n_1400),
.B(n_1394),
.Y(n_1528)
);

CKINVDCx11_ASAP7_75t_R g1529 ( 
.A(n_1362),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1375),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1359),
.B(n_1349),
.Y(n_1531)
);

BUFx2_ASAP7_75t_R g1532 ( 
.A(n_1372),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1339),
.A2(n_1399),
.B1(n_1369),
.B2(n_1347),
.Y(n_1533)
);

CKINVDCx11_ASAP7_75t_R g1534 ( 
.A(n_1368),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1315),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1447),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1387),
.A2(n_1385),
.B1(n_1388),
.B2(n_1386),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1352),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1352),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1463),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1346),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1375),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1373),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1369),
.A2(n_1410),
.B1(n_1459),
.B2(n_1448),
.Y(n_1544)
);

BUFx6f_ASAP7_75t_L g1545 ( 
.A(n_1317),
.Y(n_1545)
);

AOI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1421),
.A2(n_1419),
.B(n_1412),
.Y(n_1546)
);

AO21x1_ASAP7_75t_SL g1547 ( 
.A1(n_1411),
.A2(n_1382),
.B(n_1371),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1406),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1373),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1414),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1417),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1327),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1335),
.B(n_1465),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1425),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1436),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1410),
.A2(n_1431),
.B1(n_1448),
.B2(n_1459),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1386),
.A2(n_1400),
.B1(n_1313),
.B2(n_1350),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1326),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1326),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1420),
.A2(n_1389),
.B(n_1390),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1431),
.B(n_1313),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1337),
.Y(n_1562)
);

AO21x1_ASAP7_75t_L g1563 ( 
.A1(n_1401),
.A2(n_1420),
.B(n_1405),
.Y(n_1563)
);

OR2x6_ASAP7_75t_L g1564 ( 
.A(n_1427),
.B(n_1464),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1427),
.A2(n_1464),
.B1(n_1430),
.B2(n_1452),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1430),
.A2(n_1452),
.B1(n_1461),
.B2(n_1441),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1337),
.A2(n_1461),
.B1(n_1441),
.B2(n_1438),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1428),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1428),
.A2(n_1438),
.B1(n_1346),
.B2(n_1357),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1367),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1346),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1346),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1367),
.B(n_1376),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1357),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1408),
.Y(n_1575)
);

CKINVDCx16_ASAP7_75t_R g1576 ( 
.A(n_1350),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1357),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1364),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1364),
.A2(n_1395),
.B1(n_1418),
.B2(n_1415),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1415),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1418),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1405),
.Y(n_1582)
);

INVx8_ASAP7_75t_L g1583 ( 
.A(n_1418),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1363),
.B(n_1320),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1345),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1345),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1355),
.A2(n_1450),
.B(n_1424),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1460),
.Y(n_1588)
);

AO21x1_ASAP7_75t_L g1589 ( 
.A1(n_1311),
.A2(n_1184),
.B(n_1179),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1310),
.B(n_1433),
.Y(n_1590)
);

OA21x2_ASAP7_75t_L g1591 ( 
.A1(n_1322),
.A2(n_1328),
.B(n_1374),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1445),
.A2(n_1456),
.B1(n_1003),
.B2(n_1282),
.Y(n_1592)
);

OA21x2_ASAP7_75t_L g1593 ( 
.A1(n_1322),
.A2(n_1328),
.B(n_1374),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1345),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1363),
.A2(n_1184),
.B1(n_1323),
.B2(n_1278),
.Y(n_1595)
);

BUFx2_ASAP7_75t_R g1596 ( 
.A(n_1354),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1320),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1432),
.Y(n_1598)
);

CKINVDCx11_ASAP7_75t_R g1599 ( 
.A(n_1460),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1345),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1317),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1310),
.B(n_1433),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1437),
.B(n_1336),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1445),
.A2(n_1456),
.B1(n_1429),
.B2(n_1453),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1460),
.Y(n_1605)
);

AOI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1454),
.A2(n_1289),
.B(n_1283),
.Y(n_1606)
);

OA21x2_ASAP7_75t_L g1607 ( 
.A1(n_1322),
.A2(n_1328),
.B(n_1374),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1355),
.A2(n_1450),
.B(n_1424),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1531),
.B(n_1530),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1604),
.A2(n_1584),
.B1(n_1496),
.B2(n_1499),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1477),
.B(n_1597),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1541),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1531),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1583),
.Y(n_1614)
);

AOI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1507),
.A2(n_1511),
.B(n_1514),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1506),
.B(n_1494),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1583),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1552),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1530),
.B(n_1542),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1541),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1479),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1534),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1506),
.B(n_1491),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1592),
.A2(n_1478),
.B(n_1490),
.Y(n_1624)
);

OR2x6_ASAP7_75t_L g1625 ( 
.A(n_1469),
.B(n_1583),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1587),
.A2(n_1608),
.B(n_1528),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1530),
.B(n_1542),
.Y(n_1627)
);

OR2x6_ASAP7_75t_L g1628 ( 
.A(n_1469),
.B(n_1583),
.Y(n_1628)
);

OR2x6_ASAP7_75t_L g1629 ( 
.A(n_1469),
.B(n_1526),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1551),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1606),
.A2(n_1546),
.B(n_1591),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1554),
.Y(n_1632)
);

AO21x2_ASAP7_75t_L g1633 ( 
.A1(n_1524),
.A2(n_1589),
.B(n_1550),
.Y(n_1633)
);

NAND2x1p5_ASAP7_75t_L g1634 ( 
.A(n_1498),
.B(n_1581),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1469),
.B(n_1526),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1513),
.B(n_1515),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1534),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1533),
.B(n_1508),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1492),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1555),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1480),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1590),
.Y(n_1642)
);

OA21x2_ASAP7_75t_L g1643 ( 
.A1(n_1563),
.A2(n_1548),
.B(n_1483),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1533),
.B(n_1602),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1599),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1591),
.A2(n_1593),
.B(n_1607),
.Y(n_1646)
);

BUFx12f_ASAP7_75t_L g1647 ( 
.A(n_1599),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1481),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1482),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1485),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1605),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1488),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1489),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1493),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1497),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1501),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1523),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1560),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1603),
.B(n_1510),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1523),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1505),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1568),
.Y(n_1662)
);

OA21x2_ASAP7_75t_L g1663 ( 
.A1(n_1575),
.A2(n_1517),
.B(n_1486),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1582),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1580),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1575),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1581),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1549),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1468),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1526),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1584),
.B(n_1547),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1543),
.B(n_1522),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1473),
.Y(n_1673)
);

AO21x1_ASAP7_75t_L g1674 ( 
.A1(n_1527),
.A2(n_1537),
.B(n_1557),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1503),
.Y(n_1675)
);

OA21x2_ASAP7_75t_L g1676 ( 
.A1(n_1517),
.A2(n_1544),
.B(n_1579),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1504),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1585),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1586),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1564),
.B(n_1556),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1520),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1564),
.B(n_1556),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1594),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1538),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1520),
.B(n_1544),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1487),
.B(n_1519),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1600),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1520),
.Y(n_1688)
);

NOR3xp33_ASAP7_75t_L g1689 ( 
.A(n_1576),
.B(n_1474),
.C(n_1571),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1564),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1598),
.B(n_1535),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1484),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1591),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1593),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1539),
.B(n_1538),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1593),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1607),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1607),
.B(n_1595),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1572),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1521),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1574),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1553),
.B(n_1595),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1516),
.B(n_1578),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_SL g1704 ( 
.A(n_1577),
.B(n_1498),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1536),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1540),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1570),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1570),
.Y(n_1708)
);

CKINVDCx6p67_ASAP7_75t_R g1709 ( 
.A(n_1605),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1570),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1484),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1566),
.A2(n_1565),
.B(n_1518),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1484),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1512),
.Y(n_1714)
);

NAND2x1_ASAP7_75t_L g1715 ( 
.A(n_1569),
.B(n_1567),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1545),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1545),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1545),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1609),
.B(n_1475),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1709),
.B(n_1472),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1609),
.B(n_1561),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1613),
.B(n_1561),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1611),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1619),
.B(n_1512),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1619),
.B(n_1601),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1638),
.B(n_1601),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1611),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1627),
.B(n_1601),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1627),
.B(n_1545),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1641),
.B(n_1649),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1644),
.B(n_1588),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1685),
.B(n_1562),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1618),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1699),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1632),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1656),
.B(n_1588),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1681),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1701),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1685),
.B(n_1562),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1671),
.B(n_1559),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1648),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1648),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1633),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1657),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1656),
.B(n_1472),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1617),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1650),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1667),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1610),
.B(n_1562),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1650),
.B(n_1558),
.Y(n_1750)
);

NAND2x1p5_ASAP7_75t_L g1751 ( 
.A(n_1670),
.B(n_1715),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1652),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1667),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1652),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1629),
.B(n_1509),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1671),
.B(n_1573),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1634),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1653),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_R g1759 ( 
.A(n_1645),
.B(n_1525),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1698),
.B(n_1505),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1653),
.B(n_1529),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1633),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1654),
.B(n_1476),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1657),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1634),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1654),
.B(n_1529),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1681),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1640),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1684),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1655),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1614),
.B(n_1525),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1707),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1624),
.A2(n_1623),
.B1(n_1616),
.B2(n_1702),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1664),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1664),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1643),
.B(n_1500),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1633),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1709),
.B(n_1495),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1643),
.B(n_1495),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1665),
.Y(n_1780)
);

INVx2_ASAP7_75t_R g1781 ( 
.A(n_1660),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1660),
.Y(n_1782)
);

OAI31xp33_ASAP7_75t_L g1783 ( 
.A1(n_1686),
.A2(n_1471),
.A3(n_1502),
.B(n_1596),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1665),
.B(n_1532),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1626),
.B(n_1470),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1626),
.B(n_1470),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1626),
.B(n_1710),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1636),
.B(n_1672),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1629),
.B(n_1635),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_L g1790 ( 
.A(n_1617),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1708),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1626),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1741),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1779),
.B(n_1643),
.C(n_1689),
.Y(n_1794)
);

OAI21xp33_ASAP7_75t_SL g1795 ( 
.A1(n_1760),
.A2(n_1695),
.B(n_1621),
.Y(n_1795)
);

OAI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1773),
.A2(n_1703),
.B1(n_1643),
.B2(n_1691),
.C(n_1672),
.Y(n_1796)
);

NAND3xp33_ASAP7_75t_SL g1797 ( 
.A(n_1783),
.B(n_1674),
.C(n_1651),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1779),
.A2(n_1663),
.B1(n_1676),
.B2(n_1712),
.Y(n_1798)
);

OAI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1783),
.A2(n_1703),
.B1(n_1663),
.B2(n_1715),
.C(n_1668),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1760),
.B(n_1658),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1723),
.B(n_1659),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1719),
.A2(n_1663),
.B1(n_1674),
.B2(n_1676),
.Y(n_1802)
);

AOI221x1_ASAP7_75t_SL g1803 ( 
.A1(n_1730),
.A2(n_1688),
.B1(n_1696),
.B2(n_1694),
.C(n_1693),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1727),
.B(n_1642),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1741),
.Y(n_1805)
);

OAI21xp33_ASAP7_75t_L g1806 ( 
.A1(n_1787),
.A2(n_1662),
.B(n_1688),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1733),
.B(n_1662),
.Y(n_1807)
);

OAI21xp33_ASAP7_75t_L g1808 ( 
.A1(n_1787),
.A2(n_1710),
.B(n_1693),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1735),
.B(n_1711),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1721),
.B(n_1658),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1721),
.B(n_1622),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1740),
.B(n_1622),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1731),
.A2(n_1637),
.B1(n_1645),
.B2(n_1684),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1768),
.B(n_1711),
.Y(n_1814)
);

NAND3xp33_ASAP7_75t_L g1815 ( 
.A(n_1776),
.B(n_1718),
.C(n_1713),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1776),
.A2(n_1713),
.B(n_1716),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1732),
.B(n_1680),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1730),
.B(n_1668),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1731),
.A2(n_1637),
.B1(n_1661),
.B2(n_1647),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1740),
.B(n_1661),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1738),
.B(n_1718),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_L g1822 ( 
.A(n_1738),
.B(n_1716),
.C(n_1697),
.Y(n_1822)
);

NAND4xp25_ASAP7_75t_L g1823 ( 
.A(n_1761),
.B(n_1766),
.C(n_1745),
.D(n_1736),
.Y(n_1823)
);

NAND3xp33_ASAP7_75t_L g1824 ( 
.A(n_1774),
.B(n_1697),
.C(n_1696),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1732),
.B(n_1680),
.Y(n_1825)
);

NAND3xp33_ASAP7_75t_L g1826 ( 
.A(n_1775),
.B(n_1694),
.C(n_1663),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1734),
.B(n_1704),
.Y(n_1827)
);

NAND3xp33_ASAP7_75t_L g1828 ( 
.A(n_1780),
.B(n_1679),
.C(n_1683),
.Y(n_1828)
);

OAI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1785),
.A2(n_1634),
.B(n_1676),
.Y(n_1829)
);

OAI221xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1749),
.A2(n_1629),
.B1(n_1635),
.B2(n_1628),
.C(n_1625),
.Y(n_1830)
);

OA21x2_ASAP7_75t_L g1831 ( 
.A1(n_1743),
.A2(n_1646),
.B(n_1631),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1719),
.A2(n_1675),
.B1(n_1687),
.B2(n_1683),
.C(n_1679),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1739),
.B(n_1682),
.Y(n_1833)
);

NAND3xp33_ASAP7_75t_L g1834 ( 
.A(n_1763),
.B(n_1726),
.C(n_1791),
.Y(n_1834)
);

NAND3xp33_ASAP7_75t_L g1835 ( 
.A(n_1763),
.B(n_1726),
.C(n_1785),
.Y(n_1835)
);

OAI21xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1786),
.A2(n_1771),
.B(n_1766),
.Y(n_1836)
);

NAND4xp25_ASAP7_75t_L g1837 ( 
.A(n_1761),
.B(n_1620),
.C(n_1612),
.D(n_1687),
.Y(n_1837)
);

NAND2xp33_ASAP7_75t_SL g1838 ( 
.A(n_1759),
.B(n_1617),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1734),
.B(n_1704),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1722),
.B(n_1675),
.Y(n_1840)
);

NAND3xp33_ASAP7_75t_L g1841 ( 
.A(n_1786),
.B(n_1717),
.C(n_1666),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1722),
.B(n_1714),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1757),
.B(n_1692),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1742),
.B(n_1747),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1742),
.B(n_1714),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1769),
.B(n_1647),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1757),
.B(n_1692),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1739),
.B(n_1682),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1747),
.B(n_1669),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1725),
.B(n_1682),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1752),
.B(n_1639),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1752),
.B(n_1673),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1749),
.A2(n_1676),
.B1(n_1712),
.B2(n_1635),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1754),
.B(n_1673),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1748),
.B(n_1789),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1754),
.B(n_1677),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1758),
.B(n_1677),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1725),
.B(n_1630),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1788),
.B(n_1636),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1765),
.B(n_1692),
.Y(n_1860)
);

NOR3xp33_ASAP7_75t_L g1861 ( 
.A(n_1737),
.B(n_1615),
.C(n_1717),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1758),
.B(n_1678),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1728),
.B(n_1690),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1770),
.B(n_1678),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1728),
.B(n_1630),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1743),
.A2(n_1700),
.B1(n_1705),
.B2(n_1706),
.C(n_1666),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_L g1867 ( 
.A(n_1750),
.B(n_1700),
.C(n_1706),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1770),
.Y(n_1868)
);

NAND4xp25_ASAP7_75t_L g1869 ( 
.A(n_1736),
.B(n_1612),
.C(n_1620),
.D(n_1705),
.Y(n_1869)
);

OAI221xp5_ASAP7_75t_SL g1870 ( 
.A1(n_1745),
.A2(n_1635),
.B1(n_1625),
.B2(n_1628),
.C(n_1690),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1831),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1801),
.B(n_1840),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1855),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1818),
.B(n_1788),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1855),
.Y(n_1875)
);

BUFx2_ASAP7_75t_L g1876 ( 
.A(n_1855),
.Y(n_1876)
);

BUFx3_ASAP7_75t_L g1877 ( 
.A(n_1831),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1793),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1803),
.B(n_1808),
.Y(n_1879)
);

INVxp67_ASAP7_75t_SL g1880 ( 
.A(n_1824),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1805),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1868),
.B(n_1744),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1831),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1844),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1810),
.B(n_1767),
.Y(n_1885)
);

AND2x2_ASAP7_75t_SL g1886 ( 
.A(n_1802),
.B(n_1789),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1810),
.B(n_1767),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1800),
.B(n_1767),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1851),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1834),
.B(n_1782),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1807),
.B(n_1809),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1850),
.B(n_1792),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1822),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1800),
.B(n_1781),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1826),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1858),
.B(n_1781),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1858),
.B(n_1781),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1814),
.B(n_1772),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1865),
.B(n_1744),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1794),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1852),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1817),
.B(n_1792),
.Y(n_1902)
);

OAI21xp5_ASAP7_75t_SL g1903 ( 
.A1(n_1797),
.A2(n_1778),
.B(n_1771),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1865),
.B(n_1792),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1863),
.B(n_1792),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1854),
.Y(n_1906)
);

INVx1_ASAP7_75t_SL g1907 ( 
.A(n_1827),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1804),
.B(n_1772),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1821),
.B(n_1835),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1806),
.B(n_1748),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1829),
.B(n_1729),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1795),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1856),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1857),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1862),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1867),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1864),
.B(n_1764),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_1838),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1842),
.B(n_1753),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1825),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1833),
.B(n_1753),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1833),
.B(n_1724),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1848),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1849),
.Y(n_1924)
);

NAND2x1_ASAP7_75t_SL g1925 ( 
.A(n_1846),
.B(n_1755),
.Y(n_1925)
);

INVx2_ASAP7_75t_SL g1926 ( 
.A(n_1843),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1859),
.B(n_1750),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1848),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1878),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1871),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1912),
.B(n_1873),
.Y(n_1931)
);

NOR3xp33_ASAP7_75t_L g1932 ( 
.A(n_1900),
.B(n_1903),
.C(n_1895),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1878),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1878),
.Y(n_1934)
);

NAND2x1_ASAP7_75t_L g1935 ( 
.A(n_1918),
.B(n_1811),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1912),
.B(n_1812),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1916),
.Y(n_1937)
);

NOR5xp2_ASAP7_75t_L g1938 ( 
.A(n_1900),
.B(n_1836),
.C(n_1799),
.D(n_1796),
.E(n_1815),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1871),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1916),
.B(n_1828),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1912),
.B(n_1820),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1881),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1881),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1872),
.B(n_1802),
.Y(n_1944)
);

NAND2x1p5_ASAP7_75t_L g1945 ( 
.A(n_1918),
.B(n_1769),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1881),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1908),
.Y(n_1947)
);

INVxp67_ASAP7_75t_SL g1948 ( 
.A(n_1893),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1882),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1909),
.B(n_1845),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1882),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1876),
.B(n_1769),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1924),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1872),
.B(n_1832),
.Y(n_1954)
);

INVx2_ASAP7_75t_SL g1955 ( 
.A(n_1925),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1876),
.B(n_1923),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1924),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1872),
.B(n_1839),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1895),
.B(n_1924),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1871),
.Y(n_1960)
);

INVx1_ASAP7_75t_SL g1961 ( 
.A(n_1908),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1913),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1876),
.B(n_1846),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1923),
.B(n_1861),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1909),
.B(n_1823),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1895),
.B(n_1816),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1884),
.Y(n_1967)
);

INVxp67_ASAP7_75t_SL g1968 ( 
.A(n_1893),
.Y(n_1968)
);

OAI33xp33_ASAP7_75t_L g1969 ( 
.A1(n_1879),
.A2(n_1895),
.A3(n_1909),
.B1(n_1890),
.B2(n_1884),
.B3(n_1913),
.Y(n_1969)
);

NAND4xp75_ASAP7_75t_L g1970 ( 
.A(n_1886),
.B(n_1784),
.C(n_1720),
.D(n_1866),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1884),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1923),
.B(n_1813),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1879),
.B(n_1819),
.Y(n_1973)
);

O2A1O1Ixp5_ASAP7_75t_L g1974 ( 
.A1(n_1880),
.A2(n_1843),
.B(n_1847),
.C(n_1860),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1927),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1913),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1917),
.Y(n_1977)
);

INVx2_ASAP7_75t_SL g1978 ( 
.A(n_1925),
.Y(n_1978)
);

NOR3xp33_ASAP7_75t_SL g1979 ( 
.A(n_1903),
.B(n_1838),
.C(n_1837),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1880),
.B(n_1869),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1923),
.B(n_1756),
.Y(n_1981)
);

AOI21x1_ASAP7_75t_L g1982 ( 
.A1(n_1918),
.A2(n_1615),
.B(n_1860),
.Y(n_1982)
);

NAND2xp33_ASAP7_75t_SL g1983 ( 
.A(n_1979),
.B(n_1925),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1948),
.B(n_1907),
.Y(n_1984)
);

INVxp67_ASAP7_75t_SL g1985 ( 
.A(n_1968),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1942),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1942),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1946),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1946),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1932),
.B(n_1907),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1941),
.B(n_1923),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1969),
.B(n_1891),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1941),
.B(n_1923),
.Y(n_1993)
);

INVxp67_ASAP7_75t_SL g1994 ( 
.A(n_1937),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1929),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1950),
.B(n_1908),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_L g1997 ( 
.A(n_1973),
.B(n_1891),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1950),
.B(n_1927),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1931),
.Y(n_1999)
);

INVxp67_ASAP7_75t_L g2000 ( 
.A(n_1940),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1947),
.B(n_1890),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1933),
.Y(n_2002)
);

INVx2_ASAP7_75t_SL g2003 ( 
.A(n_1963),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1966),
.A2(n_1886),
.B(n_1890),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1961),
.B(n_1891),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1934),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1936),
.B(n_1926),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1954),
.B(n_1889),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1975),
.B(n_1965),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1958),
.B(n_1889),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1965),
.B(n_1927),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1943),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1936),
.B(n_1931),
.Y(n_2013)
);

NAND2x1_ASAP7_75t_L g2014 ( 
.A(n_1931),
.B(n_1875),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1977),
.B(n_1874),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1981),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1977),
.B(n_1874),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1963),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_1935),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1959),
.B(n_1949),
.Y(n_2020)
);

INVxp67_ASAP7_75t_SL g2021 ( 
.A(n_1938),
.Y(n_2021)
);

A2O1A1Ixp33_ASAP7_75t_L g2022 ( 
.A1(n_1980),
.A2(n_1886),
.B(n_1853),
.C(n_1798),
.Y(n_2022)
);

INVx2_ASAP7_75t_SL g2023 ( 
.A(n_1935),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1972),
.B(n_1873),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1953),
.Y(n_2025)
);

NAND2x1p5_ASAP7_75t_L g2026 ( 
.A(n_1955),
.B(n_1873),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1945),
.B(n_1926),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1944),
.B(n_1874),
.Y(n_2028)
);

NOR2x1_ASAP7_75t_L g2029 ( 
.A(n_1970),
.B(n_1873),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1957),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1949),
.B(n_1898),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1951),
.B(n_1889),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1951),
.B(n_1898),
.Y(n_2033)
);

HB1xp67_ASAP7_75t_L g2034 ( 
.A(n_1962),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1945),
.B(n_1926),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1967),
.Y(n_2036)
);

CKINVDCx16_ASAP7_75t_R g2037 ( 
.A(n_1983),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2034),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2034),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1986),
.Y(n_2040)
);

INVx4_ASAP7_75t_L g2041 ( 
.A(n_2013),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1987),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1988),
.Y(n_2043)
);

NOR2x1_ASAP7_75t_L g2044 ( 
.A(n_2029),
.B(n_1997),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_2011),
.B(n_1971),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1997),
.B(n_1962),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_2021),
.A2(n_1992),
.B1(n_2004),
.B2(n_2000),
.Y(n_2047)
);

BUFx2_ASAP7_75t_L g2048 ( 
.A(n_2003),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_SL g2049 ( 
.A(n_2014),
.B(n_1956),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1989),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1995),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2002),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_2021),
.B(n_1945),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_2018),
.Y(n_2054)
);

CKINVDCx16_ASAP7_75t_R g2055 ( 
.A(n_1983),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2006),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_1998),
.B(n_1976),
.Y(n_2057)
);

CKINVDCx16_ASAP7_75t_R g2058 ( 
.A(n_2024),
.Y(n_2058)
);

OAI221xp5_ASAP7_75t_L g2059 ( 
.A1(n_2022),
.A2(n_1978),
.B1(n_1955),
.B2(n_1877),
.C(n_1974),
.Y(n_2059)
);

INVx1_ASAP7_75t_SL g2060 ( 
.A(n_1990),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1992),
.A2(n_1978),
.B(n_1886),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2012),
.Y(n_2062)
);

NOR2x1_ASAP7_75t_L g2063 ( 
.A(n_1984),
.B(n_1970),
.Y(n_2063)
);

BUFx3_ASAP7_75t_L g2064 ( 
.A(n_1999),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_1985),
.B(n_1972),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2016),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1991),
.B(n_1956),
.Y(n_2067)
);

NOR2x1_ASAP7_75t_L g2068 ( 
.A(n_2007),
.B(n_2009),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_2015),
.B(n_1976),
.Y(n_2069)
);

NOR2xp33_ASAP7_75t_L g2070 ( 
.A(n_1985),
.B(n_1952),
.Y(n_2070)
);

INVx1_ASAP7_75t_SL g2071 ( 
.A(n_2028),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2025),
.Y(n_2072)
);

OAI22x1_ASAP7_75t_L g2073 ( 
.A1(n_1994),
.A2(n_1964),
.B1(n_1982),
.B2(n_1960),
.Y(n_2073)
);

OAI21x1_ASAP7_75t_L g2074 ( 
.A1(n_2026),
.A2(n_1982),
.B(n_1939),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2030),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1993),
.B(n_1952),
.Y(n_2076)
);

OAI22xp33_ASAP7_75t_L g2077 ( 
.A1(n_2059),
.A2(n_2000),
.B1(n_2008),
.B2(n_2001),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2058),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2038),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2039),
.Y(n_2080)
);

NAND3xp33_ASAP7_75t_SL g2081 ( 
.A(n_2047),
.B(n_2022),
.C(n_2007),
.Y(n_2081)
);

OAI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_2061),
.A2(n_2063),
.B1(n_2044),
.B2(n_2060),
.Y(n_2082)
);

OAI21xp5_ASAP7_75t_SL g2083 ( 
.A1(n_2047),
.A2(n_2026),
.B(n_1994),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2071),
.B(n_2005),
.Y(n_2084)
);

NAND3xp33_ASAP7_75t_L g2085 ( 
.A(n_2053),
.B(n_2065),
.C(n_2070),
.Y(n_2085)
);

OAI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_2037),
.A2(n_2019),
.B1(n_2023),
.B2(n_1996),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2065),
.B(n_2020),
.Y(n_2087)
);

OAI211xp5_ASAP7_75t_SL g2088 ( 
.A1(n_2068),
.A2(n_2035),
.B(n_2027),
.C(n_2033),
.Y(n_2088)
);

AOI22xp33_ASAP7_75t_L g2089 ( 
.A1(n_2073),
.A2(n_1877),
.B1(n_1853),
.B2(n_1939),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2054),
.B(n_2017),
.Y(n_2090)
);

AOI221x1_ASAP7_75t_L g2091 ( 
.A1(n_2073),
.A2(n_2053),
.B1(n_2049),
.B2(n_2070),
.C(n_2041),
.Y(n_2091)
);

AOI222xp33_ASAP7_75t_L g2092 ( 
.A1(n_2046),
.A2(n_1877),
.B1(n_1930),
.B2(n_1960),
.C1(n_1871),
.C2(n_1883),
.Y(n_2092)
);

NAND4xp25_ASAP7_75t_L g2093 ( 
.A(n_2041),
.B(n_2027),
.C(n_2035),
.D(n_1964),
.Y(n_2093)
);

AOI211xp5_ASAP7_75t_L g2094 ( 
.A1(n_2074),
.A2(n_1877),
.B(n_1883),
.C(n_1930),
.Y(n_2094)
);

INVx2_ASAP7_75t_SL g2095 ( 
.A(n_2041),
.Y(n_2095)
);

INVxp67_ASAP7_75t_L g2096 ( 
.A(n_2064),
.Y(n_2096)
);

HB1xp67_ASAP7_75t_L g2097 ( 
.A(n_2064),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2055),
.A2(n_1784),
.B1(n_1911),
.B2(n_2010),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2040),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2048),
.B(n_2036),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2066),
.B(n_2031),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2066),
.A2(n_1911),
.B1(n_1883),
.B2(n_2032),
.Y(n_2102)
);

OAI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_2074),
.A2(n_1910),
.B(n_1926),
.Y(n_2103)
);

OAI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2045),
.A2(n_1883),
.B1(n_1875),
.B2(n_1751),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2076),
.Y(n_2105)
);

A2O1A1Ixp33_ASAP7_75t_L g2106 ( 
.A1(n_2049),
.A2(n_2069),
.B(n_2057),
.C(n_2072),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2097),
.B(n_2051),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2078),
.B(n_2076),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2090),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2096),
.B(n_2052),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_2105),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2096),
.B(n_2056),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2084),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2087),
.B(n_2062),
.Y(n_2114)
);

AOI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_2081),
.A2(n_2069),
.B1(n_2075),
.B2(n_2050),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2095),
.Y(n_2116)
);

NOR2x1_ASAP7_75t_R g2117 ( 
.A(n_2100),
.B(n_2067),
.Y(n_2117)
);

INVx1_ASAP7_75t_SL g2118 ( 
.A(n_2101),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2085),
.B(n_2042),
.Y(n_2119)
);

AOI22xp33_ASAP7_75t_L g2120 ( 
.A1(n_2081),
.A2(n_2043),
.B1(n_2067),
.B2(n_1712),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2079),
.B(n_1889),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2099),
.Y(n_2122)
);

INVx3_ASAP7_75t_L g2123 ( 
.A(n_2080),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2083),
.B(n_1910),
.Y(n_2124)
);

AOI22xp5_ASAP7_75t_L g2125 ( 
.A1(n_2082),
.A2(n_1911),
.B1(n_1894),
.B2(n_1910),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2089),
.B(n_1920),
.Y(n_2126)
);

NOR2x1_ASAP7_75t_L g2127 ( 
.A(n_2106),
.B(n_1981),
.Y(n_2127)
);

INVx1_ASAP7_75t_SL g2128 ( 
.A(n_2086),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2102),
.Y(n_2129)
);

AOI221xp5_ASAP7_75t_L g2130 ( 
.A1(n_2115),
.A2(n_2077),
.B1(n_2088),
.B2(n_2103),
.C(n_2094),
.Y(n_2130)
);

AOI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_2129),
.A2(n_2092),
.B1(n_2098),
.B2(n_2088),
.Y(n_2131)
);

AOI222xp33_ASAP7_75t_L g2132 ( 
.A1(n_2120),
.A2(n_2091),
.B1(n_2104),
.B2(n_1762),
.C1(n_1777),
.C2(n_2093),
.Y(n_2132)
);

NOR3xp33_ASAP7_75t_SL g2133 ( 
.A(n_2119),
.B(n_1870),
.C(n_1847),
.Y(n_2133)
);

AOI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_2124),
.A2(n_1875),
.B(n_1898),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2125),
.A2(n_1875),
.B1(n_1919),
.B2(n_1894),
.Y(n_2135)
);

O2A1O1Ixp33_ASAP7_75t_L g2136 ( 
.A1(n_2123),
.A2(n_1894),
.B(n_1917),
.C(n_1896),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2118),
.B(n_1920),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2108),
.B(n_2128),
.Y(n_2138)
);

AOI221x1_ASAP7_75t_SL g2139 ( 
.A1(n_2109),
.A2(n_1902),
.B1(n_1892),
.B2(n_1920),
.C(n_1928),
.Y(n_2139)
);

NAND3xp33_ASAP7_75t_SL g2140 ( 
.A(n_2113),
.B(n_1897),
.C(n_1896),
.Y(n_2140)
);

NAND4xp25_ASAP7_75t_L g2141 ( 
.A(n_2108),
.B(n_1919),
.C(n_1888),
.D(n_1899),
.Y(n_2141)
);

AOI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_2129),
.A2(n_1777),
.B1(n_1762),
.B2(n_1917),
.C(n_1915),
.Y(n_2142)
);

OAI211xp5_ASAP7_75t_SL g2143 ( 
.A1(n_2127),
.A2(n_1919),
.B(n_1928),
.C(n_1920),
.Y(n_2143)
);

OAI322xp33_ASAP7_75t_L g2144 ( 
.A1(n_2131),
.A2(n_2113),
.A3(n_2109),
.B1(n_2114),
.B2(n_2107),
.C1(n_2112),
.C2(n_2110),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2138),
.Y(n_2145)
);

AOI22x1_ASAP7_75t_SL g2146 ( 
.A1(n_2141),
.A2(n_2116),
.B1(n_2122),
.B2(n_2111),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2134),
.B(n_2111),
.Y(n_2147)
);

NAND4xp25_ASAP7_75t_L g2148 ( 
.A(n_2130),
.B(n_2111),
.C(n_2116),
.D(n_2123),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2137),
.Y(n_2149)
);

AOI211xp5_ASAP7_75t_L g2150 ( 
.A1(n_2143),
.A2(n_2140),
.B(n_2117),
.C(n_2135),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2139),
.B(n_2123),
.Y(n_2151)
);

NOR2x1_ASAP7_75t_L g2152 ( 
.A(n_2136),
.B(n_2122),
.Y(n_2152)
);

NAND3xp33_ASAP7_75t_SL g2153 ( 
.A(n_2132),
.B(n_2126),
.C(n_2121),
.Y(n_2153)
);

NAND4xp25_ASAP7_75t_L g2154 ( 
.A(n_2142),
.B(n_1888),
.C(n_1899),
.D(n_1897),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2145),
.Y(n_2155)
);

NAND3xp33_ASAP7_75t_L g2156 ( 
.A(n_2148),
.B(n_2133),
.C(n_1897),
.Y(n_2156)
);

INVx2_ASAP7_75t_SL g2157 ( 
.A(n_2147),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2152),
.Y(n_2158)
);

AND4x1_ASAP7_75t_L g2159 ( 
.A(n_2150),
.B(n_1896),
.C(n_1899),
.D(n_1888),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2149),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_2144),
.B(n_1901),
.Y(n_2161)
);

NAND4xp25_ASAP7_75t_L g2162 ( 
.A(n_2151),
.B(n_1746),
.C(n_1887),
.D(n_1885),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_2158),
.A2(n_2153),
.B1(n_2146),
.B2(n_2154),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2157),
.Y(n_2164)
);

OAI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_2156),
.A2(n_1892),
.B1(n_1902),
.B2(n_1928),
.Y(n_2165)
);

NOR2x1_ASAP7_75t_L g2166 ( 
.A(n_2155),
.B(n_1892),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2160),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2161),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2161),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2159),
.Y(n_2170)
);

NAND4xp75_ASAP7_75t_L g2171 ( 
.A(n_2164),
.B(n_2162),
.C(n_1905),
.D(n_1904),
.Y(n_2171)
);

NAND4xp25_ASAP7_75t_L g2172 ( 
.A(n_2163),
.B(n_1746),
.C(n_1887),
.D(n_1885),
.Y(n_2172)
);

NOR2x1_ASAP7_75t_L g2173 ( 
.A(n_2167),
.B(n_1921),
.Y(n_2173)
);

NOR3xp33_ASAP7_75t_L g2174 ( 
.A(n_2168),
.B(n_2169),
.C(n_2170),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2166),
.Y(n_2175)
);

NOR3xp33_ASAP7_75t_L g2176 ( 
.A(n_2165),
.B(n_1841),
.C(n_1830),
.Y(n_2176)
);

NOR2x1_ASAP7_75t_L g2177 ( 
.A(n_2175),
.B(n_1921),
.Y(n_2177)
);

AND3x2_ASAP7_75t_L g2178 ( 
.A(n_2174),
.B(n_1921),
.C(n_1922),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2173),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2171),
.Y(n_2180)
);

AOI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2179),
.A2(n_2172),
.B1(n_2176),
.B2(n_1892),
.Y(n_2181)
);

OAI22xp5_ASAP7_75t_L g2182 ( 
.A1(n_2177),
.A2(n_1892),
.B1(n_1902),
.B2(n_1906),
.Y(n_2182)
);

NOR3xp33_ASAP7_75t_L g2183 ( 
.A(n_2181),
.B(n_2180),
.C(n_2182),
.Y(n_2183)
);

AOI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_2183),
.A2(n_2178),
.B1(n_1892),
.B2(n_1902),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2183),
.A2(n_1902),
.B1(n_1905),
.B2(n_1901),
.Y(n_2185)
);

OA22x2_ASAP7_75t_L g2186 ( 
.A1(n_2184),
.A2(n_1902),
.B1(n_1904),
.B2(n_1905),
.Y(n_2186)
);

HB1xp67_ASAP7_75t_L g2187 ( 
.A(n_2185),
.Y(n_2187)
);

AOI21xp5_ASAP7_75t_SL g2188 ( 
.A1(n_2187),
.A2(n_1790),
.B(n_1746),
.Y(n_2188)
);

AOI222xp33_ASAP7_75t_SL g2189 ( 
.A1(n_2188),
.A2(n_2186),
.B1(n_1928),
.B2(n_1901),
.C1(n_1906),
.C2(n_1914),
.Y(n_2189)
);

OAI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_2189),
.A2(n_1906),
.B1(n_1915),
.B2(n_1914),
.Y(n_2190)
);

AOI221xp5_ASAP7_75t_L g2191 ( 
.A1(n_2190),
.A2(n_1915),
.B1(n_1906),
.B2(n_1914),
.C(n_1901),
.Y(n_2191)
);

AOI211xp5_ASAP7_75t_L g2192 ( 
.A1(n_2191),
.A2(n_1790),
.B(n_1692),
.C(n_1617),
.Y(n_2192)
);


endmodule