module real_aes_342_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g239 ( .A(n_0), .B(n_154), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_1), .B(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_2), .B(n_138), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_3), .B(n_156), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_4), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g145 ( .A(n_5), .Y(n_145) );
NAND2xp33_ASAP7_75t_SL g224 ( .A(n_6), .B(n_144), .Y(n_224) );
INVx1_ASAP7_75t_L g215 ( .A(n_7), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g756 ( .A(n_8), .Y(n_756) );
AND2x2_ASAP7_75t_L g132 ( .A(n_9), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g462 ( .A(n_10), .B(n_185), .Y(n_462) );
AND2x2_ASAP7_75t_L g470 ( .A(n_11), .B(n_221), .Y(n_470) );
INVx2_ASAP7_75t_L g134 ( .A(n_12), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_13), .B(n_156), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_14), .Y(n_111) );
AOI221x1_ASAP7_75t_L g218 ( .A1(n_15), .A2(n_147), .B1(n_219), .B2(n_221), .C(n_223), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_16), .B(n_138), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_17), .B(n_138), .Y(n_502) );
INVx1_ASAP7_75t_L g115 ( .A(n_18), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_19), .A2(n_90), .B1(n_138), .B2(n_189), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_20), .A2(n_72), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_20), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_21), .A2(n_147), .B(n_152), .Y(n_146) );
AOI221xp5_ASAP7_75t_SL g229 ( .A1(n_22), .A2(n_35), .B1(n_138), .B2(n_147), .C(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_23), .B(n_154), .Y(n_153) );
OR2x2_ASAP7_75t_L g135 ( .A(n_24), .B(n_89), .Y(n_135) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_24), .A2(n_89), .B(n_134), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_25), .B(n_156), .Y(n_209) );
INVxp67_ASAP7_75t_L g217 ( .A(n_26), .Y(n_217) );
AND2x2_ASAP7_75t_L g178 ( .A(n_27), .B(n_168), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_28), .A2(n_147), .B(n_238), .Y(n_237) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_29), .A2(n_221), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_30), .B(n_156), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_31), .A2(n_147), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_32), .B(n_156), .Y(n_486) );
AND2x2_ASAP7_75t_L g144 ( .A(n_33), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g148 ( .A(n_33), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g197 ( .A(n_33), .Y(n_197) );
OR2x6_ASAP7_75t_L g113 ( .A(n_34), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_36), .B(n_138), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_37), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_38), .A2(n_82), .B1(n_147), .B2(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_39), .B(n_156), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_40), .B(n_138), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_41), .B(n_154), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_42), .A2(n_147), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g242 ( .A(n_43), .B(n_168), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_44), .B(n_154), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_45), .B(n_168), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_46), .B(n_138), .Y(n_475) );
INVx1_ASAP7_75t_L g141 ( .A(n_47), .Y(n_141) );
INVx1_ASAP7_75t_L g151 ( .A(n_47), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_48), .B(n_156), .Y(n_468) );
AND2x2_ASAP7_75t_L g493 ( .A(n_49), .B(n_168), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_50), .B(n_138), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_51), .B(n_154), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_52), .B(n_154), .Y(n_485) );
AND2x2_ASAP7_75t_L g169 ( .A(n_53), .B(n_168), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_54), .B(n_138), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_55), .B(n_156), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_56), .B(n_138), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_57), .A2(n_147), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_58), .B(n_154), .Y(n_165) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_59), .B(n_133), .Y(n_210) );
AND2x2_ASAP7_75t_L g508 ( .A(n_60), .B(n_133), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_61), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_62), .A2(n_147), .B(n_174), .Y(n_173) );
AOI22xp33_ASAP7_75t_SL g101 ( .A1(n_63), .A2(n_102), .B1(n_750), .B2(n_757), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_64), .B(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_SL g200 ( .A(n_65), .B(n_185), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_66), .B(n_154), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_67), .B(n_154), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_68), .A2(n_93), .B1(n_147), .B2(n_195), .Y(n_532) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_69), .A2(n_78), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx14_ASAP7_75t_R g120 ( .A(n_69), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_70), .B(n_156), .Y(n_505) );
INVx1_ASAP7_75t_L g143 ( .A(n_71), .Y(n_143) );
INVx1_ASAP7_75t_L g149 ( .A(n_71), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_72), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_73), .B(n_154), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_74), .A2(n_147), .B(n_497), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_75), .A2(n_147), .B(n_449), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_76), .A2(n_147), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g488 ( .A(n_77), .B(n_133), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_78), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_79), .B(n_168), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_80), .B(n_138), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_81), .A2(n_84), .B1(n_138), .B2(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g116 ( .A(n_83), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_85), .B(n_154), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_86), .B(n_154), .Y(n_232) );
AND2x2_ASAP7_75t_L g452 ( .A(n_87), .B(n_185), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_88), .A2(n_147), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_91), .B(n_156), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_92), .A2(n_147), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_94), .B(n_156), .Y(n_450) );
INVxp67_ASAP7_75t_L g220 ( .A(n_95), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_96), .B(n_138), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_97), .B(n_156), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_98), .A2(n_147), .B(n_207), .Y(n_206) );
BUFx2_ASAP7_75t_L g507 ( .A(n_99), .Y(n_507) );
BUFx2_ASAP7_75t_L g105 ( .A(n_100), .Y(n_105) );
INVx1_ASAP7_75t_SL g739 ( .A(n_100), .Y(n_739) );
AO21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_106), .B(n_737), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_117), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_108), .A2(n_741), .B(n_746), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
BUFx3_ASAP7_75t_L g749 ( .A(n_110), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x6_ASAP7_75t_SL g122 ( .A(n_111), .B(n_113), .Y(n_122) );
OR2x6_ASAP7_75t_SL g437 ( .A(n_111), .B(n_112), .Y(n_437) );
OR2x2_ASAP7_75t_L g736 ( .A(n_111), .B(n_113), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AOI221x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_121), .B1(n_729), .B2(n_732), .C(n_733), .Y(n_117) );
INVxp67_ASAP7_75t_SL g732 ( .A(n_118), .Y(n_732) );
AO22x2_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_436), .B2(n_438), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_122), .B(n_124), .Y(n_731) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
XNOR2xp5_ASAP7_75t_L g742 ( .A(n_124), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_358), .Y(n_124) );
NOR3xp33_ASAP7_75t_SL g125 ( .A(n_126), .B(n_282), .C(n_332), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_262), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_201), .B(n_243), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_179), .Y(n_129) );
INVx1_ASAP7_75t_SL g368 ( .A(n_130), .Y(n_368) );
AOI32xp33_ASAP7_75t_L g399 ( .A1(n_130), .A2(n_381), .A3(n_400), .B1(n_401), .B2(n_402), .Y(n_399) );
AND2x2_ASAP7_75t_L g401 ( .A(n_130), .B(n_258), .Y(n_401) );
AND2x4_ASAP7_75t_SL g130 ( .A(n_131), .B(n_159), .Y(n_130) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
INVx5_ASAP7_75t_L g261 ( .A(n_131), .Y(n_261) );
OR2x2_ASAP7_75t_L g268 ( .A(n_131), .B(n_260), .Y(n_268) );
INVx2_ASAP7_75t_L g273 ( .A(n_131), .Y(n_273) );
AND2x2_ASAP7_75t_L g285 ( .A(n_131), .B(n_160), .Y(n_285) );
AND2x2_ASAP7_75t_L g290 ( .A(n_131), .B(n_170), .Y(n_290) );
OR2x2_ASAP7_75t_L g297 ( .A(n_131), .B(n_182), .Y(n_297) );
AND2x4_ASAP7_75t_L g306 ( .A(n_131), .B(n_171), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_SL g348 ( .A1(n_131), .A2(n_264), .B(n_299), .C(n_337), .Y(n_348) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x4_ASAP7_75t_L g158 ( .A(n_134), .B(n_135), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_146), .B(n_158), .Y(n_136) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
INVx1_ASAP7_75t_L g225 ( .A(n_139), .Y(n_225) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
AND2x6_ASAP7_75t_L g154 ( .A(n_140), .B(n_149), .Y(n_154) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g156 ( .A(n_142), .B(n_151), .Y(n_156) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx5_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
AND2x2_ASAP7_75t_L g150 ( .A(n_145), .B(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_145), .Y(n_192) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
BUFx3_ASAP7_75t_L g193 ( .A(n_148), .Y(n_193) );
INVx2_ASAP7_75t_L g199 ( .A(n_149), .Y(n_199) );
AND2x4_ASAP7_75t_L g195 ( .A(n_150), .B(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_155), .B(n_157), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_154), .B(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_157), .A2(n_164), .B(n_165), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_157), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_157), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_157), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_157), .A2(n_239), .B(n_240), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_157), .A2(n_450), .B(n_451), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_157), .A2(n_459), .B(n_460), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_157), .A2(n_467), .B(n_468), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_157), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_157), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_157), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_157), .A2(n_505), .B(n_506), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_158), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_158), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_158), .B(n_220), .Y(n_219) );
NOR3xp33_ASAP7_75t_L g223 ( .A(n_158), .B(n_224), .C(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_158), .A2(n_475), .B(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_158), .A2(n_495), .B(n_496), .Y(n_494) );
INVx3_ASAP7_75t_SL g298 ( .A(n_159), .Y(n_298) );
AND2x2_ASAP7_75t_L g344 ( .A(n_159), .B(n_261), .Y(n_344) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_170), .Y(n_159) );
AND2x2_ASAP7_75t_L g181 ( .A(n_160), .B(n_182), .Y(n_181) );
OR2x2_ASAP7_75t_L g275 ( .A(n_160), .B(n_171), .Y(n_275) );
AND2x2_ASAP7_75t_L g279 ( .A(n_160), .B(n_258), .Y(n_279) );
INVx1_ASAP7_75t_L g305 ( .A(n_160), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_160), .B(n_171), .Y(n_327) );
INVx2_ASAP7_75t_L g331 ( .A(n_160), .Y(n_331) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_160), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_160), .B(n_261), .Y(n_408) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_167), .B(n_169), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_166), .Y(n_161) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_167), .A2(n_172), .B(n_178), .Y(n_171) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_167), .A2(n_172), .B(n_178), .Y(n_260) );
AOI21x1_ASAP7_75t_L g455 ( .A1(n_167), .A2(n_456), .B(n_462), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_168), .A2(n_229), .B(n_233), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_168), .A2(n_447), .B(n_448), .Y(n_446) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_168), .A2(n_531), .B(n_532), .Y(n_530) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g342 ( .A(n_171), .B(n_182), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_177), .Y(n_172) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx1_ASAP7_75t_L g352 ( .A(n_180), .Y(n_352) );
NAND2xp33_ASAP7_75t_SL g377 ( .A(n_180), .B(n_269), .Y(n_377) );
AND2x2_ASAP7_75t_L g419 ( .A(n_181), .B(n_261), .Y(n_419) );
AND2x2_ASAP7_75t_L g330 ( .A(n_182), .B(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g393 ( .A(n_182), .Y(n_393) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
AOI21x1_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_187), .B(n_200), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_185), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_185), .A2(n_502), .B(n_503), .Y(n_501) );
BUFx4f_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx3_ASAP7_75t_L g222 ( .A(n_186), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_194), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_189), .A2(n_195), .B1(n_214), .B2(n_216), .Y(n_213) );
AND2x4_ASAP7_75t_L g189 ( .A(n_190), .B(n_193), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
NOR2x1p5_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_201), .A2(n_284), .B1(n_386), .B2(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_226), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_202), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_202), .B(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_211), .Y(n_202) );
INVx2_ASAP7_75t_L g249 ( .A(n_203), .Y(n_249) );
OR2x2_ASAP7_75t_L g253 ( .A(n_203), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_203), .B(n_266), .Y(n_271) );
AND2x4_ASAP7_75t_SL g281 ( .A(n_203), .B(n_212), .Y(n_281) );
OR2x2_ASAP7_75t_L g288 ( .A(n_203), .B(n_228), .Y(n_288) );
OR2x2_ASAP7_75t_L g300 ( .A(n_203), .B(n_212), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_203), .B(n_228), .Y(n_314) );
INVx1_ASAP7_75t_L g319 ( .A(n_203), .Y(n_319) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_203), .Y(n_337) );
AND2x2_ASAP7_75t_L g400 ( .A(n_203), .B(n_320), .Y(n_400) );
INVx2_ASAP7_75t_L g404 ( .A(n_203), .Y(n_404) );
OR2x2_ASAP7_75t_L g411 ( .A(n_203), .B(n_301), .Y(n_411) );
OR2x2_ASAP7_75t_L g433 ( .A(n_203), .B(n_434), .Y(n_433) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_210), .Y(n_203) );
AND2x2_ASAP7_75t_L g250 ( .A(n_211), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_211), .B(n_234), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_211), .B(n_310), .Y(n_372) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g269 ( .A(n_212), .Y(n_269) );
AND2x4_ASAP7_75t_L g320 ( .A(n_212), .B(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_212), .B(n_265), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_212), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_212), .B(n_254), .Y(n_413) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_218), .Y(n_212) );
INVx3_ASAP7_75t_L g481 ( .A(n_221), .Y(n_481) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AOI21x1_ASAP7_75t_L g235 ( .A1(n_222), .A2(n_236), .B(n_242), .Y(n_235) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_222), .A2(n_464), .B(n_470), .Y(n_463) );
AND2x2_ASAP7_75t_L g280 ( .A(n_226), .B(n_281), .Y(n_280) );
AO221x1_ASAP7_75t_L g354 ( .A1(n_226), .A2(n_269), .B1(n_300), .B2(n_355), .C(n_356), .Y(n_354) );
OAI322xp33_ASAP7_75t_L g406 ( .A1(n_226), .A2(n_326), .A3(n_407), .B1(n_409), .B2(n_410), .C1(n_411), .C2(n_412), .Y(n_406) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_234), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
BUFx3_ASAP7_75t_L g248 ( .A(n_228), .Y(n_248) );
INVx2_ASAP7_75t_L g254 ( .A(n_228), .Y(n_254) );
AND2x2_ASAP7_75t_L g266 ( .A(n_228), .B(n_234), .Y(n_266) );
INVx1_ASAP7_75t_L g311 ( .A(n_228), .Y(n_311) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_228), .Y(n_367) );
INVx1_ASAP7_75t_L g251 ( .A(n_234), .Y(n_251) );
OR2x2_ASAP7_75t_L g301 ( .A(n_234), .B(n_254), .Y(n_301) );
INVx2_ASAP7_75t_L g321 ( .A(n_234), .Y(n_321) );
INVx1_ASAP7_75t_L g374 ( .A(n_234), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_234), .B(n_404), .Y(n_403) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_241), .Y(n_236) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OAI21xp33_ASAP7_75t_SL g244 ( .A1(n_245), .A2(n_252), .B(n_255), .Y(n_244) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_245), .A2(n_284), .B1(n_286), .B2(n_290), .C(n_291), .Y(n_283) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_250), .Y(n_246) );
NOR2x1p5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g370 ( .A(n_249), .Y(n_370) );
INVx1_ASAP7_75t_SL g289 ( .A(n_250), .Y(n_289) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_250), .A2(n_395), .B(n_397), .Y(n_394) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_251), .Y(n_294) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_254), .Y(n_357) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
OAI211xp5_ASAP7_75t_L g332 ( .A1(n_257), .A2(n_333), .B(n_338), .C(n_349), .Y(n_332) );
OR2x2_ASAP7_75t_L g422 ( .A(n_257), .B(n_327), .Y(n_422) );
AND2x2_ASAP7_75t_L g424 ( .A(n_257), .B(n_290), .Y(n_424) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g264 ( .A(n_258), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g326 ( .A(n_258), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g364 ( .A(n_258), .B(n_331), .Y(n_364) );
OA33x2_ASAP7_75t_L g371 ( .A1(n_258), .A2(n_288), .A3(n_372), .B1(n_373), .B2(n_375), .B3(n_377), .Y(n_371) );
OR2x2_ASAP7_75t_L g382 ( .A(n_258), .B(n_367), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_258), .B(n_306), .Y(n_396) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g284 ( .A(n_260), .B(n_285), .Y(n_284) );
AOI22xp33_ASAP7_75t_SL g333 ( .A1(n_260), .A2(n_290), .B1(n_334), .B2(n_335), .Y(n_333) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_261), .B(n_341), .C(n_374), .Y(n_373) );
AOI322xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_267), .A3(n_269), .B1(n_270), .B2(n_272), .C1(n_276), .C2(n_280), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g369 ( .A(n_265), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_266), .A2(n_281), .B(n_325), .C(n_328), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_267), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
NAND4xp25_ASAP7_75t_SL g388 ( .A(n_268), .B(n_297), .C(n_389), .D(n_391), .Y(n_388) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx2_ASAP7_75t_L g278 ( .A(n_273), .Y(n_278) );
OR2x2_ASAP7_75t_L g323 ( .A(n_273), .B(n_275), .Y(n_323) );
AND2x2_ASAP7_75t_L g392 ( .A(n_274), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g397 ( .A(n_278), .B(n_392), .Y(n_397) );
BUFx2_ASAP7_75t_L g390 ( .A(n_279), .Y(n_390) );
INVx1_ASAP7_75t_SL g420 ( .A(n_280), .Y(n_420) );
AND2x4_ASAP7_75t_L g356 ( .A(n_281), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g409 ( .A(n_281), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g282 ( .A(n_283), .B(n_302), .C(n_324), .Y(n_282) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_SL g346 ( .A(n_288), .Y(n_346) );
OAI211xp5_ASAP7_75t_L g414 ( .A1(n_288), .A2(n_415), .B(n_416), .C(n_425), .Y(n_414) );
OR2x2_ASAP7_75t_L g336 ( .A(n_289), .B(n_337), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .B1(n_298), .B2(n_299), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_293), .B(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_296), .B(n_353), .Y(n_435) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g410 ( .A(n_297), .B(n_298), .Y(n_410) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g355 ( .A(n_301), .Y(n_355) );
AOI222xp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_307), .B1(n_312), .B2(n_316), .C1(n_317), .C2(n_322), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_305), .Y(n_316) );
AND2x2_ASAP7_75t_L g363 ( .A(n_306), .B(n_364), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_306), .A2(n_379), .B1(n_384), .B2(n_388), .Y(n_378) );
INVx2_ASAP7_75t_SL g431 ( .A(n_306), .Y(n_431) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g387 ( .A(n_311), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_311), .B(n_374), .Y(n_434) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g347 ( .A(n_315), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_317), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g385 ( .A(n_319), .Y(n_385) );
AND2x2_ASAP7_75t_SL g386 ( .A(n_320), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g428 ( .A(n_320), .B(n_357), .Y(n_428) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g353 ( .A(n_327), .Y(n_353) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g432 ( .A(n_330), .Y(n_432) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_331), .Y(n_376) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_343), .B(n_345), .C(n_348), .Y(n_338) );
AND2x2_ASAP7_75t_SL g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g383 ( .A(n_345), .Y(n_383) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_354), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_352), .B(n_353), .Y(n_351) );
NOR3xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_398), .C(n_414), .Y(n_358) );
NAND3xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_378), .C(n_394), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI221xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B1(n_368), .B2(n_369), .C(n_371), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_380), .B(n_383), .Y(n_379) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g407 ( .A(n_393), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g415 ( .A(n_397), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_405), .Y(n_398) );
INVx2_ASAP7_75t_L g421 ( .A(n_400), .Y(n_421) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g412 ( .A(n_403), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B1(n_421), .B2(n_422), .C(n_423), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_429), .B1(n_433), .B2(n_435), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_SL g730 ( .A(n_436), .Y(n_730) );
CKINVDCx11_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
OAI21x1_ASAP7_75t_SL g729 ( .A1(n_438), .A2(n_730), .B(n_731), .Y(n_729) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_440), .B(n_637), .Y(n_439) );
NOR3xp33_ASAP7_75t_SL g440 ( .A(n_441), .B(n_560), .C(n_595), .Y(n_440) );
OAI211xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_471), .B(n_522), .C(n_550), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_453), .Y(n_443) );
AND2x2_ASAP7_75t_L g543 ( .A(n_444), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_444), .B(n_549), .Y(n_583) );
AND2x2_ASAP7_75t_L g608 ( .A(n_444), .B(n_563), .Y(n_608) );
INVx4_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g525 ( .A(n_445), .Y(n_525) );
OR2x2_ASAP7_75t_L g546 ( .A(n_445), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g554 ( .A(n_445), .B(n_463), .Y(n_554) );
AND2x2_ASAP7_75t_L g562 ( .A(n_445), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g589 ( .A(n_445), .B(n_590), .Y(n_589) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_445), .B(n_592), .Y(n_600) );
AND2x4_ASAP7_75t_L g617 ( .A(n_445), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g655 ( .A(n_445), .Y(n_655) );
AND2x4_ASAP7_75t_SL g660 ( .A(n_445), .B(n_454), .Y(n_660) );
OR2x6_ASAP7_75t_L g445 ( .A(n_446), .B(n_452), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_453), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_453), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_463), .Y(n_453) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_454), .Y(n_555) );
INVx2_ASAP7_75t_L g591 ( .A(n_454), .Y(n_591) );
INVx1_ASAP7_75t_L g618 ( .A(n_454), .Y(n_618) );
AND2x2_ASAP7_75t_L g717 ( .A(n_454), .B(n_627), .Y(n_717) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_455), .Y(n_549) );
AND2x2_ASAP7_75t_L g563 ( .A(n_455), .B(n_463), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
INVx2_ASAP7_75t_L g592 ( .A(n_463), .Y(n_592) );
INVx2_ASAP7_75t_L g627 ( .A(n_463), .Y(n_627) );
OR2x2_ASAP7_75t_L g712 ( .A(n_463), .B(n_544), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_469), .Y(n_464) );
AOI211xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_489), .B(n_509), .C(n_516), .Y(n_471) );
INVx2_ASAP7_75t_SL g601 ( .A(n_472), .Y(n_601) );
AND2x2_ASAP7_75t_L g607 ( .A(n_472), .B(n_490), .Y(n_607) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_480), .Y(n_472) );
INVx1_ASAP7_75t_L g513 ( .A(n_473), .Y(n_513) );
INVx1_ASAP7_75t_L g519 ( .A(n_473), .Y(n_519) );
INVx2_ASAP7_75t_L g534 ( .A(n_473), .Y(n_534) );
AND2x2_ASAP7_75t_L g558 ( .A(n_473), .B(n_492), .Y(n_558) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_473), .Y(n_587) );
OR2x2_ASAP7_75t_L g667 ( .A(n_473), .B(n_500), .Y(n_667) );
AND2x2_ASAP7_75t_L g533 ( .A(n_480), .B(n_534), .Y(n_533) );
NOR2x1_ASAP7_75t_SL g565 ( .A(n_480), .B(n_500), .Y(n_565) );
AO21x1_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_482), .B(n_488), .Y(n_480) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_481), .A2(n_482), .B(n_488), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g579 ( .A(n_490), .B(n_512), .Y(n_579) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_500), .Y(n_490) );
OR2x2_ASAP7_75t_L g521 ( .A(n_491), .B(n_500), .Y(n_521) );
BUFx2_ASAP7_75t_L g535 ( .A(n_491), .Y(n_535) );
NOR2xp67_ASAP7_75t_L g586 ( .A(n_491), .B(n_587), .Y(n_586) );
INVx4_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_492), .Y(n_538) );
AND2x2_ASAP7_75t_L g564 ( .A(n_492), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g574 ( .A(n_492), .Y(n_574) );
NAND2x1_ASAP7_75t_L g612 ( .A(n_492), .B(n_500), .Y(n_612) );
OR2x2_ASAP7_75t_L g687 ( .A(n_492), .B(n_514), .Y(n_687) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx2_ASAP7_75t_SL g510 ( .A(n_500), .Y(n_510) );
AND2x2_ASAP7_75t_L g559 ( .A(n_500), .B(n_514), .Y(n_559) );
AND2x2_ASAP7_75t_L g630 ( .A(n_500), .B(n_631), .Y(n_630) );
BUFx2_ASAP7_75t_L g651 ( .A(n_500), .Y(n_651) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_508), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g573 ( .A(n_512), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
BUFx2_ASAP7_75t_L g568 ( .A(n_513), .Y(n_568) );
AND2x2_ASAP7_75t_L g540 ( .A(n_514), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g631 ( .A(n_514), .Y(n_631) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
OR2x2_ASAP7_75t_L g577 ( .A(n_518), .B(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_SL g619 ( .A(n_518), .B(n_620), .Y(n_619) );
AOI322xp5_ASAP7_75t_L g656 ( .A1(n_518), .A2(n_535), .A3(n_657), .B1(n_659), .B2(n_662), .C1(n_664), .C2(n_666), .Y(n_656) );
AND2x2_ASAP7_75t_L g721 ( .A(n_518), .B(n_722), .Y(n_721) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_519), .B(n_535), .Y(n_545) );
AOI322xp5_ASAP7_75t_L g596 ( .A1(n_520), .A2(n_597), .A3(n_601), .B1(n_602), .B2(n_605), .C1(n_607), .C2(n_608), .Y(n_596) );
INVx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g648 ( .A(n_521), .B(n_601), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_521), .A2(n_708), .B1(n_710), .B2(n_713), .Y(n_707) );
OR2x2_ASAP7_75t_L g725 ( .A(n_521), .B(n_674), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_535), .B(n_536), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_526), .Y(n_523) );
AOI221xp5_ASAP7_75t_SL g575 ( .A1(n_524), .A2(n_551), .B1(n_576), .B2(n_579), .C(n_580), .Y(n_575) );
AND2x2_ASAP7_75t_L g602 ( .A(n_524), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_525), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g644 ( .A(n_525), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g673 ( .A(n_526), .Y(n_673) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_533), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_527), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g615 ( .A(n_527), .Y(n_615) );
OR2x2_ASAP7_75t_L g622 ( .A(n_527), .B(n_623), .Y(n_622) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g665 ( .A(n_528), .B(n_627), .Y(n_665) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
AND2x4_ASAP7_75t_L g544 ( .A(n_529), .B(n_530), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_533), .B(n_594), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_533), .B(n_574), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_533), .Y(n_674) );
INVx1_ASAP7_75t_L g541 ( .A(n_534), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_542), .B1(n_545), .B2(n_546), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_SL g652 ( .A(n_540), .Y(n_652) );
AND2x2_ASAP7_75t_L g709 ( .A(n_541), .B(n_565), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_543), .B(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_SL g581 ( .A(n_543), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_543), .B(n_702), .Y(n_701) );
BUFx3_ASAP7_75t_L g569 ( .A(n_544), .Y(n_569) );
INVx2_ASAP7_75t_L g599 ( .A(n_544), .Y(n_599) );
AND2x2_ASAP7_75t_L g642 ( .A(n_544), .B(n_626), .Y(n_642) );
INVx1_ASAP7_75t_L g556 ( .A(n_546), .Y(n_556) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI21xp5_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_556), .B(n_557), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g635 ( .A(n_554), .Y(n_635) );
INVx2_ASAP7_75t_L g623 ( .A(n_555), .Y(n_623) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x2_ASAP7_75t_L g620 ( .A(n_559), .B(n_574), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_559), .A2(n_657), .B(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_561), .B(n_575), .Y(n_560) );
AOI32xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_564), .A3(n_566), .B1(n_570), .B2(n_573), .Y(n_561) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_562), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_562), .A2(n_651), .B1(n_669), .B2(n_671), .C(n_677), .Y(n_668) );
AND2x2_ASAP7_75t_L g688 ( .A(n_562), .B(n_569), .Y(n_688) );
BUFx2_ASAP7_75t_L g572 ( .A(n_563), .Y(n_572) );
INVx1_ASAP7_75t_L g697 ( .A(n_563), .Y(n_697) );
INVx1_ASAP7_75t_L g702 ( .A(n_563), .Y(n_702) );
INVx1_ASAP7_75t_SL g695 ( .A(n_564), .Y(n_695) );
INVx2_ASAP7_75t_L g578 ( .A(n_565), .Y(n_578) );
AND2x2_ASAP7_75t_L g690 ( .A(n_566), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g662 ( .A(n_568), .B(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g634 ( .A(n_569), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_569), .B(n_660), .Y(n_682) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g594 ( .A(n_574), .Y(n_594) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g584 ( .A(n_578), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g593 ( .A(n_578), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g698 ( .A(n_579), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_584), .B1(n_588), .B2(n_593), .Y(n_580) );
INVx2_ASAP7_75t_SL g672 ( .A(n_582), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_582), .B(n_711), .Y(n_713) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_584), .A2(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g629 ( .A(n_586), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g657 ( .A(n_589), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g604 ( .A(n_590), .Y(n_604) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g646 ( .A(n_592), .Y(n_646) );
INVx1_ASAP7_75t_L g691 ( .A(n_593), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_609), .C(n_632), .Y(n_595) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx2_ASAP7_75t_L g658 ( .A(n_598), .Y(n_658) );
AND2x2_ASAP7_75t_L g676 ( .A(n_598), .B(n_617), .Y(n_676) );
OR2x2_ASAP7_75t_L g715 ( .A(n_598), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_599), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g611 ( .A(n_601), .B(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g678 ( .A(n_604), .B(n_615), .Y(n_678) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_607), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g719 ( .A(n_607), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_613), .B1(n_617), .B2(n_619), .C(n_621), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_610), .A2(n_633), .B(n_636), .Y(n_632) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx3_ASAP7_75t_L g663 ( .A(n_612), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_612), .B(n_706), .Y(n_705) );
INVxp33_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g624 ( .A(n_620), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_625), .B2(n_628), .Y(n_621) );
INVx2_ASAP7_75t_L g727 ( .A(n_623), .Y(n_727) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVxp67_ASAP7_75t_L g706 ( .A(n_631), .Y(n_706) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
NOR2x1_ASAP7_75t_L g637 ( .A(n_638), .B(n_683), .Y(n_637) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_639), .B(n_656), .C(n_668), .D(n_680), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_643), .B(n_647), .C(n_649), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g679 ( .A(n_642), .Y(n_679) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_644), .A2(n_650), .B(n_653), .Y(n_649) );
INVx2_ASAP7_75t_L g728 ( .A(n_645), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_646), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g661 ( .A(n_646), .Y(n_661) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
OR2x2_ASAP7_75t_L g723 ( .A(n_651), .B(n_687), .Y(n_723) );
INVxp67_ASAP7_75t_SL g694 ( .A(n_658), .Y(n_694) );
AND2x2_ASAP7_75t_SL g659 ( .A(n_660), .B(n_661), .Y(n_659) );
AND2x2_ASAP7_75t_L g664 ( .A(n_660), .B(n_665), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_660), .A2(n_690), .B(n_692), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_660), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_SL g718 ( .A(n_660), .Y(n_718) );
INVxp67_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI22xp33_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND4xp25_ASAP7_75t_L g683 ( .A(n_684), .B(n_689), .C(n_699), .D(n_720), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .B1(n_696), .B2(n_698), .Y(n_692) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI211xp5_ASAP7_75t_SL g699 ( .A1(n_700), .A2(n_703), .B(n_707), .C(n_714), .Y(n_699) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_718), .B(n_719), .Y(n_714) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
OAI21xp5_ASAP7_75t_SL g720 ( .A1(n_721), .A2(n_724), .B(n_726), .Y(n_720) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
BUFx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx3_ASAP7_75t_L g753 ( .A(n_736), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
BUFx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx2_ASAP7_75t_L g758 ( .A(n_751), .Y(n_758) );
INVx2_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
endmodule