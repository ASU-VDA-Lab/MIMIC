module fake_jpeg_9819_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_48),
.B1(n_17),
.B2(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_47),
.Y(n_56)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_95)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_26),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_78),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_17),
.B1(n_33),
.B2(n_38),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_74),
.B1(n_91),
.B2(n_95),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_17),
.B1(n_38),
.B2(n_48),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_80),
.B(n_86),
.Y(n_118)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_94),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_47),
.B1(n_33),
.B2(n_32),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_47),
.B1(n_40),
.B2(n_36),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_67),
.B1(n_62),
.B2(n_61),
.Y(n_112)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_62),
.B1(n_56),
.B2(n_40),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_96),
.B1(n_78),
.B2(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_88),
.B1(n_23),
.B2(n_24),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_115),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_63),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_125),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_83),
.B(n_21),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_128),
.C(n_24),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_72),
.Y(n_122)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_56),
.B1(n_21),
.B2(n_23),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_29),
.B1(n_114),
.B2(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_22),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_28),
.C(n_30),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_93),
.B1(n_99),
.B2(n_26),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_142),
.B(n_146),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_146),
.B(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_104),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_140),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_143),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_75),
.C(n_77),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_152),
.C(n_30),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_84),
.B1(n_85),
.B2(n_79),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_139),
.A2(n_141),
.B1(n_148),
.B2(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_92),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_85),
.B1(n_79),
.B2(n_89),
.Y(n_141)
);

NOR2x1p5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_30),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_36),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_24),
.B(n_22),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_151),
.B1(n_154),
.B2(n_114),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_88),
.B1(n_26),
.B2(n_29),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_112),
.B1(n_103),
.B2(n_128),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_28),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_36),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_120),
.A2(n_30),
.B(n_35),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_30),
.B(n_102),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_100),
.A2(n_36),
.A3(n_35),
.B1(n_34),
.B2(n_31),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_116),
.B(n_30),
.Y(n_185)
);

OAI22x1_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_157),
.B1(n_130),
.B2(n_155),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_159),
.A2(n_164),
.B1(n_185),
.B2(n_0),
.Y(n_207)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_171),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_166),
.B1(n_174),
.B2(n_178),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_113),
.B1(n_34),
.B2(n_31),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_165),
.B(n_170),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_145),
.B1(n_129),
.B2(n_142),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_15),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_167),
.B(n_3),
.Y(n_221)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_143),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_113),
.B1(n_101),
.B2(n_31),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_177),
.B1(n_179),
.B2(n_181),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_107),
.B1(n_127),
.B2(n_101),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_148),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_107),
.B1(n_127),
.B2(n_124),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_150),
.A2(n_35),
.B1(n_100),
.B2(n_124),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_135),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_126),
.B(n_30),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_190),
.Y(n_198)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_187),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_137),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_131),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_15),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_132),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_1),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_149),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_149),
.A3(n_132),
.B1(n_144),
.B2(n_16),
.C1(n_14),
.C2(n_13),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g235 ( 
.A1(n_193),
.A2(n_176),
.B(n_161),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_194),
.B(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_190),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_204),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_144),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_213),
.C(n_183),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_16),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_202),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_16),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_14),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_211),
.B(n_178),
.Y(n_238)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_217),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_159),
.A2(n_13),
.B1(n_12),
.B2(n_2),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_12),
.C(n_1),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_221),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_0),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_185),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_167),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_189),
.B1(n_169),
.B2(n_162),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_160),
.B1(n_180),
.B2(n_165),
.Y(n_224)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_213),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_205),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_168),
.B1(n_170),
.B2(n_163),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_236),
.B1(n_211),
.B2(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_239),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_235),
.A2(n_238),
.B(n_240),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_168),
.B1(n_163),
.B2(n_186),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_219),
.B(n_195),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_175),
.B1(n_173),
.B2(n_176),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_246),
.B1(n_214),
.B2(n_222),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_244),
.C(n_245),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_177),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_3),
.C(n_4),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_210),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_220),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_247),
.B(n_6),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_198),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_252),
.Y(n_277)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_255),
.C(n_258),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_205),
.C(n_199),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_209),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_256),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_207),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_207),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_209),
.C(n_210),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_207),
.C(n_212),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_246),
.Y(n_284)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_7),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_267),
.C(n_245),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_8),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_8),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_268),
.A2(n_233),
.B1(n_228),
.B2(n_230),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_287),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_248),
.B(n_240),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_279),
.B(n_261),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_248),
.B(n_223),
.Y(n_279)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_229),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_286),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_270),
.A2(n_233),
.B1(n_229),
.B2(n_230),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_253),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_293),
.C(n_296),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_281),
.B(n_283),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_259),
.B1(n_258),
.B2(n_255),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_291),
.A2(n_297),
.B1(n_9),
.B2(n_10),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_254),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_292),
.B(n_295),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_254),
.C(n_250),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_277),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_276),
.C(n_279),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_272),
.A2(n_257),
.B1(n_266),
.B2(n_11),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_225),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_302),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_243),
.C(n_10),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_280),
.Y(n_303)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_303),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_273),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_304),
.A2(n_306),
.B(n_307),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_309),
.C(n_301),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_280),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_278),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_311),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_291),
.A2(n_278),
.B1(n_273),
.B2(n_275),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_11),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_296),
.B(n_11),
.CI(n_9),
.CON(n_312),
.SN(n_312)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_314),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_288),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_308),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_318),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_290),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_324),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_322),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_293),
.C(n_310),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_329),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_307),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_315),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_312),
.C(n_10),
.Y(n_333)
);

OAI321xp33_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_323),
.A3(n_305),
.B1(n_316),
.B2(n_312),
.C(n_313),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_331),
.B(n_328),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_326),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_333),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_327),
.Y(n_339)
);


endmodule