module fake_netlist_1_3194_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
OAI22xp5_ASAP7_75t_SL g11 ( .A1(n_7), .A2(n_10), .B1(n_4), .B2(n_0), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_4), .B(n_1), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_12), .B(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_13), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_14), .B(n_15), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_19), .B(n_16), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
BUFx2_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
OAI221xp5_ASAP7_75t_SL g25 ( .A1(n_23), .A2(n_11), .B1(n_21), .B2(n_19), .C(n_5), .Y(n_25) );
NAND2xp5_ASAP7_75t_SL g26 ( .A(n_24), .B(n_11), .Y(n_26) );
A2O1A1Ixp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_24), .B(n_21), .C(n_15), .Y(n_27) );
XNOR2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_1), .Y(n_28) );
NOR3xp33_ASAP7_75t_SL g29 ( .A(n_28), .B(n_2), .C(n_3), .Y(n_29) );
NOR2xp33_ASAP7_75t_L g30 ( .A(n_28), .B(n_2), .Y(n_30) );
AOI221xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_27), .B1(n_15), .B2(n_5), .C(n_8), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g33 ( .A(n_32), .Y(n_33) );
NAND2xp33_ASAP7_75t_L g34 ( .A(n_33), .B(n_31), .Y(n_34) );
endmodule