module real_aes_8971_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_532;
wire n_284;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_713;
wire n_735;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g508 ( .A(n_1), .Y(n_508) );
INVx1_ASAP7_75t_L g203 ( .A(n_2), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_3), .A2(n_37), .B1(n_175), .B2(n_517), .Y(n_516) );
AOI21xp33_ASAP7_75t_L g214 ( .A1(n_4), .A2(n_132), .B(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_5), .B(n_162), .Y(n_500) );
AND2x6_ASAP7_75t_L g137 ( .A(n_6), .B(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_7), .A2(n_183), .B(n_184), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_8), .B(n_38), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_9), .B(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g220 ( .A(n_10), .Y(n_220) );
INVx1_ASAP7_75t_L g158 ( .A(n_11), .Y(n_158) );
INVx1_ASAP7_75t_L g504 ( .A(n_12), .Y(n_504) );
INVx1_ASAP7_75t_L g191 ( .A(n_13), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_14), .B(n_206), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_15), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_16), .B(n_154), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_17), .A2(n_41), .B1(n_749), .B2(n_750), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_17), .Y(n_750) );
AO32x2_ASAP7_75t_L g514 ( .A1(n_18), .A2(n_153), .A3(n_162), .B1(n_486), .B2(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_19), .B(n_175), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_20), .B(n_148), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_21), .B(n_154), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_22), .A2(n_50), .B1(n_175), .B2(n_517), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_23), .B(n_132), .Y(n_131) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_24), .A2(n_76), .B1(n_175), .B2(n_206), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_25), .B(n_175), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_26), .B(n_213), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_27), .A2(n_188), .B(n_190), .C(n_192), .Y(n_187) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_28), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_29), .B(n_166), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_30), .B(n_173), .Y(n_204) );
INVx1_ASAP7_75t_L g230 ( .A(n_31), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_32), .B(n_166), .Y(n_530) );
INVx2_ASAP7_75t_L g135 ( .A(n_33), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_34), .B(n_175), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_35), .B(n_166), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_36), .A2(n_137), .B(n_140), .C(n_143), .Y(n_139) );
INVx1_ASAP7_75t_L g228 ( .A(n_39), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_40), .B(n_173), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_41), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_42), .A2(n_104), .B1(n_115), .B2(n_758), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_43), .B(n_175), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_44), .A2(n_87), .B1(n_151), .B2(n_517), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_45), .B(n_175), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_46), .B(n_175), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_47), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_48), .B(n_484), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_49), .B(n_132), .Y(n_176) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_51), .A2(n_60), .B1(n_175), .B2(n_206), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_52), .A2(n_140), .B1(n_206), .B2(n_227), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_53), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_54), .B(n_175), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g199 ( .A(n_55), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_56), .B(n_175), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_57), .A2(n_218), .B(n_219), .C(n_221), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_58), .Y(n_268) );
INVx1_ASAP7_75t_L g216 ( .A(n_59), .Y(n_216) );
INVx1_ASAP7_75t_L g138 ( .A(n_61), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_62), .B(n_175), .Y(n_509) );
INVx1_ASAP7_75t_L g157 ( .A(n_63), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_64), .Y(n_120) );
AO32x2_ASAP7_75t_L g550 ( .A1(n_65), .A2(n_162), .A3(n_165), .B1(n_486), .B2(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g482 ( .A(n_66), .Y(n_482) );
INVx1_ASAP7_75t_L g525 ( .A(n_67), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_SL g238 ( .A1(n_68), .A2(n_148), .B(n_221), .C(n_239), .Y(n_238) );
INVxp67_ASAP7_75t_L g240 ( .A(n_69), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_70), .B(n_206), .Y(n_526) );
INVx1_ASAP7_75t_L g107 ( .A(n_71), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_72), .Y(n_233) );
INVx1_ASAP7_75t_L g261 ( .A(n_73), .Y(n_261) );
OAI321xp33_ASAP7_75t_L g121 ( .A1(n_74), .A2(n_122), .A3(n_452), .B1(n_455), .B2(n_456), .C(n_458), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_74), .Y(n_455) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_75), .A2(n_89), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_75), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_77), .A2(n_137), .B(n_140), .C(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_78), .B(n_517), .Y(n_539) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_79), .A2(n_747), .B1(n_748), .B2(n_751), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_79), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_80), .B(n_206), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_81), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g155 ( .A(n_82), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_83), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_84), .B(n_206), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_85), .A2(n_137), .B(n_140), .C(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g110 ( .A(n_86), .Y(n_110) );
OR2x2_ASAP7_75t_L g454 ( .A(n_86), .B(n_111), .Y(n_454) );
OR2x2_ASAP7_75t_L g466 ( .A(n_86), .B(n_112), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_88), .A2(n_102), .B1(n_206), .B2(n_207), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_89), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_90), .B(n_166), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_91), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_92), .A2(n_137), .B(n_140), .C(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_93), .Y(n_178) );
INVx1_ASAP7_75t_L g237 ( .A(n_94), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_95), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_96), .B(n_145), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_97), .B(n_206), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_98), .B(n_162), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_99), .B(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_100), .A2(n_132), .B(n_236), .Y(n_235) );
AOI222xp33_ASAP7_75t_L g462 ( .A1(n_101), .A2(n_463), .B1(n_745), .B2(n_746), .C1(n_752), .C2(n_754), .Y(n_462) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g759 ( .A(n_105), .Y(n_759) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g753 ( .A(n_109), .Y(n_753) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g469 ( .A(n_110), .B(n_112), .Y(n_469) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_461), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g757 ( .A(n_119), .Y(n_757) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_122), .B(n_457), .Y(n_456) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_124), .B1(n_448), .B2(n_449), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_123), .A2(n_466), .B1(n_467), .B2(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_124), .A2(n_464), .B1(n_467), .B2(n_470), .Y(n_463) );
AND2x2_ASAP7_75t_SL g124 ( .A(n_125), .B(n_417), .Y(n_124) );
NOR3xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_310), .C(n_383), .Y(n_125) );
OAI211xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_195), .B(n_242), .C(n_294), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_163), .Y(n_128) );
AND2x2_ASAP7_75t_L g258 ( .A(n_129), .B(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g277 ( .A(n_129), .Y(n_277) );
INVx2_ASAP7_75t_L g292 ( .A(n_129), .Y(n_292) );
INVx1_ASAP7_75t_L g322 ( .A(n_129), .Y(n_322) );
AND2x2_ASAP7_75t_L g372 ( .A(n_129), .B(n_293), .Y(n_372) );
AOI32xp33_ASAP7_75t_L g399 ( .A1(n_129), .A2(n_327), .A3(n_400), .B1(n_402), .B2(n_403), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_129), .B(n_248), .Y(n_405) );
AND2x2_ASAP7_75t_L g432 ( .A(n_129), .B(n_275), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_129), .B(n_441), .Y(n_440) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_159), .Y(n_129) );
AOI21xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_139), .B(n_152), .Y(n_130) );
BUFx2_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_133), .B(n_137), .Y(n_200) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g484 ( .A(n_134), .Y(n_484) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx1_ASAP7_75t_L g207 ( .A(n_135), .Y(n_207) );
INVx1_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx3_ASAP7_75t_L g146 ( .A(n_136), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_136), .Y(n_148) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
INVx4_ASAP7_75t_SL g193 ( .A(n_137), .Y(n_193) );
BUFx3_ASAP7_75t_L g486 ( .A(n_137), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_137), .A2(n_493), .B(n_496), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_137), .A2(n_503), .B(n_507), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_137), .A2(n_524), .B(n_527), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_137), .A2(n_533), .B(n_537), .Y(n_532) );
INVx5_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx3_ASAP7_75t_L g151 ( .A(n_141), .Y(n_151) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
INVx1_ASAP7_75t_L g517 ( .A(n_141), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_147), .B(n_149), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_145), .A2(n_203), .B(n_204), .C(n_205), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_145), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_145), .A2(n_494), .B(n_495), .Y(n_493) );
INVx2_ASAP7_75t_L g499 ( .A(n_145), .Y(n_499) );
O2A1O1Ixp5_ASAP7_75t_SL g524 ( .A1(n_145), .A2(n_221), .B(n_525), .C(n_526), .Y(n_524) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_146), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_146), .B(n_240), .Y(n_239) );
OAI22xp5_ASAP7_75t_SL g551 ( .A1(n_146), .A2(n_173), .B1(n_552), .B2(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g536 ( .A(n_148), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_149), .A2(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g192 ( .A(n_151), .Y(n_192) );
INVx1_ASAP7_75t_L g266 ( .A(n_152), .Y(n_266) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_152), .A2(n_477), .B(n_487), .Y(n_476) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_152), .A2(n_502), .B(n_510), .Y(n_501) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_153), .A2(n_198), .B(n_208), .Y(n_197) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_153), .A2(n_225), .B(n_232), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_153), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_155), .B(n_156), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_SL g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx3_ASAP7_75t_L g213 ( .A(n_161), .Y(n_213) );
AO21x1_ASAP7_75t_L g562 ( .A1(n_161), .A2(n_563), .B(n_566), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_161), .B(n_486), .C(n_563), .Y(n_587) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_162), .A2(n_235), .B(n_241), .Y(n_234) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_162), .A2(n_492), .B(n_500), .Y(n_491) );
AND2x2_ASAP7_75t_L g321 ( .A(n_163), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g343 ( .A(n_163), .Y(n_343) );
AND2x2_ASAP7_75t_L g428 ( .A(n_163), .B(n_258), .Y(n_428) );
AND2x2_ASAP7_75t_L g431 ( .A(n_163), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_180), .Y(n_163) );
INVx2_ASAP7_75t_L g250 ( .A(n_164), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_164), .B(n_275), .Y(n_281) );
AND2x2_ASAP7_75t_L g291 ( .A(n_164), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g327 ( .A(n_164), .Y(n_327) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_167), .B(n_177), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g179 ( .A(n_166), .Y(n_179) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_166), .A2(n_182), .B(n_194), .Y(n_181) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_166), .A2(n_523), .B(n_530), .Y(n_522) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_166), .A2(n_532), .B(n_540), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_176), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_174), .Y(n_169) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g218 ( .A(n_173), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_173), .A2(n_499), .B1(n_516), .B2(n_518), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_173), .A2(n_499), .B1(n_564), .B2(n_565), .Y(n_563) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g221 ( .A(n_175), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_179), .B(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_179), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g269 ( .A(n_180), .B(n_250), .Y(n_269) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g251 ( .A(n_181), .Y(n_251) );
AND2x2_ASAP7_75t_L g293 ( .A(n_181), .B(n_275), .Y(n_293) );
AND2x2_ASAP7_75t_L g362 ( .A(n_181), .B(n_259), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .C(n_193), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_186), .A2(n_193), .B(n_216), .C(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_186), .A2(n_193), .B(n_237), .C(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_188), .B(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g506 ( .A(n_188), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_188), .A2(n_528), .B(n_529), .Y(n_527) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OAI22xp5_ASAP7_75t_SL g227 ( .A1(n_189), .A2(n_228), .B1(n_229), .B2(n_230), .Y(n_227) );
INVx2_ASAP7_75t_L g229 ( .A(n_189), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g225 ( .A1(n_193), .A2(n_200), .B1(n_226), .B2(n_231), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_210), .Y(n_195) );
OR2x2_ASAP7_75t_L g256 ( .A(n_196), .B(n_224), .Y(n_256) );
INVx1_ASAP7_75t_L g335 ( .A(n_196), .Y(n_335) );
AND2x2_ASAP7_75t_L g349 ( .A(n_196), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_196), .B(n_223), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_196), .B(n_347), .Y(n_401) );
AND2x2_ASAP7_75t_L g409 ( .A(n_196), .B(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx3_ASAP7_75t_L g246 ( .A(n_197), .Y(n_246) );
AND2x2_ASAP7_75t_L g316 ( .A(n_197), .B(n_224), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_200), .A2(n_261), .B(n_262), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_205), .A2(n_504), .B(n_505), .C(n_506), .Y(n_503) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_210), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g443 ( .A(n_210), .Y(n_443) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_223), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_211), .B(n_287), .Y(n_309) );
OR2x2_ASAP7_75t_L g338 ( .A(n_211), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g370 ( .A(n_211), .B(n_350), .Y(n_370) );
INVx1_ASAP7_75t_SL g390 ( .A(n_211), .Y(n_390) );
AND2x2_ASAP7_75t_L g394 ( .A(n_211), .B(n_255), .Y(n_394) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_SL g247 ( .A(n_212), .B(n_223), .Y(n_247) );
AND2x2_ASAP7_75t_L g254 ( .A(n_212), .B(n_234), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_212), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g297 ( .A(n_212), .B(n_279), .Y(n_297) );
INVx1_ASAP7_75t_SL g304 ( .A(n_212), .Y(n_304) );
BUFx2_ASAP7_75t_L g315 ( .A(n_212), .Y(n_315) );
AND2x2_ASAP7_75t_L g331 ( .A(n_212), .B(n_246), .Y(n_331) );
AND2x2_ASAP7_75t_L g346 ( .A(n_212), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g410 ( .A(n_212), .B(n_224), .Y(n_410) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_222), .Y(n_212) );
O2A1O1Ixp5_ASAP7_75t_L g481 ( .A1(n_218), .A2(n_482), .B(n_483), .C(n_485), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_218), .A2(n_538), .B(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_223), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g334 ( .A(n_223), .B(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_223), .A2(n_352), .B1(n_355), .B2(n_358), .C(n_363), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_223), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_234), .Y(n_223) );
INVx3_ASAP7_75t_L g279 ( .A(n_224), .Y(n_279) );
BUFx2_ASAP7_75t_L g289 ( .A(n_234), .Y(n_289) );
AND2x2_ASAP7_75t_L g303 ( .A(n_234), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g320 ( .A(n_234), .Y(n_320) );
OR2x2_ASAP7_75t_L g339 ( .A(n_234), .B(n_279), .Y(n_339) );
INVx3_ASAP7_75t_L g347 ( .A(n_234), .Y(n_347) );
AND2x2_ASAP7_75t_L g350 ( .A(n_234), .B(n_279), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_248), .B1(n_252), .B2(n_257), .C(n_270), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_245), .B(n_319), .Y(n_444) );
OR2x2_ASAP7_75t_L g447 ( .A(n_245), .B(n_278), .Y(n_447) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
OAI221xp5_ASAP7_75t_SL g270 ( .A1(n_246), .A2(n_271), .B1(n_278), .B2(n_280), .C(n_283), .Y(n_270) );
AND2x2_ASAP7_75t_L g287 ( .A(n_246), .B(n_279), .Y(n_287) );
AND2x2_ASAP7_75t_L g295 ( .A(n_246), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_246), .B(n_303), .Y(n_302) );
NAND2x1_ASAP7_75t_L g345 ( .A(n_246), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g397 ( .A(n_246), .B(n_339), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_248), .A2(n_357), .B1(n_386), .B2(n_388), .Y(n_385) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI322xp5_ASAP7_75t_L g294 ( .A1(n_249), .A2(n_258), .A3(n_295), .B1(n_298), .B2(n_301), .C1(n_305), .C2(n_308), .Y(n_294) );
OR2x2_ASAP7_75t_L g306 ( .A(n_249), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_250), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g285 ( .A(n_250), .B(n_259), .Y(n_285) );
INVx1_ASAP7_75t_L g300 ( .A(n_250), .Y(n_300) );
AND2x2_ASAP7_75t_L g366 ( .A(n_250), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g276 ( .A(n_251), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g367 ( .A(n_251), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_251), .B(n_275), .Y(n_441) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_255), .B(n_390), .Y(n_389) );
INVx3_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g341 ( .A(n_256), .B(n_288), .Y(n_341) );
OR2x2_ASAP7_75t_L g438 ( .A(n_256), .B(n_289), .Y(n_438) );
INVx1_ASAP7_75t_L g419 ( .A(n_257), .Y(n_419) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_269), .Y(n_257) );
INVx4_ASAP7_75t_L g307 ( .A(n_258), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_258), .B(n_326), .Y(n_332) );
INVx2_ASAP7_75t_L g275 ( .A(n_259), .Y(n_275) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_266), .B(n_267), .Y(n_259) );
INVx1_ASAP7_75t_L g357 ( .A(n_269), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_269), .B(n_329), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g344 ( .A1(n_271), .A2(n_345), .B(n_348), .Y(n_344) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g329 ( .A(n_275), .Y(n_329) );
INVx1_ASAP7_75t_L g356 ( .A(n_275), .Y(n_356) );
INVx1_ASAP7_75t_L g282 ( .A(n_276), .Y(n_282) );
AND2x2_ASAP7_75t_L g284 ( .A(n_276), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g380 ( .A(n_277), .B(n_366), .Y(n_380) );
AND2x2_ASAP7_75t_L g402 ( .A(n_277), .B(n_362), .Y(n_402) );
BUFx2_ASAP7_75t_L g354 ( .A(n_279), .Y(n_354) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AOI32xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_286), .A3(n_287), .B1(n_288), .B2(n_290), .Y(n_283) );
INVx1_ASAP7_75t_L g364 ( .A(n_284), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_284), .A2(n_412), .B1(n_413), .B2(n_415), .Y(n_411) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_287), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_287), .B(n_346), .Y(n_387) );
AND2x2_ASAP7_75t_L g434 ( .A(n_287), .B(n_319), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_288), .B(n_335), .Y(n_382) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g435 ( .A(n_290), .Y(n_435) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g360 ( .A(n_291), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_293), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g407 ( .A(n_293), .B(n_327), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_293), .B(n_322), .Y(n_414) );
INVx1_ASAP7_75t_SL g396 ( .A(n_295), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_296), .B(n_347), .Y(n_374) );
NOR4xp25_ASAP7_75t_L g420 ( .A(n_296), .B(n_319), .C(n_421), .D(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_297), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVxp67_ASAP7_75t_L g377 ( .A(n_300), .Y(n_377) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI21xp33_ASAP7_75t_L g427 ( .A1(n_303), .A2(n_394), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g319 ( .A(n_304), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g368 ( .A(n_307), .Y(n_368) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND4xp25_ASAP7_75t_SL g310 ( .A(n_311), .B(n_336), .C(n_351), .D(n_371), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_317), .B(n_321), .C(n_323), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g403 ( .A(n_316), .B(n_346), .Y(n_403) );
AND2x2_ASAP7_75t_L g412 ( .A(n_316), .B(n_390), .Y(n_412) );
INVx3_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_319), .B(n_354), .Y(n_416) );
AND2x2_ASAP7_75t_L g328 ( .A(n_322), .B(n_329), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_330), .B1(n_332), .B2(n_333), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g426 ( .A(n_326), .B(n_372), .Y(n_426) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_328), .B(n_377), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_329), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .B(n_342), .C(n_344), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_337), .A2(n_372), .B1(n_373), .B2(n_375), .C(n_378), .Y(n_371) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_345), .A2(n_430), .B1(n_433), .B2(n_435), .C(n_436), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_346), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_354), .B(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g384 ( .A(n_356), .Y(n_384) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_359), .A2(n_379), .B1(n_381), .B2(n_382), .Y(n_378) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI21xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B(n_369), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_368), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g442 ( .A1(n_379), .A2(n_405), .B1(n_443), .B2(n_444), .C(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g424 ( .A(n_381), .Y(n_424) );
OAI211xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_385), .B(n_391), .C(n_411), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI211xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_395), .C(n_404), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
A2O1A1Ixp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_398), .C(n_399), .Y(n_395) );
INVx1_ASAP7_75t_L g423 ( .A(n_401), .Y(n_423) );
OAI21xp5_ASAP7_75t_SL g445 ( .A1(n_402), .A2(n_428), .B(n_446), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B(n_408), .Y(n_404) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI21xp5_ASAP7_75t_SL g437 ( .A1(n_414), .A2(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_429), .C(n_442), .Y(n_417) );
OAI211xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_425), .C(n_427), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
CKINVDCx14_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g457 ( .A(n_454), .Y(n_457) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_454), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_458), .B(n_462), .C(n_756), .Y(n_461) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g755 ( .A(n_470), .Y(n_755) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR3x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_673), .C(n_722), .Y(n_471) );
NAND5xp2_ASAP7_75t_L g472 ( .A(n_473), .B(n_588), .C(n_616), .D(n_646), .E(n_660), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_511), .B1(n_541), .B2(n_546), .C(n_555), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_488), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_475), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g568 ( .A(n_476), .Y(n_568) );
AND2x2_ASAP7_75t_L g576 ( .A(n_476), .B(n_491), .Y(n_576) );
AND2x2_ASAP7_75t_L g599 ( .A(n_476), .B(n_490), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_476), .B(n_501), .Y(n_614) );
OR2x2_ASAP7_75t_L g623 ( .A(n_476), .B(n_562), .Y(n_623) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_476), .Y(n_626) );
AND2x2_ASAP7_75t_L g734 ( .A(n_476), .B(n_562), .Y(n_734) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_481), .B(n_486), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_483), .A2(n_499), .B(n_508), .C(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_488), .B(n_626), .Y(n_682) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
OAI311xp33_ASAP7_75t_L g624 ( .A1(n_489), .A2(n_625), .A3(n_626), .B1(n_627), .C1(n_642), .Y(n_624) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_501), .Y(n_489) );
AND2x2_ASAP7_75t_L g585 ( .A(n_490), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g592 ( .A(n_490), .Y(n_592) );
AND2x2_ASAP7_75t_L g713 ( .A(n_490), .B(n_545), .Y(n_713) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_491), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g569 ( .A(n_491), .B(n_501), .Y(n_569) );
AND2x2_ASAP7_75t_L g621 ( .A(n_491), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g635 ( .A(n_491), .B(n_568), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_499), .Y(n_496) );
INVx2_ASAP7_75t_L g545 ( .A(n_501), .Y(n_545) );
AND2x2_ASAP7_75t_L g584 ( .A(n_501), .B(n_568), .Y(n_584) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_519), .Y(n_511) );
OR2x2_ASAP7_75t_L g679 ( .A(n_512), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_512), .B(n_685), .Y(n_696) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_513), .B(n_692), .Y(n_691) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g554 ( .A(n_514), .Y(n_554) );
AND2x2_ASAP7_75t_L g620 ( .A(n_514), .B(n_550), .Y(n_620) );
AND2x2_ASAP7_75t_L g631 ( .A(n_514), .B(n_531), .Y(n_631) );
AND2x2_ASAP7_75t_L g640 ( .A(n_514), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_519), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_519), .B(n_581), .Y(n_625) );
INVx2_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g612 ( .A(n_520), .B(n_571), .Y(n_612) );
OR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_531), .Y(n_520) );
INVx2_ASAP7_75t_L g548 ( .A(n_521), .Y(n_548) );
AND2x2_ASAP7_75t_L g639 ( .A(n_521), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g558 ( .A(n_522), .Y(n_558) );
OR2x2_ASAP7_75t_L g656 ( .A(n_522), .B(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_522), .Y(n_719) );
AND2x2_ASAP7_75t_L g559 ( .A(n_531), .B(n_554), .Y(n_559) );
INVx1_ASAP7_75t_L g579 ( .A(n_531), .Y(n_579) );
AND2x2_ASAP7_75t_L g600 ( .A(n_531), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g641 ( .A(n_531), .Y(n_641) );
INVx1_ASAP7_75t_L g657 ( .A(n_531), .Y(n_657) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_531), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B(n_536), .Y(n_533) );
INVxp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_543), .B(n_645), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_543), .A2(n_630), .B1(n_679), .B2(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
OAI211xp5_ASAP7_75t_SL g722 ( .A1(n_544), .A2(n_723), .B(n_725), .C(n_743), .Y(n_722) );
INVx2_ASAP7_75t_L g575 ( .A(n_545), .Y(n_575) );
AND2x2_ASAP7_75t_L g633 ( .A(n_545), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g644 ( .A(n_545), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_546), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
AND2x2_ASAP7_75t_L g617 ( .A(n_547), .B(n_581), .Y(n_617) );
BUFx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g649 ( .A(n_548), .B(n_640), .Y(n_649) );
AND2x2_ASAP7_75t_L g668 ( .A(n_548), .B(n_582), .Y(n_668) );
AND2x4_ASAP7_75t_L g604 ( .A(n_549), .B(n_578), .Y(n_604) );
AND2x2_ASAP7_75t_L g742 ( .A(n_549), .B(n_718), .Y(n_742) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_550), .Y(n_571) );
INVx1_ASAP7_75t_L g582 ( .A(n_550), .Y(n_582) );
INVx1_ASAP7_75t_L g681 ( .A(n_550), .Y(n_681) );
OR2x2_ASAP7_75t_L g572 ( .A(n_554), .B(n_558), .Y(n_572) );
AND2x2_ASAP7_75t_L g581 ( .A(n_554), .B(n_582), .Y(n_581) );
NOR2xp67_ASAP7_75t_L g601 ( .A(n_554), .B(n_602), .Y(n_601) );
OAI221xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_560), .B1(n_570), .B2(n_573), .C(n_577), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g577 ( .A1(n_557), .A2(n_578), .B(n_580), .C(n_583), .Y(n_577) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g602 ( .A(n_558), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_558), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_SL g685 ( .A(n_558), .B(n_579), .Y(n_685) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_558), .Y(n_692) );
AND2x2_ASAP7_75t_L g610 ( .A(n_559), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g647 ( .A(n_559), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_569), .Y(n_560) );
INVx2_ASAP7_75t_L g638 ( .A(n_561), .Y(n_638) );
AOI222xp33_ASAP7_75t_L g687 ( .A1(n_561), .A2(n_571), .B1(n_688), .B2(n_690), .C1(n_691), .C2(n_693), .Y(n_687) );
AND2x2_ASAP7_75t_L g744 ( .A(n_561), .B(n_713), .Y(n_744) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_568), .Y(n_561) );
INVx1_ASAP7_75t_L g634 ( .A(n_562), .Y(n_634) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g586 ( .A(n_567), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g672 ( .A(n_569), .B(n_606), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_570), .A2(n_684), .B(n_686), .Y(n_683) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx2_ASAP7_75t_L g611 ( .A(n_571), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_571), .B(n_578), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_571), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx3_ASAP7_75t_L g637 ( .A(n_575), .Y(n_637) );
OR2x2_ASAP7_75t_L g689 ( .A(n_575), .B(n_611), .Y(n_689) );
AND2x2_ASAP7_75t_L g605 ( .A(n_576), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g643 ( .A(n_576), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_576), .B(n_637), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_576), .B(n_633), .Y(n_659) );
AND2x2_ASAP7_75t_L g663 ( .A(n_576), .B(n_645), .Y(n_663) );
INVxp67_ASAP7_75t_L g595 ( .A(n_578), .Y(n_595) );
BUFx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_580), .A2(n_653), .B1(n_658), .B2(n_659), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_580), .B(n_685), .Y(n_715) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g701 ( .A(n_581), .B(n_692), .Y(n_701) );
AND2x2_ASAP7_75t_L g730 ( .A(n_581), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g735 ( .A(n_581), .B(n_685), .Y(n_735) );
INVx1_ASAP7_75t_L g648 ( .A(n_582), .Y(n_648) );
BUFx2_ASAP7_75t_L g654 ( .A(n_582), .Y(n_654) );
INVx1_ASAP7_75t_L g739 ( .A(n_583), .Y(n_739) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_584), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g615 ( .A(n_585), .Y(n_615) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_586), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g598 ( .A(n_586), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g607 ( .A(n_586), .Y(n_607) );
INVx3_ASAP7_75t_L g645 ( .A(n_586), .Y(n_645) );
OR2x2_ASAP7_75t_L g711 ( .A(n_586), .B(n_712), .Y(n_711) );
AOI211xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_593), .B(n_596), .C(n_608), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_589), .A2(n_726), .B1(n_733), .B2(n_735), .C(n_736), .Y(n_725) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_597), .B(n_603), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_599), .B(n_637), .Y(n_651) );
AND2x2_ASAP7_75t_L g693 ( .A(n_599), .B(n_633), .Y(n_693) );
INVx1_ASAP7_75t_SL g706 ( .A(n_600), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_600), .B(n_654), .Y(n_709) );
INVx1_ASAP7_75t_L g727 ( .A(n_601), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_605), .A2(n_695), .B1(n_697), .B2(n_701), .C(n_702), .Y(n_694) );
AND2x2_ASAP7_75t_L g721 ( .A(n_606), .B(n_713), .Y(n_721) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g705 ( .A(n_607), .Y(n_705) );
AOI21xp33_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_612), .B(n_613), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g676 ( .A(n_611), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g662 ( .A(n_612), .Y(n_662) );
INVx1_ASAP7_75t_L g690 ( .A(n_613), .Y(n_690) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
O2A1O1Ixp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_621), .C(n_624), .Y(n_616) );
OAI31xp33_ASAP7_75t_L g743 ( .A1(n_617), .A2(n_655), .A3(n_742), .B(n_744), .Y(n_743) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g717 ( .A(n_620), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g738 ( .A(n_620), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_622), .B(n_637), .Y(n_665) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g740 ( .A(n_623), .B(n_637), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_632), .B1(n_636), .B2(n_639), .Y(n_627) );
NAND2xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_631), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g667 ( .A(n_631), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g670 ( .A(n_631), .B(n_654), .Y(n_670) );
AND2x2_ASAP7_75t_L g724 ( .A(n_631), .B(n_719), .Y(n_724) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g699 ( .A(n_635), .Y(n_699) );
NOR2xp67_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
OAI32xp33_ASAP7_75t_L g702 ( .A1(n_637), .A2(n_671), .A3(n_703), .B1(n_705), .B2(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g677 ( .A(n_640), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_640), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g700 ( .A(n_644), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B(n_650), .C(n_652), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_648), .B(n_685), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_649), .A2(n_661), .B1(n_662), .B2(n_663), .C(n_664), .Y(n_660) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g661 ( .A(n_659), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_669), .B2(n_671), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND4xp25_ASAP7_75t_SL g726 ( .A(n_669), .B(n_727), .C(n_728), .D(n_729), .Y(n_726) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
NAND4xp25_ASAP7_75t_SL g673 ( .A(n_674), .B(n_687), .C(n_694), .D(n_707), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_678), .B(n_682), .C(n_683), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g704 ( .A(n_680), .Y(n_704) );
INVx2_ASAP7_75t_L g728 ( .A(n_685), .Y(n_728) );
OR2x2_ASAP7_75t_L g737 ( .A(n_692), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B(n_714), .Y(n_707) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g733 ( .A(n_713), .B(n_734), .Y(n_733) );
AOI21xp33_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_716), .B(n_720), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
CKINVDCx16_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_739), .B1(n_740), .B2(n_741), .Y(n_736) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
endmodule