module fake_jpeg_19149_n_137 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_0),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_33),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

AO22x1_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_19),
.B1(n_20),
.B2(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2x1_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_23),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_21),
.B(n_19),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_20),
.B1(n_26),
.B2(n_28),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_33),
.B1(n_35),
.B2(n_16),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_36),
.Y(n_66)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_26),
.B1(n_28),
.B2(n_34),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_58),
.B1(n_67),
.B2(n_41),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_36),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_69),
.C(n_48),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_34),
.B1(n_33),
.B2(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_63),
.Y(n_82)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_16),
.B1(n_15),
.B2(n_27),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_15),
.B(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_22),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_74),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_86),
.B1(n_63),
.B2(n_69),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_27),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_87),
.C(n_88),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_72),
.B1(n_59),
.B2(n_58),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_17),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_70),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_53),
.C(n_29),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_53),
.C(n_25),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_68),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_100),
.Y(n_113)
);

XOR2x2_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_92),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_103),
.B(n_79),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_61),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_78),
.B1(n_85),
.B2(n_77),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_76),
.Y(n_106)
);

OAI321xp33_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_107),
.A3(n_99),
.B1(n_102),
.B2(n_103),
.C(n_95),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_64),
.B1(n_60),
.B2(n_62),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_105),
.B(n_94),
.C(n_83),
.D(n_98),
.Y(n_121)
);

OAI22x1_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_80),
.B1(n_90),
.B2(n_88),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_115),
.B1(n_101),
.B2(n_103),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_104),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_113),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_113),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_104),
.C(n_87),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_118),
.C(n_114),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_107),
.B1(n_106),
.B2(n_96),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_122),
.B1(n_111),
.B2(n_109),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_17),
.B(n_10),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_110),
.C(n_111),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_128),
.B(n_1),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_1),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_127),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_133),
.B(n_134),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_126),
.B(n_123),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_7),
.C(n_5),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_6),
.Y(n_137)
);


endmodule