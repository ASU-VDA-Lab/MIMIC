module fake_jpeg_20780_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_10),
.B(n_4),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_44),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_58),
.B1(n_57),
.B2(n_54),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_18),
.B1(n_26),
.B2(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_55),
.A2(n_45),
.B1(n_18),
.B2(n_25),
.Y(n_80)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_26),
.B1(n_18),
.B2(n_30),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_17),
.B1(n_25),
.B2(n_28),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

NAND2x1p5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_36),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_65),
.B(n_66),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_43),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_36),
.C(n_27),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_20),
.B(n_27),
.C(n_35),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_71),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_38),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_38),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_21),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_88),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_96),
.B1(n_53),
.B2(n_25),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_58),
.B1(n_57),
.B2(n_20),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_39),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_85),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_45),
.B1(n_26),
.B2(n_39),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_86),
.B1(n_28),
.B2(n_57),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_39),
.C(n_31),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_31),
.C(n_30),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_40),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_27),
.B1(n_20),
.B2(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_31),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_54),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_40),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_91),
.B(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_56),
.B(n_22),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_31),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_101),
.A2(n_118),
.B1(n_121),
.B2(n_126),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_63),
.B(n_62),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_72),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_82),
.C(n_70),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_101),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_61),
.A2(n_58),
.B1(n_35),
.B2(n_21),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_22),
.B1(n_30),
.B2(n_24),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_84),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_75),
.B(n_22),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_64),
.A2(n_35),
.B1(n_24),
.B2(n_30),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_79),
.A2(n_35),
.B1(n_24),
.B2(n_33),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_133),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_139),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_140),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_129),
.B(n_85),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_135),
.B(n_149),
.Y(n_174)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_97),
.Y(n_136)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_99),
.B(n_100),
.Y(n_168)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_103),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_153),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_119),
.B1(n_157),
.B2(n_136),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_35),
.B(n_33),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_119),
.A2(n_71),
.B1(n_63),
.B2(n_62),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_91),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_151),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_95),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_106),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_97),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_73),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_155),
.Y(n_186)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_93),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_83),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_33),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_158),
.A2(n_163),
.B1(n_166),
.B2(n_169),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_154),
.B(n_136),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_179),
.B(n_183),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_102),
.B1(n_123),
.B2(n_122),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_123),
.B1(n_117),
.B2(n_122),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_173),
.B1(n_180),
.B2(n_133),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_118),
.B1(n_112),
.B2(n_127),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_172),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_112),
.B1(n_125),
.B2(n_128),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_121),
.B1(n_109),
.B2(n_128),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_128),
.B1(n_113),
.B2(n_115),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_175),
.A2(n_32),
.B1(n_29),
.B2(n_23),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_124),
.A3(n_92),
.B1(n_90),
.B2(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_184),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_104),
.B1(n_120),
.B2(n_76),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_179),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_120),
.B(n_104),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_74),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_74),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_137),
.B(n_76),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_197),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_155),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_212),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_218),
.B1(n_220),
.B2(n_169),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_199),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_143),
.Y(n_201)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_SL g236 ( 
.A(n_202),
.B(n_204),
.C(n_89),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_152),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_208),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_142),
.C(n_138),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_214),
.C(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_211),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_162),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_89),
.C(n_76),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_161),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_32),
.Y(n_240)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_216),
.B(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_159),
.B(n_19),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_176),
.B(n_11),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_187),
.B1(n_160),
.B2(n_186),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_32),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_227),
.C(n_233),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_193),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_202),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_187),
.B1(n_159),
.B2(n_188),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_158),
.B1(n_178),
.B2(n_160),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_192),
.C(n_205),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_228),
.B(n_198),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_183),
.C(n_175),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_196),
.A2(n_89),
.B1(n_32),
.B2(n_29),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_197),
.B1(n_219),
.B2(n_204),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_236),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_29),
.C(n_23),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_193),
.C(n_212),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_211),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_191),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_254),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_256),
.B1(n_261),
.B2(n_263),
.Y(n_271)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_238),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_251),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_250),
.B(n_253),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_196),
.B1(n_216),
.B2(n_191),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_259),
.C(n_241),
.Y(n_270)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_195),
.C(n_217),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_260),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_9),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_210),
.C(n_207),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_225),
.A2(n_195),
.B1(n_200),
.B2(n_29),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_224),
.B(n_8),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_264),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_23),
.B1(n_19),
.B2(n_9),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_0),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_233),
.C(n_231),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_267),
.Y(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_222),
.B(n_231),
.C(n_240),
.D(n_234),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_237),
.C(n_244),
.Y(n_267)
);

XOR2x1_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_236),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_268),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_241),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_12),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_277),
.C(n_252),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_23),
.C(n_19),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_19),
.C(n_9),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_7),
.C(n_14),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_250),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_6),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.C1(n_11),
.C2(n_15),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_264),
.B(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_288),
.Y(n_299)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_291),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_275),
.B(n_282),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_1),
.C(n_2),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_293),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_1),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_2),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_296),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_2),
.C(n_3),
.Y(n_296)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_284),
.A2(n_271),
.B1(n_289),
.B2(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_266),
.B1(n_279),
.B2(n_277),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_278),
.B(n_4),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_306),
.A2(n_292),
.B(n_296),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_298),
.C(n_300),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_314),
.C(n_304),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_3),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_3),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_305),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_3),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

AOI21x1_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_302),
.B(n_297),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_319),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_308),
.B(n_310),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_314),
.B(n_4),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_321),
.C(n_320),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_4),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_5),
.Y(n_327)
);


endmodule