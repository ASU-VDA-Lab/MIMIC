module fake_jpeg_24751_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_2),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_6),
.B(n_1),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_1),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_19),
.Y(n_24)
);

AO22x2_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_17),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_23)
);

AND2x2_ASAP7_75t_SL g18 ( 
.A(n_7),
.B(n_0),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_20),
.B(n_12),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_2),
.C(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_5),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_18),
.B(n_17),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_17),
.C(n_12),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_11),
.B(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_28),
.C(n_11),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_18),
.B(n_17),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_24),
.B1(n_15),
.B2(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.Y(n_33)
);

AOI322xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_5),
.A3(n_10),
.B1(n_22),
.B2(n_26),
.C1(n_28),
.C2(n_27),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_10),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_33),
.C(n_22),
.Y(n_36)
);


endmodule