module fake_jpeg_15074_n_286 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_155;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_18),
.C(n_23),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_62),
.C(n_30),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_27),
.B1(n_21),
.B2(n_29),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_42),
.B1(n_41),
.B2(n_32),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_27),
.B1(n_21),
.B2(n_29),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_27),
.B1(n_16),
.B2(n_29),
.Y(n_68)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_16),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_77),
.B1(n_78),
.B2(n_63),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_73),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_47),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_84),
.Y(n_90)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_42),
.B1(n_41),
.B2(n_37),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_63),
.B1(n_54),
.B2(n_46),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_61),
.B(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_45),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_99),
.B1(n_102),
.B2(n_86),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_62),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_92),
.A2(n_109),
.B(n_25),
.Y(n_134)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_33),
.B1(n_28),
.B2(n_24),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_58),
.B1(n_55),
.B2(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_52),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_72),
.B1(n_85),
.B2(n_70),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_58),
.B1(n_43),
.B2(n_56),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_28),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_64),
.B(n_24),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_37),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_30),
.C(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_64),
.B(n_24),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_45),
.Y(n_109)
);

AOI32xp33_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_53),
.A3(n_83),
.B1(n_77),
.B2(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_121),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_83),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_117),
.C(n_129),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_65),
.B1(n_72),
.B2(n_83),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_91),
.B1(n_108),
.B2(n_111),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_44),
.B(n_70),
.C(n_22),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_134),
.B(n_105),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_122),
.B(n_90),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_65),
.B1(n_82),
.B2(n_81),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_131),
.B1(n_117),
.B2(n_132),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_135),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_87),
.C(n_18),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_80),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_133),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_94),
.A2(n_30),
.B1(n_32),
.B2(n_22),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_91),
.B1(n_109),
.B2(n_89),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_18),
.C(n_71),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_23),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_18),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_91),
.B1(n_97),
.B2(n_101),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_153),
.Y(n_175)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_111),
.B(n_109),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_151),
.B(n_162),
.Y(n_169)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_23),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_152),
.B1(n_119),
.B2(n_115),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_91),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_89),
.B1(n_98),
.B2(n_106),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_154),
.A2(n_156),
.B1(n_112),
.B2(n_32),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_98),
.B1(n_106),
.B2(n_104),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_159),
.B(n_164),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_119),
.A2(n_106),
.B(n_33),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_163),
.Y(n_165)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_167),
.B1(n_185),
.B2(n_187),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_134),
.B1(n_136),
.B2(n_96),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_103),
.C(n_96),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_178),
.C(n_180),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_26),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_177),
.B(n_162),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_112),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_103),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_139),
.A2(n_31),
.B1(n_25),
.B2(n_20),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_185),
.B1(n_187),
.B2(n_176),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_163),
.B1(n_150),
.B2(n_157),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_31),
.B1(n_20),
.B2(n_0),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_141),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_155),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_194),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_146),
.B(n_139),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_147),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_201),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_156),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_197),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_172),
.B1(n_175),
.B2(n_166),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_4),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_164),
.C(n_153),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_207),
.C(n_177),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_140),
.C(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_204),
.Y(n_212)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_1),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_206),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_26),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_217),
.C(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_172),
.B(n_184),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_223),
.B(n_205),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_167),
.C(n_168),
.Y(n_217)
);

OAI22x1_ASAP7_75t_SL g220 ( 
.A1(n_203),
.A2(n_168),
.B1(n_1),
.B2(n_4),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_1),
.C(n_2),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_2),
.C(n_4),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_199),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_226),
.Y(n_227)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_194),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_230),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_216),
.A2(n_209),
.B1(n_204),
.B2(n_207),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_229),
.A2(n_240),
.B1(n_218),
.B2(n_215),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_200),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_220),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_238),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_234),
.A2(n_218),
.B(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_237),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_224),
.B(n_223),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_239),
.A2(n_211),
.B1(n_192),
.B2(n_222),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_236),
.B(n_206),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_249),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_239),
.A2(n_219),
.B(n_191),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_217),
.C(n_213),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_230),
.C(n_228),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_6),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_255),
.C(n_242),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_229),
.C(n_214),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_258),
.B(n_260),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_5),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_262),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_15),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_243),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_265),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_252),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_267),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_249),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_255),
.A2(n_242),
.B1(n_9),
.B2(n_10),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_264),
.A2(n_261),
.B(n_253),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_275),
.B(n_9),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_270),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_13),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_8),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_278),
.B(n_279),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_269),
.B(n_11),
.Y(n_278)
);

FAx1_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_274),
.CI(n_276),
.CON(n_281),
.SN(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_281),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_280),
.B(n_12),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_13),
.B(n_10),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_12),
.Y(n_286)
);


endmodule