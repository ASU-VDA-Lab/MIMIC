module fake_netlist_6_2008_n_573 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_77, n_92, n_42, n_8, n_90, n_24, n_54, n_0, n_87, n_32, n_66, n_85, n_78, n_84, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_95, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_573);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_77;
input n_92;
input n_42;
input n_8;
input n_90;
input n_24;
input n_54;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_78;
input n_84;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_95;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_573;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_111;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_119;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_96;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_109;
wire n_529;
wire n_445;
wire n_425;
wire n_122;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_112;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_107;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_356;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_513;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_570;
wire n_406;
wire n_483;
wire n_102;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_124;
wire n_548;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_523;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_41),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_42),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_8),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_1),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_29),
.Y(n_111)
);

NOR2xp67_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_60),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_46),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_25),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_11),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_11),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_21),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_37),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_33),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_3),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_7),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_32),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_27),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_14),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_57),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_66),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_88),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_31),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_54),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_16),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_62),
.Y(n_149)
);

BUFx2_ASAP7_75t_SL g150 ( 
.A(n_0),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_48),
.B(n_55),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_10),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_91),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_45),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_5),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_4),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_49),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_24),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_17),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_78),
.B(n_77),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_17),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_12),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_92),
.Y(n_165)
);

NOR2xp67_ASAP7_75t_L g166 ( 
.A(n_15),
.B(n_68),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_35),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_53),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_85),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_67),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_20),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_20),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_23),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_86),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_69),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_L g176 ( 
.A(n_38),
.B(n_8),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_79),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_6),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_26),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_52),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_10),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_18),
.Y(n_183)
);

NOR2xp67_ASAP7_75t_L g184 ( 
.A(n_9),
.B(n_19),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_2),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

AND2x4_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_164),
.Y(n_188)
);

BUFx8_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g193 ( 
.A1(n_105),
.A2(n_84),
.B(n_83),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_105),
.B(n_0),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g197 ( 
.A(n_105),
.B(n_64),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

AND2x4_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_110),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_103),
.B(n_6),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_9),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_103),
.A2(n_34),
.B(n_58),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_102),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_12),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_110),
.A2(n_13),
.B1(n_15),
.B2(n_19),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_100),
.B(n_116),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_97),
.A2(n_13),
.B1(n_40),
.B2(n_51),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_61),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_158),
.B(n_174),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_120),
.B(n_123),
.Y(n_222)
);

CKINVDCx6p67_ASAP7_75t_R g223 ( 
.A(n_143),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_118),
.Y(n_224)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_158),
.B(n_174),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_111),
.B(n_98),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_169),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_121),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_151),
.B(n_180),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_124),
.B(n_185),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_134),
.B(n_183),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_99),
.B(n_167),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g235 ( 
.A(n_161),
.B(n_145),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_108),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_114),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_117),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_147),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_125),
.B(n_144),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_127),
.B(n_129),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_128),
.A2(n_132),
.B(n_181),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_155),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_156),
.B(n_162),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g245 ( 
.A(n_126),
.B(n_135),
.C(n_183),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_152),
.A2(n_126),
.B1(n_135),
.B2(n_178),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_172),
.Y(n_247)
);

INVxp33_ASAP7_75t_SL g248 ( 
.A(n_150),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_104),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_152),
.A2(n_184),
.B1(n_166),
.B2(n_176),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_104),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_133),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_119),
.A2(n_142),
.B1(n_149),
.B2(n_177),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_137),
.B(n_179),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_138),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_157),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_159),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_119),
.A2(n_142),
.B1(n_149),
.B2(n_170),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_106),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_173),
.B(n_175),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_96),
.Y(n_261)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_199),
.B(n_112),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_168),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_223),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g265 ( 
.A(n_199),
.B(n_208),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_222),
.B(n_250),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_225),
.A2(n_106),
.B1(n_177),
.B2(n_170),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_165),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_198),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_195),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_225),
.A2(n_141),
.B1(n_131),
.B2(n_130),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_190),
.Y(n_274)
);

AO22x2_ASAP7_75t_L g275 ( 
.A1(n_215),
.A2(n_141),
.B1(n_131),
.B2(n_130),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_251),
.Y(n_276)
);

AND2x6_ASAP7_75t_L g277 ( 
.A(n_208),
.B(n_113),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_115),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_230),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_190),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_222),
.B(n_196),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_235),
.A2(n_136),
.B1(n_146),
.B2(n_153),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_190),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_258),
.B(n_248),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_192),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_201),
.A2(n_253),
.B1(n_246),
.B2(n_215),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_216),
.B(n_259),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_192),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_202),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_205),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_188),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_205),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_209),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_204),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_206),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_235),
.A2(n_186),
.B1(n_220),
.B2(n_210),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_211),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_203),
.B(n_219),
.Y(n_298)
);

BUFx8_ASAP7_75t_SL g299 ( 
.A(n_232),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_209),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_187),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_187),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_196),
.B(n_228),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_207),
.B(n_214),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_220),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_207),
.B(n_214),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_233),
.B(n_260),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_245),
.B(n_186),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_240),
.B(n_242),
.Y(n_309)
);

OR2x6_ASAP7_75t_L g310 ( 
.A(n_201),
.B(n_245),
.Y(n_310)
);

NAND2xp33_ASAP7_75t_L g311 ( 
.A(n_235),
.B(n_230),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_227),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_227),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_256),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_257),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_213),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_235),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_269),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_265),
.B(n_240),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_265),
.B(n_287),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_282),
.B(n_218),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_188),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_316),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_270),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

NOR3x1_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_258),
.C(n_244),
.Y(n_331)
);

NOR2x2_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_253),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_304),
.A2(n_241),
.B1(n_254),
.B2(n_221),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_264),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_R g335 ( 
.A(n_264),
.B(n_189),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_261),
.B(n_252),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_262),
.B(n_234),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_262),
.B(n_291),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_281),
.B(n_218),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_191),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_234),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_263),
.B(n_254),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_234),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_281),
.B(n_306),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_303),
.A2(n_221),
.B1(n_238),
.B2(n_237),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_283),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_268),
.B(n_194),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_283),
.Y(n_349)
);

A2O1A1Ixp33_ASAP7_75t_L g350 ( 
.A1(n_303),
.A2(n_244),
.B(n_193),
.C(n_308),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_271),
.B(n_243),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_231),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_280),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_299),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_266),
.B(n_237),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_299),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_266),
.A2(n_217),
.B1(n_246),
.B2(n_197),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_276),
.B(n_243),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_277),
.A2(n_309),
.B1(n_267),
.B2(n_273),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_285),
.Y(n_360)
);

NAND2x1p5_ASAP7_75t_L g361 ( 
.A(n_272),
.B(n_212),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_289),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_277),
.B(n_238),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_277),
.B(n_236),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_284),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_294),
.B(n_224),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_365),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_296),
.Y(n_368)
);

CKINVDCx8_ASAP7_75t_R g369 ( 
.A(n_354),
.Y(n_369)
);

OAI21xp33_ASAP7_75t_L g370 ( 
.A1(n_327),
.A2(n_310),
.B(n_275),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_L g371 ( 
.A1(n_357),
.A2(n_310),
.B1(n_312),
.B2(n_247),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_344),
.A2(n_311),
.B(n_272),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_342),
.A2(n_311),
.B(n_297),
.C(n_295),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_341),
.A2(n_343),
.B(n_322),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_319),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_320),
.Y(n_376)
);

O2A1O1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_326),
.A2(n_229),
.B(n_310),
.C(n_239),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_336),
.B(n_305),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_323),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_329),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_350),
.A2(n_302),
.B(n_301),
.C(n_239),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_305),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_329),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_328),
.B(n_292),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_333),
.B(n_279),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_334),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_340),
.B(n_362),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_366),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_318),
.A2(n_275),
.B1(n_286),
.B2(n_314),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_338),
.A2(n_275),
.B1(n_290),
.B2(n_293),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_321),
.B(n_362),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

AOI21x1_ASAP7_75t_L g397 ( 
.A1(n_337),
.A2(n_290),
.B(n_288),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_332),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_332),
.A2(n_280),
.B1(n_293),
.B2(n_300),
.Y(n_399)
);

A2O1A1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_350),
.A2(n_313),
.B(n_300),
.C(n_288),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_313),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

A2O1A1Ixp33_ASAP7_75t_L g403 ( 
.A1(n_346),
.A2(n_313),
.B(n_363),
.C(n_364),
.Y(n_403)
);

OR2x6_ASAP7_75t_L g404 ( 
.A(n_324),
.B(n_356),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_324),
.B(n_335),
.Y(n_405)
);

BUFx8_ASAP7_75t_SL g406 ( 
.A(n_354),
.Y(n_406)
);

NAND3xp33_ASAP7_75t_L g407 ( 
.A(n_345),
.B(n_349),
.C(n_347),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_324),
.A2(n_360),
.B1(n_325),
.B2(n_361),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_327),
.B(n_278),
.C(n_307),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_344),
.A2(n_343),
.B(n_341),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_326),
.A2(n_342),
.B1(n_327),
.B2(n_344),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_320),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_327),
.B(n_359),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_344),
.A2(n_343),
.B(n_341),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_326),
.A2(n_342),
.B1(n_327),
.B2(n_344),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_327),
.B(n_291),
.Y(n_416)
);

O2A1O1Ixp5_ASAP7_75t_L g417 ( 
.A1(n_344),
.A2(n_326),
.B(n_339),
.C(n_306),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_342),
.A2(n_327),
.B(n_326),
.C(n_355),
.Y(n_418)
);

A2O1A1Ixp33_ASAP7_75t_SL g419 ( 
.A1(n_355),
.A2(n_342),
.B(n_327),
.C(n_348),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_353),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_326),
.A2(n_342),
.B1(n_344),
.B2(n_306),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_365),
.Y(n_422)
);

O2A1O1Ixp33_ASAP7_75t_L g423 ( 
.A1(n_344),
.A2(n_326),
.B(n_304),
.C(n_306),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_344),
.A2(n_343),
.B(n_341),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_319),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_SL g426 ( 
.A(n_405),
.B(n_389),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_389),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_367),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_413),
.A2(n_409),
.B1(n_421),
.B2(n_411),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_368),
.B(n_422),
.Y(n_430)
);

OAI221xp5_ASAP7_75t_L g431 ( 
.A1(n_415),
.A2(n_370),
.B1(n_391),
.B2(n_386),
.C(n_396),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_392),
.Y(n_432)
);

A2O1A1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_423),
.A2(n_417),
.B(n_377),
.C(n_424),
.Y(n_433)
);

AO31x2_ASAP7_75t_L g434 ( 
.A1(n_381),
.A2(n_400),
.A3(n_373),
.B(n_403),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_383),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_376),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_390),
.B(n_388),
.Y(n_437)
);

BUFx2_ASAP7_75t_SL g438 ( 
.A(n_387),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_385),
.A2(n_408),
.B1(n_372),
.B2(n_395),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_393),
.Y(n_440)
);

AO31x2_ASAP7_75t_L g441 ( 
.A1(n_394),
.A2(n_374),
.A3(n_424),
.B(n_410),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_378),
.B(n_382),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_398),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_406),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_420),
.Y(n_445)
);

AOI221xp5_ASAP7_75t_L g446 ( 
.A1(n_371),
.A2(n_399),
.B1(n_375),
.B2(n_379),
.C(n_425),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_412),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

INVx6_ASAP7_75t_L g449 ( 
.A(n_404),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_414),
.A2(n_402),
.B1(n_384),
.B2(n_420),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_401),
.B(n_384),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_404),
.B(n_407),
.Y(n_452)
);

AO31x2_ASAP7_75t_L g453 ( 
.A1(n_397),
.A2(n_381),
.A3(n_350),
.B(n_400),
.Y(n_453)
);

OAI22xp33_ASAP7_75t_L g454 ( 
.A1(n_369),
.A2(n_415),
.B1(n_411),
.B2(n_357),
.Y(n_454)
);

AO31x2_ASAP7_75t_L g455 ( 
.A1(n_381),
.A2(n_350),
.A3(n_400),
.B(n_418),
.Y(n_455)
);

O2A1O1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_418),
.A2(n_326),
.B(n_419),
.C(n_413),
.Y(n_456)
);

AO31x2_ASAP7_75t_L g457 ( 
.A1(n_381),
.A2(n_350),
.A3(n_400),
.B(n_418),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_411),
.B(n_342),
.Y(n_458)
);

INVx8_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

O2A1O1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_418),
.A2(n_326),
.B(n_419),
.C(n_413),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_367),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_413),
.A2(n_411),
.B1(n_415),
.B2(n_409),
.Y(n_462)
);

OAI22x1_ASAP7_75t_L g463 ( 
.A1(n_398),
.A2(n_357),
.B1(n_365),
.B2(n_393),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_411),
.B(n_342),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_392),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_380),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_387),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_411),
.B(n_342),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_413),
.A2(n_411),
.B1(n_415),
.B2(n_409),
.Y(n_471)
);

AO32x2_ASAP7_75t_L g472 ( 
.A1(n_391),
.A2(n_394),
.A3(n_399),
.B1(n_286),
.B2(n_201),
.Y(n_472)
);

A2O1A1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_423),
.A2(n_415),
.B(n_411),
.C(n_418),
.Y(n_473)
);

AO21x1_ASAP7_75t_L g474 ( 
.A1(n_413),
.A2(n_326),
.B(n_377),
.Y(n_474)
);

AO32x2_ASAP7_75t_L g475 ( 
.A1(n_391),
.A2(n_394),
.A3(n_399),
.B1(n_286),
.B2(n_201),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_392),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_411),
.B(n_342),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_411),
.B(n_342),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_464),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_477),
.Y(n_480)
);

AO31x2_ASAP7_75t_L g481 ( 
.A1(n_433),
.A2(n_473),
.A3(n_474),
.B(n_439),
.Y(n_481)
);

NAND2x1_ASAP7_75t_L g482 ( 
.A(n_427),
.B(n_445),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_469),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_478),
.A2(n_429),
.B1(n_471),
.B2(n_462),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_427),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_435),
.Y(n_487)
);

OAI21xp33_ASAP7_75t_SL g488 ( 
.A1(n_446),
.A2(n_450),
.B(n_442),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_436),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_456),
.A2(n_460),
.B(n_451),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_454),
.A2(n_431),
.B1(n_445),
.B2(n_430),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_SL g492 ( 
.A1(n_428),
.A2(n_437),
.B1(n_467),
.B2(n_459),
.Y(n_492)
);

AND3x2_ASAP7_75t_L g493 ( 
.A(n_448),
.B(n_452),
.C(n_437),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_468),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_449),
.A2(n_468),
.B1(n_447),
.B2(n_476),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_463),
.A2(n_452),
.B1(n_440),
.B2(n_467),
.Y(n_496)
);

NAND3xp33_ASAP7_75t_L g497 ( 
.A(n_432),
.B(n_466),
.C(n_467),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_443),
.B(n_449),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_441),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g500 ( 
.A1(n_455),
.A2(n_457),
.B(n_441),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_426),
.A2(n_459),
.B1(n_475),
.B2(n_472),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_465),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_444),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_434),
.B(n_453),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_438),
.B(n_472),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_475),
.A2(n_458),
.B1(n_470),
.B2(n_464),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_484),
.A2(n_490),
.B(n_491),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_499),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_506),
.B(n_479),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_485),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_504),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_479),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_501),
.A2(n_480),
.B1(n_505),
.B2(n_500),
.Y(n_513)
);

AO21x2_ASAP7_75t_L g514 ( 
.A1(n_487),
.A2(n_489),
.B(n_494),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_486),
.B(n_493),
.Y(n_515)
);

OA21x2_ASAP7_75t_L g516 ( 
.A1(n_481),
.A2(n_496),
.B(n_488),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_486),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_481),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_481),
.B(n_485),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_495),
.A2(n_497),
.B(n_498),
.Y(n_520)
);

OAI31xp33_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_498),
.A3(n_502),
.B(n_483),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_492),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_519),
.B(n_483),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_510),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_508),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_482),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_512),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_512),
.B(n_502),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_510),
.B(n_503),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_503),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_515),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_512),
.A2(n_513),
.B(n_507),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_516),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_508),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_519),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_533),
.B(n_518),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_533),
.B(n_518),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_527),
.B(n_528),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_527),
.B(n_518),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_525),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_R g541 ( 
.A(n_529),
.B(n_520),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_535),
.B(n_518),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_524),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_521),
.B(n_511),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_535),
.B(n_526),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_525),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_545),
.B(n_537),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_540),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_545),
.B(n_537),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_543),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_538),
.B(n_523),
.Y(n_551)
);

CKINVDCx8_ASAP7_75t_R g552 ( 
.A(n_541),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_550),
.B(n_539),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_552),
.B(n_521),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_552),
.B(n_530),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_547),
.B(n_536),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_547),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_549),
.B(n_542),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_557),
.Y(n_559)
);

OAI322xp33_ASAP7_75t_L g560 ( 
.A1(n_554),
.A2(n_548),
.A3(n_519),
.B1(n_530),
.B2(n_522),
.C1(n_544),
.C2(n_540),
.Y(n_560)
);

AOI21xp33_ASAP7_75t_L g561 ( 
.A1(n_555),
.A2(n_544),
.B(n_520),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_555),
.A2(n_531),
.B1(n_522),
.B2(n_520),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_559),
.B(n_558),
.Y(n_563)
);

AOI211xp5_ASAP7_75t_SL g564 ( 
.A1(n_563),
.A2(n_560),
.B(n_561),
.C(n_559),
.Y(n_564)
);

NOR3xp33_ASAP7_75t_L g565 ( 
.A(n_564),
.B(n_553),
.C(n_532),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_565),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_566),
.Y(n_567)
);

AOI22x1_ASAP7_75t_L g568 ( 
.A1(n_567),
.A2(n_515),
.B1(n_558),
.B2(n_556),
.Y(n_568)
);

AOI22x1_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_515),
.B1(n_517),
.B2(n_549),
.Y(n_569)
);

AOI222xp33_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_562),
.B1(n_532),
.B2(n_513),
.C1(n_515),
.C2(n_551),
.Y(n_570)
);

AOI222xp33_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_515),
.B1(n_513),
.B2(n_531),
.C1(n_546),
.C2(n_534),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_571),
.B(n_515),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_520),
.B1(n_515),
.B2(n_514),
.Y(n_573)
);


endmodule