module real_jpeg_1051_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_0),
.A2(n_31),
.B1(n_37),
.B2(n_83),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_0),
.A2(n_58),
.B1(n_59),
.B2(n_83),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_0),
.A2(n_74),
.B1(n_76),
.B2(n_83),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_2),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_3),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_3),
.A2(n_26),
.B1(n_31),
.B2(n_37),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_3),
.A2(n_26),
.B1(n_74),
.B2(n_76),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_4),
.A2(n_31),
.B1(n_37),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_66),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_66),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_4),
.A2(n_66),
.B1(n_74),
.B2(n_76),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_7),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_7),
.A2(n_31),
.B1(n_37),
.B2(n_135),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_135),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_7),
.A2(n_74),
.B1(n_76),
.B2(n_135),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_31),
.B1(n_37),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_8),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_63),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_8),
.A2(n_63),
.B1(n_74),
.B2(n_76),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_9),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_9),
.A2(n_31),
.B1(n_37),
.B2(n_175),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_175),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_9),
.A2(n_74),
.B1(n_76),
.B2(n_175),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_10),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_10),
.A2(n_31),
.B1(n_37),
.B2(n_113),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_113),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_10),
.A2(n_74),
.B1(n_76),
.B2(n_113),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_14),
.B(n_28),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_14),
.B(n_41),
.Y(n_212)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_14),
.A2(n_16),
.B(n_37),
.C(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_14),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_14),
.B(n_57),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_14),
.A2(n_31),
.B1(n_37),
.B2(n_225),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_14),
.B(n_71),
.C(n_74),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_225),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_14),
.B(n_103),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_14),
.B(n_92),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_15),
.Y(n_342)
);

BUFx12_ASAP7_75t_L g344 ( 
.A(n_15),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_16),
.A2(n_37),
.B(n_56),
.C(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_16),
.B(n_37),
.Y(n_56)
);

AO22x2_ASAP7_75t_L g57 ( 
.A1(n_16),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_57)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_17),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_17),
.A2(n_40),
.B1(n_74),
.B2(n_76),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_17),
.A2(n_31),
.B1(n_37),
.B2(n_40),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_342),
.B(n_343),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_45),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_42),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_23),
.B(n_341),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_24),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_24),
.B(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_39),
.B2(n_41),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_25),
.A2(n_29),
.B1(n_41),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_38)
);

AOI32xp33_ASAP7_75t_L g195 ( 
.A1(n_27),
.A2(n_34),
.A3(n_37),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_27),
.A2(n_84),
.B(n_225),
.C(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_39),
.B(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_29),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_29),
.A2(n_41),
.B1(n_134),
.B2(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_38),
.Y(n_29)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_30),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_30),
.A2(n_82),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_30),
.B(n_112),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_30),
.A2(n_84),
.B1(n_85),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_30),
.A2(n_110),
.B(n_189),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_30)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_31),
.B(n_35),
.Y(n_197)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OAI21x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_337),
.B(n_339),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_325),
.B(n_336),
.Y(n_46)
);

AO21x1_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_151),
.B(n_322),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_138),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_114),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_50),
.B(n_114),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_95),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_79),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_52),
.A2(n_53),
.B(n_67),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_52),
.B(n_79),
.C(n_95),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_67),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_64),
.B1(n_65),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_54),
.A2(n_62),
.B1(n_64),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_54),
.A2(n_64),
.B1(n_89),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_54),
.A2(n_191),
.B(n_193),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_54),
.A2(n_193),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_55),
.B(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_55),
.A2(n_57),
.B1(n_192),
.B2(n_209),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_55),
.A2(n_57),
.B(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_57),
.B(n_172),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_59),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_58),
.A2(n_61),
.B(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_59),
.B(n_270),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_64),
.A2(n_131),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_64),
.A2(n_171),
.B(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_73),
.B1(n_77),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_68),
.A2(n_73),
.B1(n_218),
.B2(n_252),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_68),
.A2(n_220),
.B(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_92),
.B1(n_108),
.B2(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_69),
.A2(n_92),
.B1(n_129),
.B2(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_69),
.A2(n_217),
.B(n_219),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_69),
.B(n_221),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_73),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_73),
.A2(n_241),
.B(n_252),
.Y(n_251)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_74),
.B(n_281),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_94),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_80),
.A2(n_81),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g149 ( 
.A(n_81),
.B(n_87),
.C(n_91),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_81),
.B(n_142),
.C(n_149),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_84),
.A2(n_133),
.B(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_90),
.A2(n_91),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_91),
.B(n_143),
.C(n_147),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_92),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_99),
.B(n_109),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_97),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_106),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_99),
.B1(n_109),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_98),
.A2(n_99),
.B1(n_106),
.B2(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_103),
.B(n_104),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_100),
.A2(n_103),
.B1(n_126),
.B2(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_100),
.A2(n_225),
.B(n_258),
.Y(n_282)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_101),
.A2(n_102),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_101),
.A2(n_102),
.B1(n_200),
.B2(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_101),
.B(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_101),
.A2(n_256),
.B(n_257),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_101),
.A2(n_102),
.B1(n_256),
.B2(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_102),
.A2(n_215),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_102),
.B(n_229),
.Y(n_258)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_103),
.A2(n_228),
.B(n_285),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_106),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.C(n_121),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_130),
.C(n_132),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_123),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_132),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_137),
.B(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_138),
.A2(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_150),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_139),
.B(n_150),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_144),
.Y(n_331)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_148),
.Y(n_329)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_176),
.B(n_321),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_153),
.B(n_156),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_162),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_169),
.C(n_173),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_164),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_165),
.B(n_167),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_166),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_168),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_202),
.B(n_320),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_178),
.B(n_180),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.C(n_187),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_181),
.B(n_185),
.Y(n_305)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_187),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_194),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_188),
.B(n_190),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_194),
.B(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_195),
.A2(n_198),
.B1(n_199),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI31xp33_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_302),
.A3(n_312),
.B(n_317),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_246),
.B(n_301),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_230),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_205),
.B(n_230),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_216),
.C(n_222),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_206),
.B(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_211),
.C(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_216),
.B(n_222),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_226),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_242),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_231),
.B(n_243),
.C(n_245),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_232),
.B(n_237),
.C(n_238),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_296),
.B(n_300),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_265),
.B(n_295),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_259),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_259),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.C(n_254),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_255),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_263),
.C(n_264),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_277),
.B(n_294),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_273),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_273),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_292),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_288),
.B(n_293),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_283),
.B(n_287),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_286),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_291),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_299),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI21xp33_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_306),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.C(n_310),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_316),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_335),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_335),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_334),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_330),
.B1(n_332),
.B2(n_333),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_328),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_330),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_332),
.C(n_334),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_338),
.Y(n_341)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);


endmodule