module fake_jpeg_22403_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_0),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_26),
.B1(n_22),
.B2(n_19),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_36),
.B1(n_39),
.B2(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_15),
.B1(n_18),
.B2(n_22),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_16),
.B1(n_29),
.B2(n_28),
.Y(n_74)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_32),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_60),
.B(n_34),
.Y(n_95)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_63),
.Y(n_83)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_37),
.B1(n_33),
.B2(n_32),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_59),
.B1(n_61),
.B2(n_64),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_57),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_37),
.B1(n_33),
.B2(n_36),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_33),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_36),
.B1(n_15),
.B2(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_69),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_23),
.B1(n_17),
.B2(n_20),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_19),
.B1(n_38),
.B2(n_39),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_45),
.B(n_21),
.C(n_34),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_30),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_16),
.B1(n_29),
.B2(n_28),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_84)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_24),
.B1(n_23),
.B2(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_92),
.B1(n_99),
.B2(n_102),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_85),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_37),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_52),
.B1(n_37),
.B2(n_24),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_37),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_95),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_37),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_101),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_34),
.C(n_42),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_97),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_34),
.C(n_42),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_35),
.B1(n_50),
.B2(n_21),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_73),
.B1(n_55),
.B2(n_63),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_27),
.B1(n_20),
.B2(n_35),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_106),
.Y(n_141)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_71),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_110),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_70),
.B1(n_69),
.B2(n_71),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_54),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_111),
.B(n_114),
.Y(n_148)
);

INVx2_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_30),
.B1(n_25),
.B2(n_3),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_74),
.A3(n_70),
.B1(n_60),
.B2(n_67),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_90),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_115),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_121),
.B(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_59),
.B(n_77),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_59),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_87),
.A2(n_59),
.B1(n_66),
.B2(n_68),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_125),
.B1(n_98),
.B2(n_92),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_81),
.A2(n_79),
.B1(n_30),
.B2(n_25),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_126),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_140),
.B1(n_126),
.B2(n_112),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_93),
.Y(n_132)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_143),
.B1(n_4),
.B2(n_6),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_122),
.C(n_120),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_144),
.C(n_145),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_120),
.B(n_124),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_30),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_116),
.A2(n_30),
.B1(n_25),
.B2(n_14),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_14),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_1),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_2),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_154),
.B(n_166),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_125),
.C(n_121),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_160),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_117),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_170),
.B1(n_143),
.B2(n_139),
.Y(n_183)
);

INVxp33_ASAP7_75t_SL g163 ( 
.A(n_147),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_163),
.Y(n_175)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_168),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_106),
.C(n_5),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_145),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_171),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_131),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_158),
.A2(n_149),
.B1(n_146),
.B2(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_165),
.A2(n_146),
.B1(n_129),
.B2(n_128),
.Y(n_173)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_167),
.B(n_142),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_180),
.C(n_157),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_183),
.B1(n_168),
.B2(n_127),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_138),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_185),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_166),
.A2(n_139),
.B(n_142),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_173),
.B1(n_181),
.B2(n_172),
.Y(n_201)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_169),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_159),
.C(n_157),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_194),
.C(n_196),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_184),
.B(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_161),
.C(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_155),
.C(n_127),
.Y(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_144),
.C(n_150),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_205),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_152),
.C(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_170),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_207),
.Y(n_210)
);

AO221x1_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_182),
.B1(n_188),
.B2(n_191),
.C(n_197),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_211),
.B(n_212),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_195),
.CI(n_192),
.CON(n_212),
.SN(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_205),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_215),
.B(n_216),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_214),
.B(n_183),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_198),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_200),
.A3(n_208),
.B1(n_213),
.B2(n_9),
.C1(n_10),
.C2(n_4),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_198),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_206),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_218),
.A2(n_210),
.B(n_134),
.C(n_216),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_223),
.B(n_12),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_12),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_12),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_225),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_7),
.C(n_8),
.Y(n_228)
);

OAI21x1_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_7),
.B(n_8),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_227),
.C(n_9),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_11),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_11),
.Y(n_232)
);


endmodule