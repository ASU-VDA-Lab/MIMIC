module fake_jpeg_15381_n_350 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_350);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_350;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_44),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_43),
.B1(n_26),
.B2(n_28),
.Y(n_56)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_34),
.B1(n_24),
.B2(n_33),
.Y(n_58)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_27),
.B1(n_24),
.B2(n_30),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_52),
.A2(n_55),
.B1(n_18),
.B2(n_32),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_27),
.B1(n_24),
.B2(n_30),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_43),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_32),
.B1(n_34),
.B2(n_26),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_69),
.B1(n_28),
.B2(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_32),
.B1(n_34),
.B2(n_26),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_75),
.A2(n_110),
.B1(n_21),
.B2(n_20),
.Y(n_134)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_77),
.A2(n_23),
.B1(n_17),
.B2(n_31),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_83),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_79),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_44),
.B(n_49),
.C(n_38),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g133 ( 
.A1(n_80),
.A2(n_20),
.B(n_17),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_19),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_38),
.B(n_43),
.C(n_39),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_84),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_38),
.B(n_43),
.C(n_32),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_89),
.Y(n_124)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_93),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_32),
.B(n_25),
.C(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_67),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_96),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_25),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_106),
.B1(n_21),
.B2(n_29),
.Y(n_130)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_29),
.B1(n_21),
.B2(n_42),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_54),
.A2(n_21),
.B1(n_29),
.B2(n_17),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_20),
.B(n_48),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_68),
.C(n_20),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_127),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_84),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_81),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_122),
.B(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_48),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_48),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_136),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_130),
.B(n_132),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_87),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_134),
.B(n_85),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_79),
.A2(n_46),
.B1(n_29),
.B2(n_20),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_135),
.A2(n_142),
.B1(n_93),
.B2(n_90),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_75),
.B(n_48),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_77),
.A2(n_46),
.B1(n_36),
.B2(n_19),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_108),
.B1(n_103),
.B2(n_90),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_112),
.C(n_100),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_147),
.B(n_154),
.Y(n_195)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_117),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_156),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_150),
.A2(n_153),
.B1(n_160),
.B2(n_131),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_75),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_171),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_86),
.B(n_76),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_157),
.A2(n_159),
.B(n_139),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_165),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_89),
.B(n_91),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_107),
.B1(n_101),
.B2(n_91),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_161),
.A2(n_163),
.B1(n_167),
.B2(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_113),
.B(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_100),
.B1(n_98),
.B2(n_94),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_113),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_104),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_170),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_92),
.B1(n_106),
.B2(n_109),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_120),
.A2(n_105),
.B1(n_111),
.B2(n_13),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_119),
.A2(n_36),
.A3(n_31),
.B1(n_23),
.B2(n_19),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_143),
.C(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_144),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_97),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_155),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_177),
.B(n_183),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_143),
.B(n_124),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_23),
.C(n_36),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_134),
.B1(n_130),
.B2(n_124),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_205),
.B1(n_174),
.B2(n_167),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_117),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_198),
.C(n_207),
.Y(n_221)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_196),
.A2(n_208),
.B1(n_31),
.B2(n_2),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_201),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_139),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_152),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_206),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_132),
.B(n_128),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_204),
.B(n_161),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_173),
.A2(n_118),
.B1(n_141),
.B2(n_122),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_158),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_115),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_173),
.A2(n_141),
.B1(n_116),
.B2(n_137),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_171),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_182),
.B(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_213),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_145),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_223),
.C(n_226),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_231),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_184),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_233),
.B1(n_187),
.B2(n_179),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_157),
.C(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_164),
.C(n_149),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_227),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_228),
.A2(n_234),
.B(n_189),
.Y(n_259)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_156),
.Y(n_232)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_160),
.B1(n_137),
.B2(n_97),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_19),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_208),
.C(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_203),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_239),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_195),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_237),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_179),
.B(n_1),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_217),
.A2(n_194),
.B1(n_209),
.B2(n_196),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_240),
.A2(n_263),
.B(n_1),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_199),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_245),
.C(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_199),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_192),
.C(n_204),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_218),
.C(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_214),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_9),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_193),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_259),
.A2(n_241),
.B(n_258),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_226),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_235),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_229),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_180),
.B(n_178),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_269),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_236),
.B1(n_231),
.B2(n_213),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_270),
.B1(n_271),
.B2(n_244),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_267),
.B(n_284),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_220),
.B1(n_225),
.B2(n_212),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_215),
.B1(n_212),
.B2(n_230),
.Y(n_271)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_263),
.B(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_257),
.A2(n_233),
.B(n_215),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_255),
.B1(n_260),
.B2(n_245),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_257),
.A2(n_239),
.B(n_180),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_178),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_279),
.C(n_242),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_242),
.B(n_190),
.C(n_2),
.Y(n_279)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_9),
.Y(n_285)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_7),
.C(n_10),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_243),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_297),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_267),
.B(n_248),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_265),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_278),
.A2(n_264),
.B1(n_256),
.B2(n_255),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_270),
.B1(n_268),
.B2(n_6),
.Y(n_307)
);

AOI221xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_274),
.B1(n_276),
.B2(n_273),
.C(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_295),
.B(n_302),
.Y(n_317)
);

AO22x1_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_250),
.B1(n_264),
.B2(n_249),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_303),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_10),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_266),
.B(n_277),
.CI(n_269),
.CON(n_303),
.SN(n_303)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_304),
.B(n_310),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_268),
.C(n_279),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_309),
.C(n_313),
.Y(n_327)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_307),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_R g308 ( 
.A(n_290),
.B(n_10),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_308),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_3),
.C(n_5),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_11),
.B1(n_14),
.B2(n_7),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_314),
.B(n_315),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_13),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_303),
.C(n_286),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_318),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_290),
.C(n_293),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_312),
.A2(n_299),
.B1(n_311),
.B2(n_305),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_318),
.B1(n_301),
.B2(n_306),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_15),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_311),
.A2(n_298),
.B(n_297),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_6),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_287),
.Y(n_328)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_294),
.Y(n_329)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_329),
.Y(n_336)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_330),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_13),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_332),
.Y(n_341)
);

XNOR2x1_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_5),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_333),
.A2(n_337),
.B1(n_323),
.B2(n_321),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_15),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_322),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_339),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_326),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_320),
.B(n_335),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_343),
.A2(n_345),
.B(n_340),
.Y(n_346)
);

NOR3xp33_ASAP7_75t_SL g345 ( 
.A(n_338),
.B(n_333),
.C(n_327),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_344),
.Y(n_347)
);

BUFx24_ASAP7_75t_SL g348 ( 
.A(n_347),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_337),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_341),
.Y(n_350)
);


endmodule