module fake_jpeg_12529_n_471 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_471);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_471;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_60),
.B(n_61),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_24),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_43),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_65),
.B(n_73),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_66),
.B(n_91),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_27),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_67),
.B(n_72),
.Y(n_144)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_50),
.Y(n_68)
);

INVx5_ASAP7_75t_SL g161 ( 
.A(n_68),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_27),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_0),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_79),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_82),
.B(n_85),
.Y(n_158)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_49),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_40),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_86),
.B(n_89),
.Y(n_159)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_17),
.B(n_14),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_17),
.B(n_14),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_92),
.B(n_94),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_40),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_12),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_96),
.B(n_108),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_99),
.B(n_102),
.Y(n_171)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_48),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_30),
.B(n_44),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_41),
.Y(n_151)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_107),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_38),
.Y(n_108)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_30),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_112),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_38),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_34),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_35),
.B(n_12),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_30),
.B1(n_31),
.B2(n_20),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_122),
.A2(n_127),
.B1(n_131),
.B2(n_136),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_53),
.B1(n_20),
.B2(n_39),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_37),
.B1(n_33),
.B2(n_47),
.Y(n_131)
);

BUFx2_ASAP7_75t_SL g132 ( 
.A(n_109),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_132),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_37),
.B1(n_57),
.B2(n_35),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_133),
.A2(n_167),
.B1(n_183),
.B2(n_107),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_64),
.B(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_156),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_69),
.A2(n_65),
.B1(n_84),
.B2(n_103),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_139),
.A2(n_151),
.B(n_9),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_69),
.A2(n_53),
.B1(n_41),
.B2(n_51),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_140),
.A2(n_172),
.B1(n_176),
.B2(n_181),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_70),
.B(n_56),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_157),
.B(n_162),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_75),
.B(n_114),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_110),
.A2(n_62),
.B1(n_80),
.B2(n_78),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_81),
.A2(n_57),
.B1(n_56),
.B2(n_46),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_83),
.B(n_98),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_180),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_65),
.A2(n_53),
.B1(n_51),
.B2(n_47),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_58),
.B(n_55),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_63),
.A2(n_46),
.B1(n_44),
.B2(n_3),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_116),
.A2(n_44),
.B1(n_2),
.B2(n_5),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_105),
.A2(n_0),
.B1(n_2),
.B2(n_6),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_79),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_SL g186 ( 
.A(n_112),
.Y(n_186)
);

BUFx24_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

NAND2x1_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_105),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_189),
.B(n_220),
.C(n_216),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_192),
.Y(n_276)
);

INVx3_ASAP7_75t_SL g193 ( 
.A(n_161),
.Y(n_193)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_193),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

INVx6_ASAP7_75t_SL g281 ( 
.A(n_194),
.Y(n_281)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_195),
.Y(n_288)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_196),
.Y(n_259)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_197),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_149),
.A2(n_76),
.B1(n_111),
.B2(n_87),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_198),
.A2(n_205),
.B1(n_207),
.B2(n_225),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_88),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_199),
.B(n_212),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_200),
.Y(n_290)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_201),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_202),
.B(n_203),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_123),
.B(n_68),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_158),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_204),
.B(n_208),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_131),
.A2(n_71),
.B1(n_100),
.B2(n_74),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_206),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_171),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_129),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_129),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_210),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_95),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_164),
.A2(n_73),
.B(n_68),
.C(n_59),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_213),
.A2(n_245),
.B(n_190),
.C(n_189),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

INVx4_ASAP7_75t_SL g279 ( 
.A(n_214),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_155),
.B(n_90),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_215),
.B(n_227),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_135),
.A2(n_175),
.B1(n_180),
.B2(n_127),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_217),
.A2(n_231),
.B1(n_234),
.B2(n_146),
.Y(n_271)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_218),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_130),
.Y(n_219)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_93),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_159),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_221),
.B(n_222),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_144),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_224),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_178),
.A2(n_77),
.B1(n_6),
.B2(n_7),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_142),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_226),
.B(n_228),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_177),
.B(n_0),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_8),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_120),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_235),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_154),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_233),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_151),
.B(n_9),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_122),
.A2(n_10),
.B1(n_181),
.B2(n_179),
.Y(n_234)
);

OR2x2_ASAP7_75t_SL g235 ( 
.A(n_187),
.B(n_10),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_134),
.B(n_118),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_236),
.B(n_237),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_148),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g238 ( 
.A(n_121),
.B(n_182),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_239),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_118),
.B(n_169),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_169),
.B(n_187),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_126),
.B(n_121),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_242),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_136),
.B(n_145),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_145),
.B1(n_146),
.B2(n_152),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_137),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_152),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_126),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_248),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_141),
.B(n_153),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_124),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_160),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_173),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_208),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_207),
.A2(n_176),
.B1(n_140),
.B2(n_124),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_254),
.A2(n_258),
.B1(n_273),
.B2(n_274),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_154),
.B1(n_153),
.B2(n_141),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_260),
.B(n_224),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_170),
.C(n_160),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_261),
.B(n_294),
.C(n_280),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_271),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_191),
.A2(n_125),
.B1(n_138),
.B2(n_165),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_211),
.A2(n_138),
.B1(n_147),
.B2(n_173),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_235),
.B(n_147),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_283),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_189),
.B(n_137),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_230),
.A2(n_202),
.B1(n_248),
.B2(n_234),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_285),
.A2(n_297),
.B1(n_194),
.B2(n_188),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_193),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_197),
.B(n_218),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_201),
.B(n_229),
.C(n_196),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_195),
.A2(n_238),
.B1(n_249),
.B2(n_247),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_295),
.A2(n_241),
.B1(n_237),
.B2(n_223),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_233),
.A2(n_203),
.B1(n_221),
.B2(n_222),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_293),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_299),
.B(n_302),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_300),
.A2(n_305),
.B(n_317),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_257),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_206),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_307),
.B(n_315),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_311),
.Y(n_339)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_309),
.Y(n_365)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_247),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_267),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_312),
.B(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_276),
.Y(n_313)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_243),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_270),
.Y(n_316)
);

AOI222xp33_ASAP7_75t_L g317 ( 
.A1(n_252),
.A2(n_204),
.B1(n_224),
.B2(n_246),
.C1(n_192),
.C2(n_241),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_318),
.A2(n_321),
.B(n_325),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_200),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g349 ( 
.A(n_319),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_219),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_320),
.B(n_328),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_283),
.A2(n_224),
.B(n_241),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_250),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_322),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_323),
.A2(n_281),
.B1(n_276),
.B2(n_290),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_327),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_246),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_285),
.A2(n_210),
.B1(n_209),
.B2(n_214),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_326),
.A2(n_333),
.B1(n_269),
.B2(n_272),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_261),
.B(n_226),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_281),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_255),
.B(n_265),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_329),
.B(n_336),
.Y(n_362)
);

AO22x1_ASAP7_75t_L g330 ( 
.A1(n_253),
.A2(n_232),
.B1(n_254),
.B2(n_258),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_330),
.A2(n_292),
.B(n_279),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_332),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_256),
.B(n_266),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_265),
.A2(n_256),
.B1(n_291),
.B2(n_264),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_266),
.B(n_277),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_335),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_259),
.C(n_296),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_282),
.Y(n_336)
);

AOI22x1_ASAP7_75t_SL g337 ( 
.A1(n_333),
.A2(n_273),
.B1(n_274),
.B2(n_298),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_311),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_340),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_308),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_341),
.A2(n_347),
.B1(n_355),
.B2(n_359),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_314),
.A2(n_296),
.B1(n_275),
.B2(n_269),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_344),
.A2(n_345),
.B1(n_310),
.B2(n_303),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_263),
.B1(n_259),
.B2(n_288),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_326),
.A2(n_263),
.B1(n_288),
.B2(n_278),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_325),
.A2(n_290),
.B1(n_292),
.B2(n_279),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_334),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_301),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_363),
.Y(n_369)
);

AND2x2_ASAP7_75t_SL g363 ( 
.A(n_315),
.B(n_287),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_324),
.C(n_307),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_375),
.C(n_348),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_341),
.A2(n_304),
.B1(n_318),
.B2(n_299),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_368),
.A2(n_371),
.B1(n_385),
.B2(n_345),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_321),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_370),
.A2(n_383),
.B1(n_357),
.B2(n_356),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_338),
.A2(n_304),
.B1(n_306),
.B2(n_330),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_332),
.C(n_301),
.Y(n_372)
);

NAND3xp33_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_376),
.C(n_384),
.Y(n_403)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_340),
.B(n_306),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_378),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_327),
.C(n_331),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_350),
.B(n_335),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_377),
.A2(n_388),
.B1(n_359),
.B2(n_355),
.Y(n_402)
);

BUFx12_ASAP7_75t_L g378 ( 
.A(n_365),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_300),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_379),
.B(n_380),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_339),
.B(n_300),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_381),
.B(n_386),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_325),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_342),
.B(n_309),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_339),
.A2(n_330),
.B1(n_317),
.B2(n_313),
.Y(n_385)
);

NOR3xp33_ASAP7_75t_L g386 ( 
.A(n_342),
.B(n_322),
.C(n_251),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_287),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_344),
.B(n_250),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_R g398 ( 
.A(n_389),
.B(n_352),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_354),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_393),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_394),
.C(n_395),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_354),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_348),
.C(n_364),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_364),
.C(n_363),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_363),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_407),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_398),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_363),
.C(n_352),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_399),
.B(n_404),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_401),
.A2(n_377),
.B1(n_389),
.B2(n_337),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_402),
.A2(n_387),
.B1(n_368),
.B2(n_371),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_361),
.C(n_349),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_406),
.A2(n_370),
.B(n_369),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_366),
.B(n_362),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_382),
.A2(n_337),
.B1(n_356),
.B2(n_347),
.Y(n_408)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_408),
.Y(n_411)
);

BUFx24_ASAP7_75t_SL g409 ( 
.A(n_381),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_409),
.Y(n_410)
);

A2O1A1O1Ixp25_ASAP7_75t_L g412 ( 
.A1(n_399),
.A2(n_382),
.B(n_369),
.C(n_370),
.D(n_385),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_395),
.C(n_397),
.Y(n_427)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_396),
.Y(n_413)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_413),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_414),
.A2(n_405),
.B1(n_394),
.B2(n_407),
.Y(n_426)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_415),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_417),
.A2(n_373),
.B1(n_403),
.B2(n_343),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_418),
.A2(n_357),
.B(n_353),
.Y(n_435)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_400),
.Y(n_421)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_421),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_404),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_393),
.Y(n_428)
);

BUFx12_ASAP7_75t_L g423 ( 
.A(n_406),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_423),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_426),
.A2(n_424),
.B1(n_422),
.B2(n_411),
.Y(n_440)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_431),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_430),
.A2(n_414),
.B1(n_424),
.B2(n_417),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_392),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_421),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_438),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_391),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_435),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_346),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_436),
.B(n_416),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_439),
.B(n_440),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_433),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_442),
.B(n_429),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_444),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_420),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_419),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_430),
.A2(n_418),
.B(n_423),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_446),
.A2(n_412),
.B(n_425),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_451),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_450),
.Y(n_458)
);

INVx11_ASAP7_75t_L g453 ( 
.A(n_448),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_438),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_445),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_455),
.B(n_456),
.C(n_446),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_428),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_459),
.B(n_460),
.C(n_461),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_454),
.A2(n_447),
.B(n_441),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_452),
.A2(n_440),
.B1(n_423),
.B2(n_442),
.Y(n_462)
);

AOI322xp5_ASAP7_75t_L g463 ( 
.A1(n_462),
.A2(n_450),
.A3(n_442),
.B1(n_453),
.B2(n_451),
.C1(n_427),
.C2(n_456),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_463),
.A2(n_464),
.B1(n_465),
.B2(n_343),
.Y(n_468)
);

AOI322xp5_ASAP7_75t_L g464 ( 
.A1(n_458),
.A2(n_378),
.A3(n_432),
.B1(n_437),
.B2(n_416),
.C1(n_353),
.C2(n_419),
.Y(n_464)
);

AOI322xp5_ASAP7_75t_L g465 ( 
.A1(n_462),
.A2(n_378),
.A3(n_455),
.B1(n_365),
.B2(n_449),
.C1(n_343),
.C2(n_251),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_457),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_467),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_469),
.A2(n_468),
.B(n_262),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_470),
.B(n_262),
.Y(n_471)
);


endmodule