module real_jpeg_32493_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_0),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_0),
.Y(n_185)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_0),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_0),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_0),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_1),
.A2(n_38),
.B1(n_158),
.B2(n_163),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_1),
.A2(n_38),
.B1(n_289),
.B2(n_292),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_1),
.A2(n_38),
.B1(n_356),
.B2(n_359),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_2),
.A2(n_94),
.B1(n_97),
.B2(n_103),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_2),
.A2(n_103),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_2),
.A2(n_103),
.B1(n_179),
.B2(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_187),
.B1(n_188),
.B2(n_191),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_3),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_3),
.A2(n_187),
.B1(n_245),
.B2(n_249),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_5),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_6),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_6),
.Y(n_192)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_6),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_7),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

INVx2_ASAP7_75t_R g220 ( 
.A(n_7),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_8),
.A2(n_61),
.B(n_64),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_8),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_8),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_8),
.A2(n_172),
.B1(n_288),
.B2(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_8),
.B(n_145),
.Y(n_373)
);

OAI32xp33_ASAP7_75t_L g390 ( 
.A1(n_8),
.A2(n_121),
.A3(n_391),
.B1(n_396),
.B2(n_397),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_8),
.A2(n_194),
.B1(n_407),
.B2(n_410),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_9),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_9),
.A2(n_88),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_10),
.A2(n_136),
.B1(n_139),
.B2(n_143),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_10),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_10),
.A2(n_143),
.B1(n_260),
.B2(n_263),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_10),
.A2(n_143),
.B1(n_296),
.B2(n_298),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_10),
.A2(n_143),
.B1(n_377),
.B2(n_379),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_147),
.B1(n_152),
.B2(n_153),
.Y(n_146)
);

INVx2_ASAP7_75t_R g152 ( 
.A(n_11),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_11),
.A2(n_152),
.B1(n_320),
.B2(n_325),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_11),
.A2(n_152),
.B1(n_414),
.B2(n_417),
.Y(n_413)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_12),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_12),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_12),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_14),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_15),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_15),
.Y(n_235)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_16),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_16),
.Y(n_168)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_279),
.B1(n_445),
.B2(n_446),
.Y(n_18)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_19),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_277),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_228),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_21),
.B(n_228),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_155),
.C(n_195),
.Y(n_21)
);

XOR2x2_ASAP7_75t_L g441 ( 
.A(n_22),
.B(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_68),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJx2_ASAP7_75t_L g251 ( 
.A(n_24),
.B(n_69),
.C(n_113),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_37),
.B1(n_46),
.B2(n_60),
.Y(n_24)
);

NOR2xp67_ASAP7_75t_SL g193 ( 
.A(n_25),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_25),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_26)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_27),
.Y(n_120)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_29),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_29),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_29),
.Y(n_151)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_30),
.Y(n_208)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_31),
.Y(n_203)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_32),
.Y(n_154)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_32),
.Y(n_199)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_37),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_47),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_52),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_56),
.Y(n_262)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_63),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_64),
.Y(n_212)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_113),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_81),
.B1(n_93),
.B2(n_104),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_70),
.A2(n_81),
.B1(n_104),
.B2(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_70),
.B(n_194),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_70),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_70),
.A2(n_104),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_71),
.Y(n_420)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AO21x2_ASAP7_75t_L g104 ( 
.A1(n_72),
.A2(n_105),
.B(n_109),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_74),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_74),
.Y(n_346)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_75),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_75),
.Y(n_190)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_91),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_92),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_92),
.Y(n_378)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_93),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_101),
.Y(n_344)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_104),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_104),
.A2(n_431),
.B(n_432),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_109),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_135),
.B1(n_144),
.B2(n_146),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_135),
.B1(n_144),
.B2(n_157),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_114),
.A2(n_144),
.B1(n_146),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_114),
.A2(n_144),
.B1(n_157),
.B2(n_406),
.Y(n_405)
);

AO21x2_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_121),
.B(n_125),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_128),
.B1(n_130),
.B2(n_132),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_127),
.Y(n_399)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_127),
.Y(n_419)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_131),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_131),
.Y(n_382)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_138),
.Y(n_409)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_142),
.Y(n_411)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_155),
.B(n_195),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_169),
.C(n_193),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_156),
.B(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_161),
.Y(n_271)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_161),
.Y(n_395)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_168),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_169),
.A2(n_170),
.B1(n_193),
.B2(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_176),
.B1(n_183),
.B2(n_186),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_186),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_171),
.A2(n_317),
.B1(n_318),
.B2(n_326),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_171),
.A2(n_176),
.B1(n_370),
.B2(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_172),
.A2(n_216),
.B1(n_232),
.B2(n_238),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_172),
.A2(n_288),
.B1(n_295),
.B2(n_302),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_172),
.A2(n_319),
.B1(n_327),
.B2(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx4f_ASAP7_75t_L g312 ( 
.A(n_175),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_182),
.Y(n_291)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_182),
.Y(n_294)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_182),
.Y(n_301)
);

BUFx2_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_184),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_192),
.Y(n_336)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_193),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_194),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_194),
.B(n_343),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_SL g349 ( 
.A1(n_194),
.A2(n_342),
.B(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_194),
.B(n_398),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_213),
.B1(n_225),
.B2(n_227),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_196),
.B(n_227),
.Y(n_276)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_200),
.A3(n_204),
.B1(n_206),
.B2(n_212),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_200),
.A3(n_204),
.B1(n_206),
.B2(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_219),
.Y(n_371)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_252),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_251),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_276),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_267),
.B2(n_268),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_279),
.Y(n_446)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_440),
.B(n_444),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_425),
.B(n_439),
.Y(n_281)
);

AOI21x1_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_386),
.B(n_424),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_365),
.B(n_385),
.Y(n_283)
);

AOI22x1_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_315),
.B1(n_363),
.B2(n_364),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_305),
.B(n_314),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_304),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_287),
.B(n_304),
.Y(n_314)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_295),
.Y(n_317)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_302),
.Y(n_401)
);

INVx4_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_330),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_316),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_348),
.B2(n_362),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_331),
.B(n_362),
.Y(n_366)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_341),
.B1(n_345),
.B2(n_347),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_354),
.B1(n_355),
.B2(n_361),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_353),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_354),
.A2(n_413),
.B1(n_420),
.B2(n_421),
.Y(n_412)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_361),
.B(n_433),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_367),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_372),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_374),
.C(n_383),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_383),
.B2(n_384),
.Y(n_372)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_373),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_374),
.Y(n_384)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_376),
.Y(n_421)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_SL g424 ( 
.A(n_387),
.B(n_388),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_404),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_412),
.C(n_423),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_400),
.B1(n_402),
.B2(n_403),
.Y(n_389)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_390),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_390),
.B(n_403),
.Y(n_435)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_400),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_412),
.B1(n_422),
.B2(n_423),
.Y(n_404)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_405),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_412),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_413),
.Y(n_431)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_427),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_436),
.Y(n_427)
);

OA22x2_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_434),
.B2(n_435),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_434),
.C(n_436),
.Y(n_443)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

NOR2x1_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_443),
.Y(n_444)
);


endmodule