module fake_netlist_5_769_n_1465 (n_137, n_210, n_168, n_294, n_260, n_164, n_191, n_298, n_286, n_91, n_208, n_82, n_122, n_194, n_282, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_299, n_268, n_303, n_182, n_143, n_83, n_132, n_61, n_296, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_281, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_291, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_271, n_284, n_46, n_233, n_21, n_94, n_203, n_245, n_274, n_205, n_304, n_113, n_38, n_123, n_139, n_105, n_280, n_246, n_80, n_4, n_179, n_125, n_35, n_269, n_167, n_128, n_73, n_234, n_277, n_17, n_92, n_19, n_267, n_149, n_120, n_285, n_232, n_297, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_266, n_272, n_219, n_157, n_258, n_302, n_265, n_29, n_79, n_193, n_293, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_288, n_247, n_188, n_190, n_8, n_201, n_292, n_158, n_263, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_264, n_283, n_300, n_109, n_112, n_212, n_85, n_159, n_163, n_276, n_95, n_119, n_183, n_185, n_243, n_239, n_275, n_175, n_252, n_169, n_59, n_262, n_26, n_255, n_133, n_238, n_215, n_295, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_290, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_273, n_287, n_270, n_222, n_230, n_81, n_118, n_28, n_89, n_301, n_279, n_70, n_115, n_68, n_93, n_253, n_261, n_72, n_174, n_186, n_199, n_289, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_305, n_204, n_50, n_250, n_52, n_278, n_88, n_110, n_216, n_1465);

input n_137;
input n_210;
input n_168;
input n_294;
input n_260;
input n_164;
input n_191;
input n_298;
input n_286;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_282;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_299;
input n_268;
input n_303;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_296;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_281;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_291;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_271;
input n_284;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_274;
input n_205;
input n_304;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_280;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_269;
input n_167;
input n_128;
input n_73;
input n_234;
input n_277;
input n_17;
input n_92;
input n_19;
input n_267;
input n_149;
input n_120;
input n_285;
input n_232;
input n_297;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_266;
input n_272;
input n_219;
input n_157;
input n_258;
input n_302;
input n_265;
input n_29;
input n_79;
input n_193;
input n_293;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_288;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_292;
input n_158;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_264;
input n_283;
input n_300;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_276;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_275;
input n_175;
input n_252;
input n_169;
input n_59;
input n_262;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_295;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_290;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_273;
input n_287;
input n_270;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_301;
input n_279;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_261;
input n_72;
input n_174;
input n_186;
input n_199;
input n_289;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_305;
input n_204;
input n_50;
input n_250;
input n_52;
input n_278;
input n_88;
input n_110;
input n_216;

output n_1465;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1314;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1078;
wire n_775;
wire n_600;
wire n_1374;
wire n_1328;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_1058;
wire n_586;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_851;
wire n_615;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_1270;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_318;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_48),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_220),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_184),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_53),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_164),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_144),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_102),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_108),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_231),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_141),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_203),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_25),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_14),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_15),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_291),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_158),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_198),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_4),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_36),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_209),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_48),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_208),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_276),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_149),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_79),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_116),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_168),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_241),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_148),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_159),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_166),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_304),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_67),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_134),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_249),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_246),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_77),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_252),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_305),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_269),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_120),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_107),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_265),
.Y(n_353)
);

BUFx8_ASAP7_75t_SL g354 ( 
.A(n_44),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_97),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_255),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_211),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_10),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_224),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_239),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_193),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_37),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_267),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_167),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_21),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_242),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_272),
.Y(n_368)
);

BUFx10_ASAP7_75t_L g369 ( 
.A(n_21),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_152),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_187),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_263),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_240),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_99),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_190),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_126),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_282),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_57),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_8),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_214),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_113),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_228),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_47),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_140),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_143),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_243),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_182),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_54),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_83),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_62),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_284),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_50),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_41),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_177),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_118),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_281),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_247),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_154),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_205),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_188),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_271),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_174),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_175),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_261),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_106),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_122),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_46),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_248),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_125),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_296),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_206),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_297),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_86),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_31),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_219),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_300),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_55),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_60),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_229),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_9),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_178),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_91),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_100),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_0),
.Y(n_424)
);

BUFx10_ASAP7_75t_L g425 ( 
.A(n_257),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_57),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_70),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_234),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_238),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_41),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_33),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_194),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_78),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_128),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_49),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_227),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_109),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_12),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_96),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_288),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_266),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_89),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_96),
.Y(n_443)
);

INVxp33_ASAP7_75t_L g444 ( 
.A(n_1),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_283),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_119),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_43),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_63),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_191),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_192),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_244),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_58),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_207),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_279),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_299),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_74),
.Y(n_456)
);

INVxp33_ASAP7_75t_SL g457 ( 
.A(n_200),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_210),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_287),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_14),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_176),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_254),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_222),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_29),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_112),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_39),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_95),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_233),
.Y(n_468)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_138),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_83),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_77),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_27),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_173),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_280),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_199),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_186),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_196),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_80),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_62),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_24),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_36),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_146),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_295),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_195),
.Y(n_484)
);

BUFx5_ASAP7_75t_L g485 ( 
.A(n_163),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_230),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_39),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_226),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_189),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_251),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_301),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_121),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_63),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_245),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_250),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_71),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_129),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_81),
.Y(n_498)
);

BUFx5_ASAP7_75t_L g499 ( 
.A(n_237),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_26),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_117),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_278),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_25),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_127),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_312),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_354),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_347),
.B(n_0),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_374),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_418),
.Y(n_509)
);

BUFx12f_ASAP7_75t_L g510 ( 
.A(n_321),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_347),
.B(n_1),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_338),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_354),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_312),
.B(n_2),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

BUFx8_ASAP7_75t_L g516 ( 
.A(n_384),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_338),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_341),
.B(n_2),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_418),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_471),
.B(n_3),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_374),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_306),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_338),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_379),
.Y(n_524)
);

BUFx12f_ASAP7_75t_L g525 ( 
.A(n_321),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_338),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_404),
.B(n_3),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_418),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_341),
.B(n_4),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_409),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_314),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_413),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_318),
.B(n_5),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_318),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_332),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_404),
.B(n_402),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_449),
.B(n_5),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_368),
.B(n_6),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_379),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_438),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_409),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_423),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_332),
.B(n_7),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_409),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_413),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_409),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_368),
.B(n_101),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_315),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_416),
.B(n_8),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_405),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_423),
.Y(n_551)
);

BUFx12f_ASAP7_75t_L g552 ( 
.A(n_369),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_423),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_457),
.B(n_9),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_405),
.B(n_10),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_469),
.B(n_444),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_441),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_441),
.B(n_11),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_459),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_416),
.B(n_11),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_444),
.B(n_12),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_423),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_426),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_459),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_491),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_491),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_455),
.B(n_13),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_426),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_455),
.B(n_15),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_327),
.B(n_391),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_426),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_479),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_479),
.B(n_16),
.Y(n_575)
);

BUFx12f_ASAP7_75t_L g576 ( 
.A(n_448),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_307),
.B(n_103),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_400),
.B(n_16),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_396),
.B(n_483),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_479),
.Y(n_580)
);

INVx6_ASAP7_75t_L g581 ( 
.A(n_425),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_311),
.Y(n_582)
);

INVx5_ASAP7_75t_L g583 ( 
.A(n_425),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_388),
.B(n_17),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_324),
.B(n_17),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_309),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_317),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_310),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_325),
.B(n_18),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_425),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_372),
.B(n_18),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_323),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_448),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_313),
.B(n_19),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_319),
.B(n_20),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_329),
.B(n_20),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_363),
.B(n_22),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_448),
.B(n_22),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_378),
.B(n_23),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_456),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_330),
.B(n_26),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_393),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_407),
.B(n_28),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_414),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_420),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_339),
.B(n_28),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_429),
.B(n_29),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_485),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_340),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_345),
.B(n_104),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_346),
.B(n_30),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_456),
.B(n_30),
.Y(n_612)
);

BUFx12f_ASAP7_75t_L g613 ( 
.A(n_465),
.Y(n_613)
);

BUFx12f_ASAP7_75t_L g614 ( 
.A(n_465),
.Y(n_614)
);

BUFx12f_ASAP7_75t_L g615 ( 
.A(n_465),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_431),
.B(n_31),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_308),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_435),
.B(n_32),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_442),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_473),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g621 ( 
.A(n_424),
.B(n_32),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_452),
.B(n_33),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_361),
.Y(n_623)
);

INVxp33_ASAP7_75t_SL g624 ( 
.A(n_322),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_473),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_367),
.B(n_34),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_460),
.B(n_34),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_467),
.B(n_35),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_453),
.B(n_35),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_478),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_476),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_370),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_476),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_487),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_476),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_490),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_485),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_371),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_493),
.B(n_37),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_485),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_490),
.B(n_38),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_496),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_503),
.B(n_38),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_485),
.Y(n_644)
);

BUFx12f_ASAP7_75t_L g645 ( 
.A(n_490),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_373),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_328),
.B(n_40),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_474),
.B(n_42),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_320),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_375),
.B(n_43),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_376),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_380),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_485),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_569),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_556),
.A2(n_428),
.B1(n_437),
.B2(n_406),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_579),
.A2(n_482),
.B1(n_495),
.B2(n_462),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_509),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_507),
.A2(n_343),
.B1(n_355),
.B2(n_331),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_536),
.B(n_326),
.Y(n_659)
);

AO22x2_ASAP7_75t_L g660 ( 
.A1(n_641),
.A2(n_422),
.B1(n_430),
.B2(n_335),
.Y(n_660)
);

AO22x2_ASAP7_75t_L g661 ( 
.A1(n_514),
.A2(n_470),
.B1(n_394),
.B2(n_398),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_520),
.A2(n_366),
.B1(n_383),
.B2(n_358),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_620),
.B(n_385),
.Y(n_663)
);

AO22x2_ASAP7_75t_L g664 ( 
.A1(n_514),
.A2(n_401),
.B1(n_408),
.B2(n_399),
.Y(n_664)
);

AO22x2_ASAP7_75t_L g665 ( 
.A1(n_533),
.A2(n_415),
.B1(n_419),
.B2(n_411),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_SL g666 ( 
.A1(n_520),
.A2(n_390),
.B1(n_392),
.B2(n_389),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_621),
.A2(n_427),
.B1(n_433),
.B2(n_417),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_617),
.B(n_333),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_515),
.Y(n_669)
);

AO22x1_ASAP7_75t_SL g670 ( 
.A1(n_568),
.A2(n_436),
.B1(n_440),
.B2(n_421),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_620),
.B(n_334),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_569),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_521),
.B(n_336),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_507),
.A2(n_443),
.B1(n_447),
.B2(n_439),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_505),
.B(n_534),
.Y(n_675)
);

AO22x2_ASAP7_75t_L g676 ( 
.A1(n_533),
.A2(n_446),
.B1(n_454),
.B2(n_445),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_593),
.B(n_480),
.Y(n_677)
);

OA22x2_ASAP7_75t_L g678 ( 
.A1(n_508),
.A2(n_498),
.B1(n_500),
.B2(n_481),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_527),
.A2(n_466),
.B1(n_472),
.B2(n_464),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_569),
.Y(n_680)
);

AO22x2_ASAP7_75t_L g681 ( 
.A1(n_543),
.A2(n_468),
.B1(n_477),
.B2(n_463),
.Y(n_681)
);

NAND3x1_ASAP7_75t_L g682 ( 
.A(n_511),
.B(n_488),
.C(n_486),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_554),
.A2(n_337),
.B1(n_344),
.B2(n_342),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_L g684 ( 
.A1(n_621),
.A2(n_501),
.B1(n_349),
.B2(n_350),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_513),
.B(n_44),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_537),
.B(n_568),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_535),
.B(n_348),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_629),
.A2(n_351),
.B1(n_353),
.B2(n_352),
.Y(n_688)
);

OA22x2_ASAP7_75t_L g689 ( 
.A1(n_532),
.A2(n_356),
.B1(n_359),
.B2(n_357),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_542),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_593),
.B(n_360),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_648),
.A2(n_362),
.B1(n_365),
.B2(n_364),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_551),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_562),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_572),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_574),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_573),
.Y(n_697)
);

AO22x2_ASAP7_75t_L g698 ( 
.A1(n_543),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_624),
.B(n_377),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_522),
.B(n_381),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_573),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_573),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_519),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_557),
.B(n_45),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_SL g705 ( 
.A1(n_581),
.A2(n_382),
.B1(n_387),
.B2(n_386),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_531),
.B(n_548),
.Y(n_706)
);

AO22x2_ASAP7_75t_L g707 ( 
.A1(n_555),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_519),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_557),
.B(n_52),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_528),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_SL g711 ( 
.A1(n_647),
.A2(n_591),
.B1(n_529),
.B2(n_538),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_506),
.Y(n_712)
);

AOI22x1_ASAP7_75t_L g713 ( 
.A1(n_570),
.A2(n_504),
.B1(n_502),
.B2(n_395),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_528),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_512),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_553),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_566),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_585),
.A2(n_461),
.B1(n_497),
.B2(n_494),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_589),
.A2(n_451),
.B1(n_492),
.B2(n_489),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_512),
.Y(n_720)
);

OAI22xp33_ASAP7_75t_SL g721 ( 
.A1(n_518),
.A2(n_529),
.B1(n_549),
.B2(n_538),
.Y(n_721)
);

AO22x2_ASAP7_75t_L g722 ( 
.A1(n_555),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_583),
.B(n_397),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_583),
.B(n_403),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_561),
.A2(n_458),
.B1(n_410),
.B2(n_484),
.Y(n_725)
);

AO22x2_ASAP7_75t_L g726 ( 
.A1(n_558),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_726)
);

AO22x2_ASAP7_75t_L g727 ( 
.A1(n_558),
.A2(n_56),
.B1(n_59),
.B2(n_61),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_583),
.B(n_590),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_589),
.A2(n_450),
.B1(n_412),
.B2(n_475),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_512),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_517),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_517),
.Y(n_732)
);

AO22x2_ASAP7_75t_L g733 ( 
.A1(n_578),
.A2(n_59),
.B1(n_61),
.B2(n_64),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_650),
.A2(n_560),
.B1(n_600),
.B2(n_590),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_517),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_587),
.B(n_432),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_523),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_523),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_625),
.B(n_434),
.Y(n_739)
);

AO22x2_ASAP7_75t_L g740 ( 
.A1(n_578),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_625),
.B(n_485),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_607),
.A2(n_499),
.B1(n_316),
.B2(n_67),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_650),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_625),
.B(n_499),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_550),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_550),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_649),
.B(n_316),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_675),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_684),
.B(n_721),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_655),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_730),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_728),
.B(n_633),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_711),
.B(n_567),
.Y(n_753)
);

XNOR2x1_ASAP7_75t_L g754 ( 
.A(n_679),
.B(n_584),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_730),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_712),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_731),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_698),
.B(n_510),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_720),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_732),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_735),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_673),
.Y(n_762)
);

AOI21x1_ASAP7_75t_L g763 ( 
.A1(n_747),
.A2(n_637),
.B(n_608),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_737),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_738),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_677),
.B(n_567),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_672),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_657),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_672),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_712),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_686),
.A2(n_610),
.B(n_577),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_659),
.B(n_633),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_656),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_662),
.B(n_633),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_701),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_701),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_687),
.B(n_635),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_702),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_654),
.Y(n_779)
);

INVx3_ASAP7_75t_R g780 ( 
.A(n_691),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_669),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_654),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_745),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_746),
.Y(n_784)
);

XOR2x2_ASAP7_75t_L g785 ( 
.A(n_666),
.B(n_598),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_680),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_715),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_691),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_678),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_688),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_700),
.A2(n_541),
.B(n_530),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_716),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_715),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_736),
.A2(n_541),
.B(n_530),
.Y(n_794)
);

INVxp67_ASAP7_75t_SL g795 ( 
.A(n_715),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_668),
.B(n_635),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_708),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_714),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_690),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_689),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_693),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_671),
.B(n_636),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_694),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_695),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_696),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_703),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_703),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_710),
.Y(n_808)
);

AND2x2_ASAP7_75t_SL g809 ( 
.A(n_742),
.B(n_570),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_661),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_744),
.A2(n_706),
.B(n_741),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_SL g812 ( 
.A(n_658),
.B(n_612),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_710),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_692),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_697),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_697),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_697),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_699),
.B(n_636),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_685),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_717),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_667),
.B(n_571),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_725),
.B(n_571),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_663),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_704),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_709),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_682),
.Y(n_826)
);

XNOR2x2_ASAP7_75t_L g827 ( 
.A(n_733),
.B(n_596),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_670),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_664),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_664),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_665),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_665),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_686),
.B(n_723),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_683),
.B(n_541),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_676),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_676),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_724),
.B(n_550),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_681),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_686),
.B(n_594),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_718),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_837),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_806),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_748),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_839),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_768),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_839),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_823),
.B(n_681),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_753),
.B(n_661),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_766),
.B(n_686),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_753),
.B(n_660),
.Y(n_850)
);

AND2x2_ASAP7_75t_SL g851 ( 
.A(n_749),
.B(n_809),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_807),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_839),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_788),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_788),
.B(n_800),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_768),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_749),
.B(n_739),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_781),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_770),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_789),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_811),
.B(n_719),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_796),
.B(n_660),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_793),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_808),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_781),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_813),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_762),
.B(n_733),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_751),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_755),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_792),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_818),
.B(n_729),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_821),
.B(n_740),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_767),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_821),
.B(n_740),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_800),
.B(n_595),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_763),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_769),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_770),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_799),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_815),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_801),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_833),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_816),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_824),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_825),
.B(n_698),
.Y(n_885)
);

AND2x2_ASAP7_75t_SL g886 ( 
.A(n_809),
.B(n_595),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_772),
.B(n_707),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_775),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_829),
.B(n_601),
.Y(n_889)
);

INVx4_ASAP7_75t_L g890 ( 
.A(n_776),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_803),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_777),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_756),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_759),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_804),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_822),
.B(n_707),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_760),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_774),
.B(n_713),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_830),
.B(n_601),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_822),
.B(n_790),
.Y(n_900)
);

AND2x6_ASAP7_75t_L g901 ( 
.A(n_831),
.B(n_606),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_805),
.Y(n_902)
);

AND2x4_ASAP7_75t_SL g903 ( 
.A(n_758),
.B(n_685),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_832),
.B(n_606),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_797),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_820),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_812),
.A2(n_674),
.B1(n_577),
.B2(n_610),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_835),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_817),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_798),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_761),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_764),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_810),
.B(n_734),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_802),
.B(n_722),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_765),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_836),
.B(n_722),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_826),
.B(n_834),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_838),
.B(n_726),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_812),
.B(n_713),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_810),
.B(n_726),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_778),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_757),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_752),
.B(n_786),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_783),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_758),
.B(n_727),
.Y(n_925)
);

NAND2x1p5_ASAP7_75t_L g926 ( 
.A(n_784),
.B(n_611),
.Y(n_926)
);

AND2x2_ASAP7_75t_SL g927 ( 
.A(n_827),
.B(n_611),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_758),
.B(n_727),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_771),
.A2(n_610),
.B(n_577),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_779),
.Y(n_930)
);

INVxp67_ASAP7_75t_SL g931 ( 
.A(n_787),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_782),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_785),
.B(n_545),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_827),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_795),
.B(n_577),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_790),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_814),
.B(n_524),
.Y(n_937)
);

BUFx4f_ASAP7_75t_L g938 ( 
.A(n_936),
.Y(n_938)
);

OR2x6_ASAP7_75t_L g939 ( 
.A(n_936),
.B(n_819),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_855),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_937),
.B(n_754),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_853),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_936),
.B(n_934),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_937),
.B(n_750),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_853),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_855),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_845),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_853),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_857),
.B(n_814),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_853),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_841),
.B(n_840),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_841),
.B(n_840),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_854),
.B(n_582),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_SL g954 ( 
.A(n_886),
.B(n_927),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_854),
.B(n_780),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_845),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_898),
.B(n_882),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_882),
.B(n_773),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_853),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_855),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_893),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_900),
.B(n_773),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_846),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_842),
.B(n_626),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_844),
.B(n_559),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_856),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_860),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_884),
.Y(n_968)
);

NOR2x1_ASAP7_75t_L g969 ( 
.A(n_849),
.B(n_844),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_844),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_856),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_842),
.B(n_626),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_843),
.B(n_592),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_888),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_843),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_888),
.Y(n_976)
);

NAND2xp33_ASAP7_75t_L g977 ( 
.A(n_846),
.B(n_610),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_878),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_858),
.Y(n_979)
);

NAND2x1_ASAP7_75t_SL g980 ( 
.A(n_925),
.B(n_605),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_892),
.B(n_602),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_888),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_858),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_865),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_908),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_888),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_865),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_892),
.B(n_604),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_892),
.B(n_619),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_932),
.B(n_634),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_932),
.B(n_828),
.Y(n_991)
);

BUFx8_ASAP7_75t_L g992 ( 
.A(n_925),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_868),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_888),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_889),
.B(n_828),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_852),
.B(n_705),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_889),
.B(n_904),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_889),
.B(n_596),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_884),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_904),
.B(n_870),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_904),
.B(n_852),
.Y(n_1001)
);

INVx4_ASAP7_75t_L g1002 ( 
.A(n_863),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_864),
.B(n_875),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_893),
.Y(n_1004)
);

BUFx4f_ASAP7_75t_SL g1005 ( 
.A(n_859),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_L g1006 ( 
.A(n_861),
.B(n_791),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_882),
.B(n_743),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_864),
.B(n_597),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_875),
.B(n_597),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_868),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_936),
.B(n_630),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_882),
.B(n_640),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_882),
.B(n_919),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_863),
.Y(n_1014)
);

INVxp67_ASAP7_75t_SL g1015 ( 
.A(n_931),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_936),
.B(n_630),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_875),
.B(n_599),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_877),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_967),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_980),
.Y(n_1020)
);

OR2x6_ASAP7_75t_L g1021 ( 
.A(n_943),
.B(n_958),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1010),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1010),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_1005),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_948),
.Y(n_1025)
);

CKINVDCx11_ASAP7_75t_R g1026 ( 
.A(n_961),
.Y(n_1026)
);

BUFx12f_ASAP7_75t_L g1027 ( 
.A(n_1004),
.Y(n_1027)
);

BUFx4_ASAP7_75t_SL g1028 ( 
.A(n_939),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_971),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_978),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_971),
.Y(n_1031)
);

INVx6_ASAP7_75t_L g1032 ( 
.A(n_948),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_938),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_979),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_979),
.Y(n_1035)
);

BUFx2_ASAP7_75t_SL g1036 ( 
.A(n_975),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_985),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_938),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_984),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_984),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_982),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_987),
.Y(n_1042)
);

BUFx12f_ASAP7_75t_L g1043 ( 
.A(n_992),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_1011),
.Y(n_1044)
);

INVx8_ASAP7_75t_L g1045 ( 
.A(n_948),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1008),
.B(n_851),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1008),
.B(n_851),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_949),
.A2(n_886),
.B1(n_934),
.B2(n_871),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_987),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_947),
.Y(n_1050)
);

BUFx4_ASAP7_75t_SL g1051 ( 
.A(n_939),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_950),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_943),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_993),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_944),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_992),
.Y(n_1056)
);

BUFx4f_ASAP7_75t_L g1057 ( 
.A(n_950),
.Y(n_1057)
);

INVxp67_ASAP7_75t_SL g1058 ( 
.A(n_950),
.Y(n_1058)
);

AO21x2_ASAP7_75t_L g1059 ( 
.A1(n_957),
.A2(n_929),
.B(n_907),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_956),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1018),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_959),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_974),
.B(n_866),
.Y(n_1063)
);

BUFx4_ASAP7_75t_SL g1064 ( 
.A(n_941),
.Y(n_1064)
);

INVx3_ASAP7_75t_SL g1065 ( 
.A(n_995),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_974),
.B(n_866),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_970),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_982),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_970),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_1016),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_959),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_951),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_962),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_966),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_1014),
.Y(n_1075)
);

BUFx12f_ASAP7_75t_L g1076 ( 
.A(n_995),
.Y(n_1076)
);

OR2x6_ASAP7_75t_L g1077 ( 
.A(n_958),
.B(n_906),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_951),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_982),
.Y(n_1079)
);

NAND2x1p5_ASAP7_75t_L g1080 ( 
.A(n_976),
.B(n_866),
.Y(n_1080)
);

OR2x6_ASAP7_75t_L g1081 ( 
.A(n_959),
.B(n_906),
.Y(n_1081)
);

INVxp67_ASAP7_75t_SL g1082 ( 
.A(n_986),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_983),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_952),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_952),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_1014),
.Y(n_1086)
);

BUFx12f_ASAP7_75t_L g1087 ( 
.A(n_991),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_986),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1003),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_986),
.Y(n_1090)
);

BUFx4f_ASAP7_75t_SL g1091 ( 
.A(n_991),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1039),
.Y(n_1092)
);

INVx6_ASAP7_75t_L g1093 ( 
.A(n_1045),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_SL g1094 ( 
.A1(n_1073),
.A2(n_954),
.B1(n_933),
.B2(n_896),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1039),
.Y(n_1095)
);

BUFx8_ASAP7_75t_SL g1096 ( 
.A(n_1027),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1022),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1075),
.B(n_1086),
.Y(n_1098)
);

BUFx4f_ASAP7_75t_L g1099 ( 
.A(n_1027),
.Y(n_1099)
);

CKINVDCx11_ASAP7_75t_R g1100 ( 
.A(n_1026),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1048),
.A2(n_1007),
.B1(n_957),
.B2(n_896),
.Y(n_1101)
);

CKINVDCx16_ASAP7_75t_R g1102 ( 
.A(n_1043),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_1019),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1033),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1046),
.A2(n_1007),
.B1(n_874),
.B2(n_872),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_1067),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1040),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_1030),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_1030),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1047),
.A2(n_933),
.B1(n_874),
.B2(n_872),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1019),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_SL g1112 ( 
.A1(n_1044),
.A2(n_850),
.B(n_848),
.Y(n_1112)
);

BUFx4_ASAP7_75t_SL g1113 ( 
.A(n_1075),
.Y(n_1113)
);

BUFx8_ASAP7_75t_SL g1114 ( 
.A(n_1043),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1023),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1021),
.A2(n_1013),
.B1(n_972),
.B2(n_964),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1040),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1049),
.Y(n_1118)
);

INVx6_ASAP7_75t_L g1119 ( 
.A(n_1045),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1049),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1029),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1021),
.A2(n_1013),
.B1(n_996),
.B2(n_1015),
.Y(n_1122)
);

INVx6_ASAP7_75t_L g1123 ( 
.A(n_1045),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_SL g1124 ( 
.A1(n_1055),
.A2(n_1091),
.B1(n_1085),
.B2(n_1065),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_1070),
.A2(n_850),
.B1(n_848),
.B2(n_1001),
.Y(n_1125)
);

OAI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1055),
.A2(n_917),
.B1(n_968),
.B2(n_999),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1077),
.A2(n_1001),
.B1(n_1000),
.B2(n_998),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1031),
.Y(n_1128)
);

CKINVDCx11_ASAP7_75t_R g1129 ( 
.A(n_1026),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1077),
.A2(n_1000),
.B1(n_998),
.B2(n_1009),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_SL g1131 ( 
.A1(n_1087),
.A2(n_756),
.B1(n_516),
.B2(n_614),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1050),
.Y(n_1132)
);

CKINVDCx6p67_ASAP7_75t_R g1133 ( 
.A(n_1056),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_1024),
.Y(n_1134)
);

INVx6_ASAP7_75t_L g1135 ( 
.A(n_1045),
.Y(n_1135)
);

INVx6_ASAP7_75t_L g1136 ( 
.A(n_1033),
.Y(n_1136)
);

BUFx10_ASAP7_75t_L g1137 ( 
.A(n_1085),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1072),
.Y(n_1138)
);

CKINVDCx11_ASAP7_75t_R g1139 ( 
.A(n_1056),
.Y(n_1139)
);

OAI21xp33_ASAP7_75t_SL g1140 ( 
.A1(n_1077),
.A2(n_1035),
.B(n_1034),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_SL g1141 ( 
.A1(n_1065),
.A2(n_955),
.B1(n_615),
.B2(n_631),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1021),
.A2(n_1017),
.B1(n_997),
.B2(n_847),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1020),
.A2(n_847),
.B1(n_988),
.B2(n_981),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1042),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1078),
.A2(n_988),
.B1(n_989),
.B2(n_981),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_SL g1146 ( 
.A1(n_1087),
.A2(n_516),
.B1(n_645),
.B2(n_613),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1089),
.A2(n_989),
.B1(n_940),
.B2(n_946),
.Y(n_1147)
);

BUFx4_ASAP7_75t_R g1148 ( 
.A(n_1038),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1050),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1060),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1060),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_1037),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1086),
.Y(n_1153)
);

BUFx4f_ASAP7_75t_L g1154 ( 
.A(n_1076),
.Y(n_1154)
);

BUFx12f_ASAP7_75t_L g1155 ( 
.A(n_1076),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1083),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1084),
.A2(n_973),
.B1(n_867),
.B2(n_862),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1053),
.A2(n_990),
.B1(n_953),
.B2(n_960),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_SL g1159 ( 
.A1(n_1036),
.A2(n_903),
.B1(n_928),
.B2(n_885),
.Y(n_1159)
);

INVx8_ASAP7_75t_L g1160 ( 
.A(n_1081),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1054),
.A2(n_990),
.B1(n_953),
.B2(n_960),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1094),
.B(n_920),
.Y(n_1162)
);

BUFx4f_ASAP7_75t_SL g1163 ( 
.A(n_1108),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_1111),
.Y(n_1164)
);

INVx6_ASAP7_75t_L g1165 ( 
.A(n_1093),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1094),
.A2(n_1002),
.B1(n_1038),
.B2(n_1014),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1105),
.A2(n_1101),
.B1(n_1110),
.B2(n_1125),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1092),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1095),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1100),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1107),
.Y(n_1171)
);

AND2x4_ASAP7_75t_SL g1172 ( 
.A(n_1109),
.B(n_1137),
.Y(n_1172)
);

OAI222xp33_ASAP7_75t_L g1173 ( 
.A1(n_1101),
.A2(n_639),
.B1(n_616),
.B2(n_622),
.C1(n_627),
.C2(n_603),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1112),
.B(n_913),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1145),
.A2(n_1081),
.B1(n_1057),
.B2(n_1066),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1142),
.A2(n_873),
.B1(n_890),
.B2(n_869),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1097),
.Y(n_1177)
);

INVx6_ASAP7_75t_L g1178 ( 
.A(n_1093),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1154),
.A2(n_928),
.B1(n_525),
.B2(n_552),
.Y(n_1179)
);

OAI21xp33_ASAP7_75t_L g1180 ( 
.A1(n_1143),
.A2(n_923),
.B(n_895),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1157),
.A2(n_575),
.B1(n_618),
.B2(n_616),
.Y(n_1181)
);

BUFx12f_ASAP7_75t_L g1182 ( 
.A(n_1139),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1152),
.B(n_1158),
.Y(n_1183)
);

INVx5_ASAP7_75t_SL g1184 ( 
.A(n_1133),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_1134),
.B(n_1057),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1117),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1159),
.A2(n_1130),
.B1(n_1161),
.B2(n_1126),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1115),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1121),
.Y(n_1189)
);

AOI222xp33_ASAP7_75t_L g1190 ( 
.A1(n_1124),
.A2(n_642),
.B1(n_622),
.B2(n_643),
.C1(n_627),
.C2(n_639),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1159),
.A2(n_1081),
.B1(n_1057),
.B2(n_1066),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1128),
.Y(n_1192)
);

NOR2x1_ASAP7_75t_SL g1193 ( 
.A(n_1116),
.B(n_1081),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1118),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1144),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1098),
.B(n_1025),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1131),
.A2(n_576),
.B1(n_1064),
.B2(n_913),
.Y(n_1197)
);

INVx4_ASAP7_75t_L g1198 ( 
.A(n_1148),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_L g1199 ( 
.A(n_1147),
.B(n_628),
.C(n_642),
.Y(n_1199)
);

INVx6_ASAP7_75t_L g1200 ( 
.A(n_1093),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1122),
.A2(n_881),
.B1(n_891),
.B2(n_879),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1127),
.A2(n_1063),
.B1(n_1080),
.B2(n_976),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1122),
.A2(n_1061),
.B1(n_539),
.B2(n_924),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1129),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1149),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1136),
.A2(n_1080),
.B1(n_1063),
.B2(n_926),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1138),
.B(n_885),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1151),
.A2(n_539),
.B1(n_924),
.B2(n_902),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1156),
.A2(n_902),
.B1(n_891),
.B2(n_1059),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1120),
.A2(n_1059),
.B1(n_910),
.B2(n_905),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1153),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1155),
.A2(n_910),
.B1(n_905),
.B2(n_969),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1136),
.A2(n_926),
.B1(n_963),
.B2(n_1067),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1113),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1096),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1114),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1132),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1098),
.B(n_887),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1154),
.A2(n_969),
.B1(n_877),
.B2(n_883),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1136),
.A2(n_926),
.B1(n_963),
.B2(n_1067),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1103),
.B(n_887),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1150),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1104),
.B(n_914),
.Y(n_1223)
);

OAI222xp33_ASAP7_75t_L g1224 ( 
.A1(n_1187),
.A2(n_1146),
.B1(n_1074),
.B2(n_540),
.C1(n_1102),
.C2(n_914),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1197),
.A2(n_1160),
.B1(n_1099),
.B2(n_1141),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1174),
.B(n_1104),
.Y(n_1226)
);

NOR3xp33_ASAP7_75t_L g1227 ( 
.A(n_1173),
.B(n_1140),
.C(n_540),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1205),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1162),
.A2(n_1160),
.B1(n_1099),
.B2(n_1104),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1167),
.A2(n_915),
.B1(n_921),
.B2(n_911),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1190),
.A2(n_547),
.B1(n_963),
.B2(n_564),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1198),
.A2(n_1123),
.B1(n_1135),
.B2(n_1119),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1181),
.A2(n_565),
.B1(n_915),
.B2(n_911),
.Y(n_1233)
);

AO22x1_ASAP7_75t_L g1234 ( 
.A1(n_1191),
.A2(n_1058),
.B1(n_1082),
.B2(n_1106),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1164),
.B(n_1083),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_L g1236 ( 
.A(n_1181),
.B(n_1199),
.C(n_1203),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1183),
.A2(n_1123),
.B1(n_1135),
.B2(n_1119),
.Y(n_1237)
);

NOR3xp33_ASAP7_75t_L g1238 ( 
.A(n_1179),
.B(n_1006),
.C(n_897),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1193),
.A2(n_1106),
.B1(n_1059),
.B2(n_1069),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1180),
.A2(n_565),
.B1(n_883),
.B2(n_880),
.Y(n_1240)
);

NAND2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1185),
.B(n_1175),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1211),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1166),
.A2(n_909),
.B1(n_880),
.B2(n_897),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1221),
.A2(n_909),
.B1(n_894),
.B2(n_922),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1163),
.A2(n_1069),
.B1(n_901),
.B2(n_1119),
.Y(n_1245)
);

NOR3xp33_ASAP7_75t_L g1246 ( 
.A(n_1179),
.B(n_894),
.C(n_912),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1218),
.A2(n_930),
.B1(n_922),
.B2(n_912),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1203),
.B(n_1090),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1201),
.A2(n_930),
.B1(n_912),
.B2(n_901),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1212),
.A2(n_901),
.B1(n_316),
.B2(n_499),
.Y(n_1250)
);

OAI211xp5_ASAP7_75t_L g1251 ( 
.A1(n_1207),
.A2(n_918),
.B(n_916),
.C(n_586),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1177),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1176),
.A2(n_901),
.B1(n_316),
.B2(n_499),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1188),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1219),
.A2(n_901),
.B1(n_316),
.B2(n_499),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1163),
.A2(n_316),
.B1(n_499),
.B2(n_945),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1223),
.A2(n_942),
.B1(n_945),
.B2(n_965),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1202),
.A2(n_942),
.B1(n_994),
.B2(n_1012),
.Y(n_1258)
);

NOR3xp33_ASAP7_75t_L g1259 ( 
.A(n_1206),
.B(n_1052),
.C(n_1025),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1208),
.A2(n_994),
.B1(n_1012),
.B2(n_1090),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1168),
.B(n_918),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1208),
.A2(n_977),
.B1(n_1135),
.B2(n_1123),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1172),
.A2(n_994),
.B1(n_1032),
.B2(n_1025),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1169),
.B(n_1088),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1189),
.A2(n_1069),
.B1(n_899),
.B2(n_1032),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1182),
.A2(n_1032),
.B1(n_1052),
.B2(n_1062),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1171),
.B(n_1088),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1192),
.A2(n_1195),
.B1(n_1184),
.B2(n_1196),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1213),
.A2(n_899),
.B1(n_1032),
.B2(n_1041),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1184),
.A2(n_1052),
.B1(n_1062),
.B2(n_1088),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1214),
.A2(n_1062),
.B1(n_1068),
.B2(n_1079),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1184),
.A2(n_646),
.B1(n_652),
.B2(n_586),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1217),
.A2(n_646),
.B1(n_652),
.B2(n_588),
.Y(n_1273)
);

NAND3xp33_ASAP7_75t_L g1274 ( 
.A(n_1209),
.B(n_609),
.C(n_588),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1209),
.A2(n_1194),
.B1(n_1186),
.B2(n_1210),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1210),
.A2(n_638),
.B1(n_651),
.B2(n_588),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1222),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1220),
.A2(n_899),
.B1(n_1079),
.B2(n_1068),
.Y(n_1278)
);

OAI222xp33_ASAP7_75t_L g1279 ( 
.A1(n_1170),
.A2(n_1028),
.B1(n_1051),
.B2(n_644),
.C1(n_653),
.C2(n_544),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1165),
.A2(n_1071),
.B1(n_632),
.B2(n_623),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1165),
.A2(n_623),
.B1(n_609),
.B2(n_632),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1178),
.A2(n_623),
.B1(n_609),
.B2(n_632),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1178),
.A2(n_638),
.B1(n_651),
.B2(n_1071),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1204),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1178),
.B(n_1071),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1226),
.B(n_1200),
.Y(n_1286)
);

NAND3xp33_ASAP7_75t_L g1287 ( 
.A(n_1227),
.B(n_651),
.C(n_638),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1252),
.B(n_1200),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1254),
.B(n_68),
.Y(n_1289)
);

AOI21xp33_ASAP7_75t_L g1290 ( 
.A1(n_1236),
.A2(n_1071),
.B(n_935),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_SL g1291 ( 
.A(n_1279),
.B(n_1215),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1252),
.B(n_1200),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1254),
.B(n_69),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1242),
.B(n_69),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1228),
.B(n_70),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1238),
.B(n_1216),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1228),
.B(n_71),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1268),
.B(n_72),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1277),
.B(n_72),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1277),
.B(n_73),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1224),
.A2(n_73),
.B(n_74),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1235),
.B(n_75),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1248),
.B(n_76),
.Y(n_1303)
);

AND2x2_ASAP7_75t_SL g1304 ( 
.A(n_1246),
.B(n_523),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_L g1305 ( 
.A(n_1256),
.B(n_653),
.C(n_526),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1229),
.B(n_76),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1225),
.A2(n_78),
.B(n_79),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1241),
.A2(n_876),
.B1(n_82),
.B2(n_84),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1230),
.B(n_1275),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1264),
.B(n_81),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1267),
.B(n_82),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1239),
.B(n_84),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1234),
.B(n_85),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1285),
.B(n_1237),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1241),
.A2(n_876),
.B1(n_87),
.B2(n_88),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1231),
.B(n_526),
.C(n_876),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1234),
.B(n_86),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1233),
.A2(n_876),
.B1(n_88),
.B2(n_89),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1240),
.B(n_1261),
.Y(n_1319)
);

NAND3xp33_ASAP7_75t_L g1320 ( 
.A(n_1272),
.B(n_580),
.C(n_563),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1260),
.B(n_90),
.Y(n_1321)
);

OAI22x1_ASAP7_75t_L g1322 ( 
.A1(n_1278),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1258),
.B(n_1265),
.Y(n_1323)
);

NAND3xp33_ASAP7_75t_L g1324 ( 
.A(n_1244),
.B(n_580),
.C(n_563),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1251),
.B(n_546),
.C(n_794),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1245),
.A2(n_1284),
.B(n_1232),
.Y(n_1326)
);

NAND4xp25_ASAP7_75t_SL g1327 ( 
.A(n_1263),
.B(n_92),
.C(n_93),
.D(n_94),
.Y(n_1327)
);

AOI221xp5_ASAP7_75t_L g1328 ( 
.A1(n_1274),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.C(n_99),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1278),
.B(n_98),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1259),
.B(n_546),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1257),
.B(n_100),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1262),
.B(n_105),
.Y(n_1332)
);

NAND3xp33_ASAP7_75t_L g1333 ( 
.A(n_1250),
.B(n_546),
.C(n_110),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1286),
.B(n_1302),
.Y(n_1334)
);

XNOR2xp5_ASAP7_75t_L g1335 ( 
.A(n_1306),
.B(n_1266),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1288),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1292),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1301),
.A2(n_1243),
.B1(n_1247),
.B2(n_1249),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1307),
.A2(n_1276),
.B1(n_1255),
.B2(n_1269),
.Y(n_1339)
);

NOR3xp33_ASAP7_75t_L g1340 ( 
.A(n_1296),
.B(n_1271),
.C(n_1280),
.Y(n_1340)
);

INVx4_ASAP7_75t_SL g1341 ( 
.A(n_1289),
.Y(n_1341)
);

NOR3xp33_ASAP7_75t_L g1342 ( 
.A(n_1296),
.B(n_1269),
.C(n_1270),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1314),
.B(n_1283),
.Y(n_1343)
);

NAND3xp33_ASAP7_75t_L g1344 ( 
.A(n_1329),
.B(n_1282),
.C(n_1281),
.Y(n_1344)
);

OA211x2_ASAP7_75t_L g1345 ( 
.A1(n_1330),
.A2(n_1253),
.B(n_1273),
.C(n_115),
.Y(n_1345)
);

NAND3xp33_ASAP7_75t_L g1346 ( 
.A(n_1308),
.B(n_111),
.C(n_114),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1303),
.B(n_1323),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1289),
.B(n_123),
.Y(n_1348)
);

NAND3xp33_ASAP7_75t_SL g1349 ( 
.A(n_1308),
.B(n_124),
.C(n_130),
.Y(n_1349)
);

NAND4xp75_ASAP7_75t_L g1350 ( 
.A(n_1312),
.B(n_131),
.C(n_132),
.D(n_133),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1294),
.B(n_135),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1309),
.B(n_136),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1293),
.B(n_1295),
.Y(n_1353)
);

AO21x2_ASAP7_75t_L g1354 ( 
.A1(n_1330),
.A2(n_137),
.B(n_139),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1293),
.Y(n_1355)
);

AOI211xp5_ASAP7_75t_L g1356 ( 
.A1(n_1327),
.A2(n_142),
.B(n_145),
.C(n_147),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1295),
.B(n_150),
.Y(n_1357)
);

AND3x1_ASAP7_75t_L g1358 ( 
.A(n_1291),
.B(n_1326),
.C(n_1312),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1297),
.B(n_1298),
.Y(n_1359)
);

AND2x6_ASAP7_75t_L g1360 ( 
.A(n_1313),
.B(n_151),
.Y(n_1360)
);

AO21x2_ASAP7_75t_L g1361 ( 
.A1(n_1317),
.A2(n_153),
.B(n_155),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1299),
.B(n_156),
.Y(n_1362)
);

NAND4xp75_ASAP7_75t_L g1363 ( 
.A(n_1328),
.B(n_157),
.C(n_160),
.D(n_161),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1300),
.B(n_162),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1310),
.B(n_165),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1311),
.B(n_169),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1319),
.B(n_170),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1336),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1337),
.Y(n_1369)
);

XOR2x2_ASAP7_75t_L g1370 ( 
.A(n_1358),
.B(n_1315),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1355),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1353),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1347),
.B(n_1332),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1353),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1341),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1334),
.B(n_1290),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1341),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1360),
.Y(n_1378)
);

NAND4xp75_ASAP7_75t_L g1379 ( 
.A(n_1339),
.B(n_1304),
.C(n_1321),
.D(n_1331),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1359),
.B(n_1343),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1361),
.B(n_1322),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1360),
.B(n_1322),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1361),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1360),
.Y(n_1384)
);

NAND4xp75_ASAP7_75t_SL g1385 ( 
.A(n_1362),
.B(n_1304),
.C(n_1287),
.D(n_1316),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1360),
.B(n_1324),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1335),
.Y(n_1387)
);

XOR2x2_ASAP7_75t_L g1388 ( 
.A(n_1356),
.B(n_1318),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1357),
.Y(n_1389)
);

NAND4xp75_ASAP7_75t_SL g1390 ( 
.A(n_1364),
.B(n_1325),
.C(n_1305),
.D(n_1320),
.Y(n_1390)
);

XNOR2x2_ASAP7_75t_L g1391 ( 
.A(n_1370),
.B(n_1363),
.Y(n_1391)
);

XOR2x2_ASAP7_75t_L g1392 ( 
.A(n_1370),
.B(n_1350),
.Y(n_1392)
);

AO22x2_ASAP7_75t_L g1393 ( 
.A1(n_1383),
.A2(n_1381),
.B1(n_1379),
.B2(n_1382),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1368),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1379),
.A2(n_1339),
.B1(n_1346),
.B2(n_1344),
.Y(n_1395)
);

XOR2x2_ASAP7_75t_L g1396 ( 
.A(n_1387),
.B(n_1349),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1371),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1377),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1374),
.B(n_1342),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1372),
.B(n_1351),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1371),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1374),
.B(n_1352),
.Y(n_1402)
);

INVx5_ASAP7_75t_L g1403 ( 
.A(n_1378),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1375),
.Y(n_1404)
);

INVxp67_ASAP7_75t_SL g1405 ( 
.A(n_1383),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_1378),
.Y(n_1406)
);

OA22x2_ASAP7_75t_L g1407 ( 
.A1(n_1387),
.A2(n_1338),
.B1(n_1348),
.B2(n_1365),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1374),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1381),
.Y(n_1409)
);

AOI22x1_ASAP7_75t_L g1410 ( 
.A1(n_1393),
.A2(n_1406),
.B1(n_1378),
.B2(n_1384),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1394),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1409),
.Y(n_1412)
);

OA22x2_ASAP7_75t_L g1413 ( 
.A1(n_1395),
.A2(n_1384),
.B1(n_1376),
.B2(n_1388),
.Y(n_1413)
);

XNOR2x1_ASAP7_75t_L g1414 ( 
.A(n_1392),
.B(n_1396),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1394),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1409),
.Y(n_1416)
);

XNOR2x1_ASAP7_75t_L g1417 ( 
.A(n_1396),
.B(n_1389),
.Y(n_1417)
);

OA22x2_ASAP7_75t_L g1418 ( 
.A1(n_1395),
.A2(n_1386),
.B1(n_1369),
.B2(n_1338),
.Y(n_1418)
);

AOI22x1_ASAP7_75t_SL g1419 ( 
.A1(n_1406),
.A2(n_1385),
.B1(n_1340),
.B2(n_1390),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1403),
.Y(n_1420)
);

XNOR2x1_ASAP7_75t_SL g1421 ( 
.A(n_1393),
.B(n_1366),
.Y(n_1421)
);

XNOR2x1_ASAP7_75t_L g1422 ( 
.A(n_1393),
.B(n_1380),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1398),
.Y(n_1423)
);

INVx3_ASAP7_75t_SL g1424 ( 
.A(n_1403),
.Y(n_1424)
);

OA22x2_ASAP7_75t_L g1425 ( 
.A1(n_1404),
.A2(n_1367),
.B1(n_1373),
.B2(n_1345),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1412),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1416),
.Y(n_1427)
);

OAI22x1_ASAP7_75t_L g1428 ( 
.A1(n_1410),
.A2(n_1403),
.B1(n_1399),
.B2(n_1408),
.Y(n_1428)
);

NOR2x1_ASAP7_75t_L g1429 ( 
.A(n_1414),
.B(n_1400),
.Y(n_1429)
);

OAI322xp33_ASAP7_75t_L g1430 ( 
.A1(n_1413),
.A2(n_1407),
.A3(n_1391),
.B1(n_1405),
.B2(n_1401),
.C1(n_1397),
.C2(n_1402),
.Y(n_1430)
);

INVx5_ASAP7_75t_SL g1431 ( 
.A(n_1419),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1429),
.Y(n_1432)
);

OAI322xp33_ASAP7_75t_L g1433 ( 
.A1(n_1426),
.A2(n_1413),
.A3(n_1418),
.B1(n_1422),
.B2(n_1417),
.C1(n_1421),
.C2(n_1425),
.Y(n_1433)
);

AOI22x1_ASAP7_75t_L g1434 ( 
.A1(n_1428),
.A2(n_1424),
.B1(n_1420),
.B2(n_1418),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1431),
.A2(n_1418),
.B1(n_1417),
.B2(n_1419),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1435),
.A2(n_1425),
.B1(n_1423),
.B2(n_1427),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1435),
.A2(n_1420),
.B1(n_1430),
.B2(n_1415),
.Y(n_1437)
);

O2A1O1Ixp5_ASAP7_75t_SL g1438 ( 
.A1(n_1432),
.A2(n_1420),
.B(n_1415),
.C(n_1411),
.Y(n_1438)
);

NOR4xp25_ASAP7_75t_L g1439 ( 
.A(n_1433),
.B(n_1411),
.C(n_1333),
.D(n_1354),
.Y(n_1439)
);

NOR2x1_ASAP7_75t_L g1440 ( 
.A(n_1436),
.B(n_1434),
.Y(n_1440)
);

AOI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1439),
.A2(n_171),
.B1(n_172),
.B2(n_179),
.C(n_180),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1437),
.A2(n_181),
.B1(n_183),
.B2(n_185),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1438),
.A2(n_197),
.B1(n_201),
.B2(n_202),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1440),
.A2(n_1442),
.B(n_1441),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1443),
.B(n_204),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1445),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1444),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1446),
.A2(n_221),
.B1(n_223),
.B2(n_225),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1447),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1449),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1448),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1448),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1451),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1452),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1450),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1453),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_1456)
);

AOI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1454),
.A2(n_260),
.B1(n_262),
.B2(n_264),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1456),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1457),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1458),
.A2(n_1455),
.B1(n_270),
.B2(n_275),
.Y(n_1460)
);

OA22x2_ASAP7_75t_L g1461 ( 
.A1(n_1459),
.A2(n_268),
.B1(n_277),
.B2(n_286),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1460),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1461),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1462),
.A2(n_1463),
.B1(n_290),
.B2(n_292),
.C(n_294),
.Y(n_1464)
);

AOI211xp5_ASAP7_75t_L g1465 ( 
.A1(n_1464),
.A2(n_289),
.B(n_298),
.C(n_302),
.Y(n_1465)
);


endmodule