module fake_jpeg_11643_n_374 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_374);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_374;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_47),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_9),
.C(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_56),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_52),
.Y(n_92)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_9),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_58),
.Y(n_95)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_65),
.Y(n_87)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_67),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_18),
.B(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_68),
.Y(n_89)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_26),
.B(n_8),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_31),
.B(n_8),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_36),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_71),
.B(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_20),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_78),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_20),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_79),
.B(n_82),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_24),
.B1(n_38),
.B2(n_30),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_84),
.A2(n_104),
.B1(n_35),
.B2(n_22),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_69),
.B1(n_48),
.B2(n_62),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_100),
.B1(n_24),
.B2(n_38),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_96),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_45),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_36),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_31),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_48),
.A2(n_38),
.B1(n_30),
.B2(n_24),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_64),
.B1(n_67),
.B2(n_30),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_54),
.B(n_28),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_59),
.B(n_28),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_107),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_21),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_21),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_57),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_114),
.B(n_147),
.C(n_95),
.Y(n_169)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_131),
.Y(n_166)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_124),
.B1(n_138),
.B2(n_142),
.Y(n_156)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_24),
.B1(n_38),
.B2(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_82),
.A2(n_28),
.B1(n_34),
.B2(n_26),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_129),
.A2(n_134),
.B1(n_153),
.B2(n_83),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_72),
.A2(n_22),
.B(n_37),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_133),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_34),
.B1(n_22),
.B2(n_43),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_95),
.Y(n_173)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_139),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_18),
.B1(n_41),
.B2(n_34),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_143),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_94),
.B1(n_86),
.B2(n_98),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_87),
.A2(n_35),
.B1(n_41),
.B2(n_53),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_107),
.A2(n_35),
.B1(n_37),
.B2(n_33),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_149),
.B1(n_142),
.B2(n_131),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_91),
.A2(n_37),
.B(n_33),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_148),
.B(n_154),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_81),
.A2(n_33),
.B1(n_49),
.B2(n_39),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_81),
.B(n_0),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_90),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_104),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_163),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_89),
.B1(n_79),
.B2(n_84),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_114),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_164),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_170),
.B1(n_172),
.B2(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_117),
.B(n_89),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_162),
.B(n_180),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_83),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_149),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_173),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_101),
.B1(n_98),
.B2(n_86),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_96),
.C(n_92),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_181),
.C(n_184),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_101),
.B1(n_105),
.B2(n_73),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_174),
.B(n_176),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_118),
.B(n_105),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_113),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_183),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_73),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_98),
.C(n_86),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_80),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_112),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_151),
.A2(n_80),
.B1(n_93),
.B2(n_112),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_115),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_178),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_187),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_200),
.Y(n_231)
);

BUFx12_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_182),
.Y(n_247)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_203),
.B(n_207),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_130),
.B(n_147),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_213),
.B(n_163),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_166),
.A2(n_151),
.B(n_126),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_205),
.B(n_221),
.Y(n_226)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_164),
.A2(n_141),
.B1(n_146),
.B2(n_130),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_212),
.B1(n_218),
.B2(n_158),
.Y(n_228)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_159),
.B(n_188),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_150),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_215),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_211),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_161),
.A2(n_156),
.B1(n_160),
.B2(n_162),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_144),
.B(n_126),
.C(n_114),
.D(n_154),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_155),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_159),
.B(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_182),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_156),
.A2(n_144),
.B1(n_143),
.B2(n_137),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_148),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_171),
.B(n_140),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_223),
.B(n_163),
.Y(n_240)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_136),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_208),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g277 ( 
.A1(n_229),
.A2(n_202),
.B(n_220),
.C(n_219),
.D(n_194),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_184),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_230),
.B(n_234),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_191),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_233),
.B(n_253),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_155),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_216),
.A2(n_155),
.B1(n_163),
.B2(n_159),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_235),
.A2(n_242),
.B(n_252),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_240),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_157),
.B1(n_170),
.B2(n_119),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_243),
.B1(n_246),
.B2(n_199),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_127),
.B1(n_128),
.B2(n_123),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_168),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_230),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_204),
.A2(n_93),
.B1(n_168),
.B2(n_102),
.Y(n_246)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_102),
.B1(n_122),
.B2(n_108),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_251),
.A2(n_207),
.B1(n_215),
.B2(n_196),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_216),
.A2(n_108),
.B1(n_39),
.B2(n_11),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_10),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_214),
.A2(n_0),
.B(n_1),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_214),
.B(n_235),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_197),
.B1(n_192),
.B2(n_193),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_255),
.A2(n_261),
.B1(n_266),
.B2(n_202),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_256),
.A2(n_251),
.B1(n_252),
.B2(n_232),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_257),
.B(n_250),
.Y(n_298)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_206),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_245),
.C(n_225),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_227),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_222),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_264),
.B(n_272),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_236),
.A2(n_202),
.B1(n_213),
.B2(n_206),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_203),
.Y(n_267)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_274),
.B(n_277),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_231),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_276),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_226),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_229),
.A2(n_244),
.B(n_236),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_249),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_275),
.B(n_237),
.Y(n_292)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_279),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_288),
.Y(n_302)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

HAxp5_ASAP7_75t_SL g284 ( 
.A(n_269),
.B(n_226),
.CON(n_284),
.SN(n_284)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_289),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_227),
.Y(n_286)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_286),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_243),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_240),
.B(n_246),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_291),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_267),
.Y(n_291)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_259),
.B1(n_279),
.B2(n_260),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_268),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_244),
.C(n_237),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_257),
.C(n_274),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_299),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_241),
.Y(n_299)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_304),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_282),
.A2(n_294),
.B1(n_256),
.B2(n_297),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_303),
.A2(n_307),
.B1(n_308),
.B2(n_281),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_266),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_305),
.B(n_224),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_282),
.A2(n_259),
.B1(n_258),
.B2(n_275),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_255),
.C(n_278),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_315),
.C(n_287),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_278),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_299),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_238),
.C(n_270),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_261),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_273),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_323),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_329),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_321),
.A2(n_301),
.B(n_315),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_322),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_293),
.B1(n_300),
.B2(n_290),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_310),
.A2(n_283),
.B1(n_286),
.B2(n_287),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_332),
.C(n_314),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_289),
.C(n_284),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_328),
.C(n_304),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_316),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_327),
.A2(n_321),
.B(n_324),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_270),
.C(n_239),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_254),
.Y(n_329)
);

NOR3xp33_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_333),
.C(n_303),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_328),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_307),
.A2(n_285),
.B1(n_198),
.B2(n_200),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_313),
.B(n_285),
.Y(n_333)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_334),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_337),
.B(n_341),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_342),
.Y(n_353)
);

AOI21xp33_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_312),
.B(n_317),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_340),
.A2(n_329),
.B(n_12),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_343),
.A2(n_10),
.B1(n_16),
.B2(n_4),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_306),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_39),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_306),
.C(n_201),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_345),
.B(n_39),
.C(n_12),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_346),
.B(n_347),
.Y(n_358)
);

AO21x1_ASAP7_75t_L g362 ( 
.A1(n_348),
.A2(n_349),
.B(n_14),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_13),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_13),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_354),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_345),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_5),
.C(n_7),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_352),
.A2(n_336),
.B(n_342),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_356),
.A2(n_360),
.B(n_362),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_335),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_335),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_336),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_361),
.B(n_347),
.Y(n_366)
);

FAx1_ASAP7_75t_SL g363 ( 
.A(n_356),
.B(n_354),
.CI(n_349),
.CON(n_363),
.SN(n_363)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_363),
.B(n_366),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_357),
.B(n_358),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_365),
.A2(n_367),
.B(n_14),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_364),
.A2(n_351),
.B(n_14),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_369),
.A2(n_370),
.B(n_366),
.Y(n_371)
);

AOI322xp5_ASAP7_75t_L g372 ( 
.A1(n_371),
.A2(n_1),
.A3(n_3),
.B1(n_15),
.B2(n_16),
.C1(n_368),
.C2(n_365),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_15),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_16),
.B(n_1),
.Y(n_374)
);


endmodule