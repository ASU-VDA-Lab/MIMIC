module fake_jpeg_10636_n_76 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_76);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_76;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_38;
wire n_36;
wire n_74;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx11_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_26),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_5),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_52)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_2),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_51),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_33),
.B(n_36),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_52),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_31),
.B1(n_39),
.B2(n_3),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_54),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_12),
.B(n_13),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_18),
.C(n_20),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_23),
.Y(n_58)
);

FAx1_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_59),
.CI(n_56),
.CON(n_60),
.SN(n_60)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_24),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_61),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_63),
.B(n_68),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_62),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_66),
.B1(n_52),
.B2(n_63),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_60),
.C(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);


endmodule