module fake_jpeg_32102_n_45 (n_3, n_2, n_1, n_0, n_4, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_11),
.B(n_1),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_3),
.C(n_5),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_18),
.A2(n_6),
.B(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_23),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_21),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_3),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_6),
.B(n_12),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_21),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_15),
.A2(n_7),
.B1(n_14),
.B2(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_31),
.B1(n_20),
.B2(n_7),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_18),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_27),
.C(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_14),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_35),
.B1(n_33),
.B2(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_39),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_41),
.C(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);


endmodule