module fake_netlist_6_3219_n_746 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_746);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_746;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_449;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_198;
wire n_300;
wire n_248;
wire n_222;
wire n_517;
wire n_718;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_611;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_692;
wire n_733;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_501;
wire n_531;
wire n_508;
wire n_663;
wire n_361;
wire n_379;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_144),
.Y(n_195)
);

BUFx8_ASAP7_75t_SL g196 ( 
.A(n_88),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_188),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_17),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_13),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_109),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_65),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_95),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_62),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_35),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_133),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_5),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_81),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_51),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_84),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_94),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_137),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_91),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_105),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_18),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_36),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_92),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_70),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_79),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_74),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_178),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_119),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_61),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_130),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_101),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_97),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_26),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_12),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_66),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_82),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_156),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_99),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_167),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_140),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_45),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_42),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_163),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_55),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_154),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_131),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_58),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_1),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_59),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_186),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_34),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_104),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_43),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_33),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_60),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_75),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_63),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_187),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_159),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_190),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_4),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_71),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_191),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_83),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_151),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_57),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_53),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_162),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_153),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_2),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_116),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_164),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_175),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_40),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_155),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_106),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_89),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_112),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_139),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_145),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_113),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_135),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_141),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_189),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_136),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_174),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_80),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_69),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_128),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_123),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_67),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_103),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_138),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_193),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_121),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_192),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_77),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_19),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_98),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_64),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_12),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_24),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_160),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_120),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_117),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_48),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_102),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_184),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_185),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_143),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_168),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_49),
.Y(n_310)
);

BUFx8_ASAP7_75t_SL g311 ( 
.A(n_17),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_50),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_18),
.Y(n_313)
);

INVxp33_ASAP7_75t_R g314 ( 
.A(n_152),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_170),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_100),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_182),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_110),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_68),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_171),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_158),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_166),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_107),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_93),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_126),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_194),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_169),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_22),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_25),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_239),
.B(n_0),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_207),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_300),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_0),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_208),
.Y(n_335)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_197),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_258),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_258),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_196),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_197),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_258),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_220),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_2),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_220),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_220),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_229),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_286),
.B(n_3),
.Y(n_348)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_238),
.Y(n_349)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_244),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_232),
.B(n_242),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_244),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_257),
.B(n_3),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_258),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_317),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_245),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_287),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_217),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_287),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_246),
.Y(n_360)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_287),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_269),
.B(n_5),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_299),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_306),
.B(n_6),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_221),
.B(n_6),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_317),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_254),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_317),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_235),
.B(n_7),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_308),
.B(n_7),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_248),
.B(n_8),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_318),
.B(n_8),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_263),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_263),
.B(n_9),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_259),
.B(n_9),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_288),
.Y(n_378)
);

BUFx8_ASAP7_75t_SL g379 ( 
.A(n_199),
.Y(n_379)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_298),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_298),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_313),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_201),
.B(n_10),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_305),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_320),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_11),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

INVx5_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_204),
.B(n_11),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_212),
.B(n_14),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_230),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_213),
.B(n_14),
.Y(n_393)
);

BUFx8_ASAP7_75t_SL g394 ( 
.A(n_225),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_214),
.B(n_15),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_216),
.B(n_16),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_222),
.B(n_19),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_271),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_262),
.B(n_20),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_227),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_233),
.B(n_20),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_304),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_304),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_316),
.B(n_21),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_240),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_241),
.Y(n_407)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_314),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_247),
.B(n_22),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_268),
.Y(n_410)
);

BUFx10_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_343),
.A2(n_226),
.B1(n_236),
.B2(n_228),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_L g414 ( 
.A1(n_376),
.A2(n_200),
.B1(n_328),
.B2(n_296),
.Y(n_414)
);

AO22x2_ASAP7_75t_L g415 ( 
.A1(n_405),
.A2(n_253),
.B1(n_260),
.B2(n_252),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_330),
.A2(n_275),
.B1(n_291),
.B2(n_272),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_365),
.A2(n_372),
.B1(n_400),
.B2(n_370),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_331),
.A2(n_302),
.B1(n_307),
.B2(n_301),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_394),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

AO22x2_ASAP7_75t_L g421 ( 
.A1(n_362),
.A2(n_266),
.B1(n_270),
.B2(n_265),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_333),
.A2(n_315),
.B1(n_198),
.B2(n_202),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

AO22x2_ASAP7_75t_L g424 ( 
.A1(n_362),
.A2(n_279),
.B1(n_282),
.B2(n_277),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_195),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_203),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_351),
.B(n_353),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_340),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_346),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_L g430 ( 
.A1(n_356),
.A2(n_290),
.B1(n_292),
.B2(n_289),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_367),
.A2(n_206),
.B1(n_209),
.B2(n_205),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_399),
.B(n_210),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_342),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_408),
.A2(n_349),
.B1(n_374),
.B2(n_358),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_351),
.B(n_293),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_403),
.B(n_211),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_392),
.A2(n_327),
.B1(n_215),
.B2(n_218),
.Y(n_438)
);

AO22x2_ASAP7_75t_L g439 ( 
.A1(n_377),
.A2(n_326),
.B1(n_325),
.B2(n_324),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_352),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_371),
.A2(n_323),
.B1(n_322),
.B2(n_321),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_352),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_SL g443 ( 
.A(n_373),
.B(n_219),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_364),
.A2(n_267),
.B1(n_223),
.B2(n_224),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_342),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_404),
.B(n_23),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_357),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_349),
.A2(n_319),
.B1(n_310),
.B2(n_309),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_404),
.B(n_231),
.Y(n_452)
);

NAND3x1_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_24),
.C(n_25),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_359),
.Y(n_454)
);

OA22x2_ASAP7_75t_L g455 ( 
.A1(n_335),
.A2(n_297),
.B1(n_295),
.B2(n_294),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_410),
.B(n_234),
.Y(n_456)
);

OAI22xp33_ASAP7_75t_L g457 ( 
.A1(n_383),
.A2(n_398),
.B1(n_393),
.B2(n_397),
.Y(n_457)
);

AO22x2_ASAP7_75t_L g458 ( 
.A1(n_390),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_345),
.A2(n_285),
.B1(n_284),
.B2(n_283),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_368),
.Y(n_460)
);

OAI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_391),
.A2(n_281),
.B1(n_280),
.B2(n_278),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_406),
.B(n_336),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_387),
.A2(n_276),
.B1(n_274),
.B2(n_273),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_395),
.A2(n_249),
.B1(n_261),
.B2(n_256),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_336),
.B(n_237),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_402),
.A2(n_264),
.B1(n_255),
.B2(n_251),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_378),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_332),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_427),
.B(n_407),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_457),
.B(n_395),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_428),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_418),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_433),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_434),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_445),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_451),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_460),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_417),
.B(n_375),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_413),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_334),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_429),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_447),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_440),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_442),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_449),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g487 ( 
.A(n_416),
.B(n_336),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_467),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_447),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_454),
.Y(n_492)
);

OR2x6_ASAP7_75t_L g493 ( 
.A(n_458),
.B(n_348),
.Y(n_493)
);

BUFx6f_ASAP7_75t_SL g494 ( 
.A(n_411),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_436),
.B(n_375),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_420),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_420),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_425),
.B(n_380),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_436),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_414),
.B(n_380),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_455),
.A2(n_338),
.B(n_337),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_465),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_446),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_443),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_421),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_426),
.Y(n_507)
);

XNOR2x1_ASAP7_75t_L g508 ( 
.A(n_458),
.B(n_379),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_412),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_424),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_439),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_464),
.A2(n_463),
.B(n_441),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_422),
.B(n_401),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_415),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_415),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_437),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_435),
.B(n_243),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_438),
.B(n_347),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_450),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_432),
.B(n_347),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_430),
.Y(n_522)
);

INVxp33_ASAP7_75t_L g523 ( 
.A(n_459),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_456),
.Y(n_524)
);

XNOR2x2_ASAP7_75t_L g525 ( 
.A(n_453),
.B(n_360),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_466),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_444),
.B(n_341),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_431),
.B(n_363),
.Y(n_528)
);

BUFx5_ASAP7_75t_L g529 ( 
.A(n_411),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_507),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_502),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_512),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_472),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_469),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_498),
.B(n_461),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_468),
.B(n_419),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_483),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_501),
.A2(n_355),
.B(n_354),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

AND2x2_ASAP7_75t_SL g540 ( 
.A(n_510),
.B(n_366),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_499),
.B(n_382),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_524),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_479),
.B(n_401),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_521),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_470),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_515),
.B(n_516),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_481),
.Y(n_547)
);

AND2x2_ASAP7_75t_SL g548 ( 
.A(n_526),
.B(n_369),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_475),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_505),
.B(n_388),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_491),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_476),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_519),
.B(n_401),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_481),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_506),
.B(n_396),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_494),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_477),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_503),
.B(n_378),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_478),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_489),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_514),
.B(n_527),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_480),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_521),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_482),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_484),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_514),
.B(n_517),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_485),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_486),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_471),
.B(n_250),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_488),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_500),
.B(n_28),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_490),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_529),
.B(n_381),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_501),
.B(n_32),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_495),
.B(n_389),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_528),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_509),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_500),
.B(n_384),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_496),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_497),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_513),
.A2(n_389),
.B(n_386),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_504),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_513),
.B(n_350),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_511),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_544),
.B(n_522),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_538),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_538),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_533),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_532),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_585),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_544),
.B(n_487),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_585),
.Y(n_593)
);

INVx6_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_533),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_547),
.B(n_543),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_539),
.Y(n_597)
);

BUFx12f_ASAP7_75t_L g598 ( 
.A(n_556),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_563),
.B(n_520),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_554),
.B(n_493),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_539),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_561),
.B(n_523),
.Y(n_602)
);

OR2x6_ASAP7_75t_L g603 ( 
.A(n_563),
.B(n_493),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_553),
.B(n_548),
.Y(n_604)
);

NAND2x1p5_ASAP7_75t_L g605 ( 
.A(n_563),
.B(n_574),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_540),
.B(n_473),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_566),
.B(n_518),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_530),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_579),
.B(n_385),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_537),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_531),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_534),
.B(n_525),
.Y(n_612)
);

NOR2x1_ASAP7_75t_L g613 ( 
.A(n_536),
.B(n_508),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_531),
.B(n_385),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_589),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_596),
.B(n_571),
.Y(n_616)
);

BUFx12f_ASAP7_75t_L g617 ( 
.A(n_598),
.Y(n_617)
);

BUFx4f_ASAP7_75t_SL g618 ( 
.A(n_598),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_605),
.B(n_574),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_599),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_589),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_608),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_595),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_586),
.B(n_577),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_591),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_603),
.B(n_577),
.Y(n_626)
);

BUFx12f_ASAP7_75t_L g627 ( 
.A(n_612),
.Y(n_627)
);

CKINVDCx11_ASAP7_75t_R g628 ( 
.A(n_603),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_595),
.Y(n_629)
);

BUFx12f_ASAP7_75t_L g630 ( 
.A(n_599),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_599),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_586),
.Y(n_632)
);

NAND2x1_ASAP7_75t_L g633 ( 
.A(n_611),
.B(n_537),
.Y(n_633)
);

BUFx12f_ASAP7_75t_L g634 ( 
.A(n_617),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_616),
.A2(n_602),
.B1(n_607),
.B2(n_604),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_617),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_615),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_625),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_621),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_621),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_L g641 ( 
.A1(n_627),
.A2(n_606),
.B1(n_605),
.B2(n_600),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_623),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_623),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_618),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_629),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_632),
.A2(n_584),
.B1(n_582),
.B2(n_531),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_620),
.B(n_590),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_624),
.A2(n_540),
.B1(n_613),
.B2(n_630),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_629),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_635),
.A2(n_584),
.B1(n_632),
.B2(n_628),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_638),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_641),
.A2(n_624),
.B1(n_631),
.B2(n_583),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_641),
.A2(n_535),
.B1(n_592),
.B2(n_569),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_648),
.A2(n_626),
.B1(n_619),
.B2(n_541),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_639),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_647),
.A2(n_541),
.B1(n_593),
.B2(n_609),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_640),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_646),
.A2(n_542),
.B1(n_564),
.B2(n_570),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_636),
.A2(n_542),
.B1(n_594),
.B2(n_558),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_634),
.A2(n_565),
.B1(n_568),
.B2(n_567),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_642),
.A2(n_562),
.B1(n_575),
.B2(n_552),
.Y(n_661)
);

OAI222xp33_ASAP7_75t_L g662 ( 
.A1(n_645),
.A2(n_614),
.B1(n_580),
.B2(n_560),
.C1(n_572),
.C2(n_557),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_649),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_637),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_644),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_637),
.A2(n_557),
.B1(n_559),
.B2(n_545),
.Y(n_666)
);

OAI222xp33_ASAP7_75t_L g667 ( 
.A1(n_643),
.A2(n_572),
.B1(n_560),
.B2(n_559),
.C1(n_549),
.C2(n_545),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_650),
.A2(n_653),
.B1(n_652),
.B2(n_654),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_656),
.A2(n_550),
.B1(n_555),
.B2(n_573),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_655),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_660),
.A2(n_622),
.B1(n_551),
.B2(n_581),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_667),
.A2(n_633),
.B(n_588),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_657),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_663),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_664),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_661),
.A2(n_555),
.B1(n_550),
.B2(n_601),
.Y(n_676)
);

AOI222xp33_ASAP7_75t_L g677 ( 
.A1(n_662),
.A2(n_578),
.B1(n_546),
.B2(n_597),
.C1(n_601),
.C2(n_29),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_665),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_666),
.B(n_658),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_666),
.A2(n_546),
.B1(n_576),
.B2(n_610),
.Y(n_680)
);

OA21x2_ASAP7_75t_L g681 ( 
.A1(n_653),
.A2(n_587),
.B(n_588),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_651),
.Y(n_682)
);

OAI22x1_ASAP7_75t_L g683 ( 
.A1(n_659),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_683)
);

OAI221xp5_ASAP7_75t_SL g684 ( 
.A1(n_668),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.C(n_41),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_674),
.B(n_44),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_682),
.B(n_46),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_682),
.B(n_47),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_670),
.B(n_52),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_675),
.B(n_54),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_673),
.B(n_56),
.Y(n_690)
);

AOI21xp33_ASAP7_75t_L g691 ( 
.A1(n_677),
.A2(n_72),
.B(n_73),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_679),
.B(n_76),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_683),
.B(n_78),
.Y(n_693)
);

OA21x2_ASAP7_75t_L g694 ( 
.A1(n_672),
.A2(n_85),
.B(n_86),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_678),
.B(n_87),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_686),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_687),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_690),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_694),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_695),
.B(n_681),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_691),
.A2(n_669),
.B1(n_681),
.B2(n_671),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_685),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_684),
.B(n_676),
.C(n_680),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_692),
.B(n_90),
.Y(n_704)
);

AND2x4_ASAP7_75t_SL g705 ( 
.A(n_688),
.B(n_96),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_689),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_696),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_697),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_700),
.B(n_693),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_698),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_702),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_699),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_706),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_704),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_713),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_707),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_710),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_711),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_708),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_L g720 ( 
.A1(n_714),
.A2(n_703),
.B1(n_701),
.B2(n_705),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_712),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_709),
.Y(n_722)
);

AO22x1_ASAP7_75t_L g723 ( 
.A1(n_721),
.A2(n_361),
.B1(n_111),
.B2(n_114),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_722),
.B(n_108),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_720),
.A2(n_115),
.B1(n_118),
.B2(n_122),
.Y(n_725)
);

OAI22x1_ASAP7_75t_L g726 ( 
.A1(n_718),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_715),
.A2(n_129),
.B1(n_132),
.B2(n_134),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_716),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_717),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_728),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_729),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_731),
.Y(n_732)
);

AND4x1_ASAP7_75t_L g733 ( 
.A(n_730),
.B(n_725),
.C(n_727),
.D(n_724),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_732),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_734),
.A2(n_733),
.B1(n_726),
.B2(n_719),
.Y(n_735)
);

NOR2x1_ASAP7_75t_L g736 ( 
.A(n_735),
.B(n_723),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_736),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_737),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_738),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_739),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_740),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_741),
.Y(n_742)
);

AO22x2_ASAP7_75t_L g743 ( 
.A1(n_742),
.A2(n_740),
.B1(n_149),
.B2(n_150),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_743),
.Y(n_744)
);

AOI221xp5_ASAP7_75t_L g745 ( 
.A1(n_744),
.A2(n_157),
.B1(n_161),
.B2(n_165),
.C(n_173),
.Y(n_745)
);

AOI211xp5_ASAP7_75t_L g746 ( 
.A1(n_745),
.A2(n_177),
.B(n_180),
.C(n_181),
.Y(n_746)
);


endmodule