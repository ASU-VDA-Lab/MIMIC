module real_jpeg_22184_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_335, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_335;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_0),
.A2(n_70),
.B1(n_71),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_0),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_0),
.A2(n_47),
.B1(n_49),
.B2(n_122),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_0),
.A2(n_36),
.B1(n_37),
.B2(n_122),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_122),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_1),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_1),
.A2(n_30),
.B1(n_70),
.B2(n_71),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_1),
.A2(n_30),
.B1(n_47),
.B2(n_49),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_2),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_2),
.A2(n_52),
.B1(n_70),
.B2(n_71),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_47),
.B1(n_49),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_3),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_70),
.B1(n_71),
.B2(n_117),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_117),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_117),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_4),
.A2(n_39),
.B1(n_70),
.B2(n_71),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_4),
.A2(n_39),
.B1(n_47),
.B2(n_49),
.Y(n_282)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_6),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_6),
.A2(n_70),
.B1(n_71),
.B2(n_84),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_6),
.A2(n_47),
.B1(n_49),
.B2(n_84),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_84),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_7),
.A2(n_49),
.B(n_66),
.C(n_102),
.D(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_7),
.B(n_49),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_7),
.B(n_46),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_7),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_7),
.A2(n_123),
.B(n_125),
.Y(n_147)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_7),
.A2(n_36),
.B(n_43),
.C(n_162),
.D(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_7),
.B(n_36),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_7),
.B(n_40),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_7),
.A2(n_37),
.B(n_202),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_141),
.Y(n_219)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_10),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_10),
.A2(n_63),
.B1(n_70),
.B2(n_71),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_10),
.A2(n_47),
.B1(n_49),
.B2(n_63),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_63),
.Y(n_275)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_12),
.A2(n_47),
.B1(n_49),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_12),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_12),
.A2(n_70),
.B1(n_71),
.B2(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_105),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_105),
.Y(n_222)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_14),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_92),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_90),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_76),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_53),
.B1(n_54),
.B2(n_75),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_22),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_41),
.B2(n_42),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_38),
.B2(n_40),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_26),
.A2(n_32),
.B1(n_35),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_33),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_28),
.A2(n_33),
.B(n_141),
.C(n_201),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_31),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_31),
.B(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_32),
.A2(n_35),
.B1(n_62),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_32),
.A2(n_35),
.B1(n_230),
.B2(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_32),
.A2(n_221),
.B(n_259),
.Y(n_277)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_33),
.Y(n_202)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_35),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_35),
.A2(n_83),
.B(n_231),
.Y(n_301)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_44),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_40),
.B(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_50),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_43),
.B(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_43),
.A2(n_46),
.B1(n_256),
.B2(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_43),
.A2(n_46),
.B1(n_89),
.B2(n_275),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_45),
.Y(n_170)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_47),
.B(n_48),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_49),
.A2(n_162),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.C(n_64),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_56),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_57),
.A2(n_59),
.B1(n_181),
.B2(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_57),
.A2(n_216),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_59),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_59),
.A2(n_181),
.B(n_182),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_59),
.A2(n_182),
.B(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_61),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_64),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_73),
.B(n_74),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_65),
.A2(n_73),
.B1(n_116),
.B2(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_65),
.A2(n_160),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_65),
.A2(n_73),
.B1(n_213),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_65),
.A2(n_73),
.B1(n_241),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_65),
.A2(n_73),
.B1(n_250),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_66),
.B(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_66),
.A2(n_69),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

CKINVDCx9p33_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_71),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_70),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NAND2x1_ASAP7_75t_SL g123 ( 
.A(n_70),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_71),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_116),
.B(n_118),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_73),
.B(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_73),
.A2(n_118),
.B(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_74),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.C(n_85),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_320),
.Y(n_326)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.C(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_82),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_82),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_85),
.B(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI321xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_317),
.A3(n_327),
.B1(n_332),
.B2(n_333),
.C(n_335),
.Y(n_92)
);

AOI321xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_267),
.A3(n_305),
.B1(n_311),
.B2(n_316),
.C(n_336),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_224),
.C(n_263),
.Y(n_94)
);

AOI21x1_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_194),
.B(n_223),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_175),
.B(n_193),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_154),
.B(n_174),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_129),
.B(n_153),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_100),
.B(n_110),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_106),
.B1(n_107),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_103),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_115),
.C(n_120),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_123),
.B(n_125),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_127),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_123),
.A2(n_124),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_123),
.A2(n_150),
.B1(n_206),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_123),
.A2(n_143),
.B1(n_239),
.B2(n_248),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_123),
.A2(n_124),
.B(n_248),
.Y(n_280)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_128),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_145),
.B(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_128),
.A2(n_134),
.B1(n_172),
.B2(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_138),
.B(n_152),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_131),
.B(n_136),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_146),
.B(n_151),
.Y(n_138)
);

NOR2x1_ASAP7_75t_R g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_142),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_155),
.B(n_156),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_167),
.B2(n_173),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_161),
.B1(n_165),
.B2(n_166),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_166),
.C(n_173),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_163),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_167),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_177),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_189),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_190),
.C(n_191),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_184),
.B2(n_188),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_185),
.C(n_186),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_196),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_210),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_198),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_198),
.B(n_209),
.C(n_210),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_204),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_217),
.C(n_218),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g312 ( 
.A1(n_225),
.A2(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_243),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_226),
.B(n_243),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_237),
.C(n_242),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_236),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_232),
.B1(n_233),
.B2(n_235),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_242),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_240),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_261),
.B2(n_262),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_251),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_246),
.B(n_251),
.C(n_262),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_249),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_257),
.C(n_260),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_257),
.B1(n_258),
.B2(n_260),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_254),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_261),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_265),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_285),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_268),
.B(n_285),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_278),
.C(n_284),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_269),
.A2(n_270),
.B1(n_278),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_274),
.C(n_276),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_283),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_280),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_279),
.A2(n_297),
.B(n_301),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_281),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_281),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_282),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_303),
.B2(n_304),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_295),
.B2(n_296),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_296),
.C(n_304),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_293),
.B(n_294),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_293),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_294),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_294),
.A2(n_319),
.B1(n_323),
.B2(n_331),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_302),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_303),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_306),
.A2(n_312),
.B(n_315),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_308),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_325),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_325),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.C(n_324),
.Y(n_318)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);


endmodule