module fake_jpeg_16797_n_46 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_46);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_17;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx12_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_8),
.B(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_3),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_29),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_32),
.B(n_33),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_19),
.A2(n_16),
.B1(n_18),
.B2(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_27),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_21),
.A2(n_27),
.B1(n_20),
.B2(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_22),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_31),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_36),
.B1(n_34),
.B2(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_35),
.C(n_43),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_22),
.B(n_36),
.Y(n_46)
);


endmodule