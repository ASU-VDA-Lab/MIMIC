module real_jpeg_28685_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_0),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_0),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_1),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_2),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_107),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_107),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_2),
.A2(n_48),
.B1(n_50),
.B2(n_107),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_3),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_SL g118 ( 
.A1(n_3),
.A2(n_28),
.B(n_32),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_117),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_30),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_3),
.A2(n_54),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_3),
.B(n_54),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_3),
.B(n_66),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_3),
.A2(n_85),
.B1(n_242),
.B2(n_246),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_3),
.A2(n_31),
.B(n_258),
.Y(n_257)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_5),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_113),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_113),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_113),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_6),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_6),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_36),
.B1(n_54),
.B2(n_55),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_8),
.A2(n_36),
.B1(n_48),
.B2(n_50),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_10),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_97),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_97),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_10),
.A2(n_48),
.B1(n_50),
.B2(n_97),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_11),
.A2(n_50),
.A3(n_54),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_12),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_104),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_12),
.A2(n_48),
.B1(n_50),
.B2(n_104),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_104),
.Y(n_262)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_14),
.B(n_31),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_14),
.A2(n_54),
.B1(n_55),
.B2(n_61),
.Y(n_63)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_14),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_15),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_15),
.A2(n_26),
.B1(n_48),
.B2(n_50),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_15),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_138)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_16),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_17),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g179 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_102),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_17),
.A2(n_54),
.B1(n_55),
.B2(n_102),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_17),
.A2(n_48),
.B1(n_50),
.B2(n_102),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_76),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_21),
.B(n_37),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_23),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_25),
.A2(n_34),
.B(n_117),
.C(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_27),
.A2(n_30),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_27),
.A2(n_30),
.B1(n_103),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_27),
.A2(n_30),
.B1(n_112),
.B2(n_185),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_31),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

OAI32xp33_ASAP7_75t_L g266 ( 
.A1(n_31),
.A2(n_55),
.A3(n_259),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_32),
.B(n_117),
.Y(n_259)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_67),
.C(n_69),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_38),
.A2(n_39),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_57),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_40),
.B(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_42),
.A2(n_71),
.B1(n_73),
.B2(n_165),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_46),
.A2(n_308),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_46),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_46),
.A2(n_57),
.B1(n_311),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_52),
.B(n_56),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_47),
.A2(n_52),
.B1(n_95),
.B2(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_47),
.A2(n_52),
.B1(n_98),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_47),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_47),
.A2(n_52),
.B1(n_56),
.B2(n_138),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_47),
.A2(n_52),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_47),
.A2(n_52),
.B1(n_216),
.B2(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_47),
.B(n_117),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_47),
.A2(n_52),
.B1(n_183),
.B2(n_286),
.Y(n_285)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_48),
.B(n_51),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_48),
.B(n_248),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_52),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_54),
.B(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_57),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_58),
.A2(n_66),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_58),
.A2(n_66),
.B1(n_108),
.B2(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_58),
.A2(n_66),
.B1(n_179),
.B2(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_58),
.A2(n_64),
.B1(n_66),
.B2(n_309),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_63),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_59),
.A2(n_63),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_59),
.A2(n_63),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_59),
.A2(n_63),
.B1(n_123),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_59),
.A2(n_63),
.B1(n_191),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_67),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_73),
.B1(n_111),
.B2(n_114),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_71),
.A2(n_73),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_326),
.B(n_332),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_302),
.A3(n_321),
.B1(n_324),
.B2(n_325),
.C(n_336),
.Y(n_77)
);

AOI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_149),
.A3(n_171),
.B1(n_296),
.B2(n_301),
.C(n_337),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_80),
.A2(n_297),
.B(n_300),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_130),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_81),
.B(n_130),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_109),
.C(n_125),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_82),
.B(n_125),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_99),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_83),
.B(n_100),
.C(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_94),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_84),
.B(n_94),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B1(n_90),
.B2(n_93),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_92),
.B1(n_93),
.B2(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_85),
.A2(n_90),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_85),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_85),
.A2(n_92),
.B1(n_236),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_85),
.A2(n_230),
.B1(n_231),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_89),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_86),
.A2(n_91),
.B1(n_120),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_86),
.A2(n_91),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g231 ( 
.A(n_91),
.Y(n_231)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_96),
.A2(n_136),
.B1(n_139),
.B2(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_109),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.C(n_122),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_110),
.B(n_122),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_115),
.B(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_116),
.B(n_119),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_117),
.B(n_246),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_128),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_129),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_148),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_142),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_142),
.C(n_148),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_140),
.B2(n_141),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_133),
.B(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_139),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_136),
.A2(n_139),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_141),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_140),
.A2(n_163),
.B(n_166),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_142),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_145),
.CI(n_147),
.CON(n_142),
.SN(n_142)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_145),
.C(n_147),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_150),
.B(n_151),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_169),
.B2(n_170),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_154),
.B(n_160),
.C(n_170),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_158),
.B(n_159),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_158),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_157),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_159),
.B(n_304),
.C(n_313),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_159),
.B(n_304),
.CI(n_313),
.CON(n_323),
.SN(n_323)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_169),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_201),
.C(n_206),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_195),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_173),
.B(n_195),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_186),
.C(n_187),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_174),
.B(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_184),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_181),
.C(n_184),
.Y(n_198)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_186),
.Y(n_294)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_189),
.B(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_192),
.B(n_194),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_193),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_198),
.C(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_202),
.A2(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_203),
.B(n_204),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_290),
.B(n_295),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_276),
.B(n_289),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_252),
.B(n_275),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_232),
.B(n_251),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_221),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_211),
.B(n_221),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_212),
.A2(n_213),
.B1(n_217),
.B2(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_226),
.C(n_228),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_227),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_229),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_239),
.B(n_250),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_244),
.B(n_249),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_253),
.B(n_254),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_265),
.B1(n_273),
.B2(n_274),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_255)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_264),
.C(n_274),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_262),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_265),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_271),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_271),
.Y(n_284)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_285),
.C(n_287),
.Y(n_291)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_288),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_314),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_314),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_312),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_306),
.B1(n_316),
.B2(n_319),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_308),
.C(n_311),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_319),
.C(n_320),
.Y(n_327)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_308),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_322),
.B(n_323),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_323),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule