module fake_netlist_6_2244_n_1337 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_321, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1337);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_321;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1337;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_680;
wire n_367;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g322 ( 
.A(n_179),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_127),
.B(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_5),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_30),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_185),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_238),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_272),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_319),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_226),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_198),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_98),
.B(n_312),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_24),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_93),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_154),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_155),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_112),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_135),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_98),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_53),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_303),
.Y(n_343)
);

BUFx2_ASAP7_75t_SL g344 ( 
.A(n_148),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_174),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_39),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_186),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_294),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_206),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_146),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_293),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_53),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_291),
.B(n_181),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_247),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_306),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_229),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_32),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_214),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_122),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_210),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_212),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_64),
.Y(n_363)
);

BUFx10_ASAP7_75t_L g364 ( 
.A(n_152),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_59),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_263),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_269),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_208),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_72),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_314),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_248),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_167),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_137),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_211),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_76),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_136),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_156),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_239),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_255),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_157),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_281),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_38),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_5),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_250),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_182),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_233),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_217),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_292),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_83),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_45),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_313),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_121),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_188),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_320),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_126),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_237),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_130),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_166),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_91),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_61),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_205),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_191),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_7),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_59),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_266),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_80),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_66),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_254),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_252),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_289),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_249),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_270),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_227),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_257),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_241),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_140),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_196),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_27),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_298),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_159),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_207),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_284),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_290),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_244),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_216),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_128),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_299),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_277),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_151),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_82),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_271),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_39),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_253),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_4),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_50),
.B(n_93),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_163),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_268),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_168),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_9),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_118),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_117),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_41),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_51),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_176),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_224),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_192),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_288),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_22),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_28),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_8),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_22),
.B(n_195),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_103),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_51),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_162),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_190),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_180),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_318),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_321),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_199),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_258),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_84),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_131),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_18),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_260),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_70),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_315),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_138),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_134),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_240),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_309),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_144),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_45),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_287),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_139),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_296),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_275),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_125),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_302),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_209),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_261),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_183),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_274),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_194),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_251),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_19),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_109),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_259),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_200),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_29),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_1),
.Y(n_491)
);

INVxp33_ASAP7_75t_SL g492 ( 
.A(n_112),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_243),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_365),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_380),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_380),
.B(n_0),
.Y(n_496)
);

BUFx12f_ASAP7_75t_L g497 ( 
.A(n_362),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_365),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_391),
.B(n_0),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_369),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_391),
.B(n_1),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_422),
.Y(n_502)
);

CKINVDCx6p67_ASAP7_75t_R g503 ( 
.A(n_431),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_362),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_369),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_368),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_360),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_368),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_384),
.B(n_2),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_360),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_360),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_360),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_368),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_368),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_341),
.B(n_2),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_L g516 ( 
.A(n_334),
.B(n_3),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_422),
.Y(n_517)
);

OA21x2_ASAP7_75t_L g518 ( 
.A1(n_415),
.A2(n_3),
.B(n_4),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_341),
.B(n_6),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_466),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_390),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_445),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_325),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_338),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_423),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_423),
.B(n_6),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_428),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_428),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_346),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_445),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_466),
.B(n_7),
.Y(n_531)
);

OA21x2_ASAP7_75t_L g532 ( 
.A1(n_415),
.A2(n_8),
.B(n_9),
.Y(n_532)
);

CKINVDCx6p67_ASAP7_75t_R g533 ( 
.A(n_412),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_360),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_340),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_448),
.B(n_10),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_456),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_456),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_360),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_340),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_489),
.B(n_10),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_489),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_364),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_364),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_348),
.A2(n_115),
.B(n_114),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_353),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_363),
.Y(n_547)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_488),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_363),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_416),
.A2(n_11),
.B(n_12),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_355),
.B(n_455),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_404),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_386),
.A2(n_119),
.B(n_116),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_382),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_335),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_355),
.B(n_13),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_488),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_404),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_481),
.B(n_14),
.Y(n_559)
);

CKINVDCx6p67_ASAP7_75t_R g560 ( 
.A(n_413),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_486),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_326),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_486),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_435),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_444),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_450),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_327),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_449),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_401),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_372),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_481),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_470),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_490),
.A2(n_25),
.B1(n_20),
.B2(n_21),
.Y(n_573)
);

OAI22x1_ASAP7_75t_R g574 ( 
.A1(n_375),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_469),
.B(n_455),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_407),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_416),
.B(n_120),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_517),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_506),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_506),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_506),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_508),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_508),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_SL g584 ( 
.A(n_515),
.B(n_484),
.Y(n_584)
);

AOI21x1_ASAP7_75t_L g585 ( 
.A1(n_507),
.A2(n_430),
.B(n_417),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_508),
.Y(n_586)
);

INVxp33_ASAP7_75t_SL g587 ( 
.A(n_520),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_551),
.B(n_484),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_513),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_559),
.B(n_417),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_572),
.B(n_430),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_575),
.B(n_418),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_513),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_514),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_514),
.Y(n_595)
);

CKINVDCx6p67_ASAP7_75t_R g596 ( 
.A(n_533),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_517),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_547),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_551),
.A2(n_519),
.B1(n_531),
.B2(n_509),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_549),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_522),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_510),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_549),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_558),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_509),
.A2(n_492),
.B1(n_440),
.B2(n_453),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g606 ( 
.A1(n_511),
.A2(n_459),
.B(n_442),
.Y(n_606)
);

INVxp67_ASAP7_75t_SL g607 ( 
.A(n_525),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_558),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_520),
.B(n_452),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_515),
.A2(n_454),
.B1(n_462),
.B2(n_433),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_548),
.Y(n_612)
);

INVxp33_ASAP7_75t_L g613 ( 
.A(n_521),
.Y(n_613)
);

INVxp33_ASAP7_75t_L g614 ( 
.A(n_535),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_568),
.Y(n_615)
);

NOR2x1p5_ASAP7_75t_L g616 ( 
.A(n_497),
.B(n_357),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_568),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_543),
.B(n_333),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_569),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_512),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_539),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_569),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_548),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_543),
.B(n_333),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_525),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_534),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_543),
.B(n_388),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_543),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_572),
.B(n_442),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_582),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_580),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_599),
.B(n_544),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_605),
.A2(n_556),
.B1(n_571),
.B2(n_536),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_588),
.B(n_541),
.C(n_536),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_579),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_581),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_580),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_592),
.Y(n_638)
);

BUFx5_ASAP7_75t_L g639 ( 
.A(n_590),
.Y(n_639)
);

OAI221xp5_ASAP7_75t_L g640 ( 
.A1(n_611),
.A2(n_541),
.B1(n_556),
.B2(n_554),
.C(n_516),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_607),
.B(n_572),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_581),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_580),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_614),
.B(n_544),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_591),
.A2(n_357),
.B(n_496),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_583),
.Y(n_646)
);

BUFx12f_ASAP7_75t_L g647 ( 
.A(n_616),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_613),
.B(n_544),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_612),
.B(n_562),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_L g650 ( 
.A(n_584),
.B(n_573),
.C(n_564),
.Y(n_650)
);

BUFx4f_ASAP7_75t_L g651 ( 
.A(n_596),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_587),
.B(n_504),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_610),
.A2(n_560),
.B1(n_358),
.B2(n_567),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g654 ( 
.A(n_601),
.B(n_530),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_586),
.Y(n_655)
);

OR2x6_ASAP7_75t_L g656 ( 
.A(n_612),
.B(n_573),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_623),
.B(n_567),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_590),
.A2(n_499),
.B1(n_501),
.B2(n_496),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_587),
.A2(n_570),
.B1(n_499),
.B2(n_526),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_586),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_601),
.B(n_530),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_593),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_SL g663 ( 
.A(n_623),
.B(n_328),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_628),
.B(n_570),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_627),
.B(n_527),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_618),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_624),
.B(n_503),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_578),
.B(n_527),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_594),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_594),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_597),
.B(n_548),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_629),
.A2(n_526),
.B(n_501),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_595),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_580),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_625),
.A2(n_436),
.B1(n_377),
.B2(n_392),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_615),
.B(n_495),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_620),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_621),
.A2(n_545),
.B(n_553),
.C(n_516),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_580),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_590),
.A2(n_565),
.B1(n_555),
.B2(n_406),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_621),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_596),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_602),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_619),
.B(n_495),
.Y(n_684)
);

AO221x1_ASAP7_75t_L g685 ( 
.A1(n_602),
.A2(n_350),
.B1(n_330),
.B2(n_329),
.C(n_323),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_617),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_619),
.B(n_502),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_589),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_617),
.B(n_528),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_589),
.Y(n_690)
);

O2A1O1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_622),
.A2(n_554),
.B(n_524),
.C(n_529),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_631),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_634),
.B(n_352),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_658),
.B(n_626),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_634),
.A2(n_324),
.B(n_354),
.C(n_459),
.Y(n_695)
);

NOR2x1_ASAP7_75t_L g696 ( 
.A(n_652),
.B(n_411),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_683),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_638),
.B(n_458),
.Y(n_698)
);

O2A1O1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_640),
.A2(n_487),
.B(n_546),
.C(n_523),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_677),
.Y(n_700)
);

O2A1O1Ixp5_ASAP7_75t_L g701 ( 
.A1(n_645),
.A2(n_606),
.B(n_585),
.C(n_474),
.Y(n_701)
);

BUFx4f_ASAP7_75t_L g702 ( 
.A(n_647),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_684),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_633),
.A2(n_482),
.B1(n_461),
.B2(n_457),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_686),
.B(n_598),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_632),
.B(n_600),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_666),
.A2(n_476),
.B1(n_493),
.B2(n_432),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_681),
.B(n_603),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_648),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_659),
.B(n_408),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_678),
.A2(n_608),
.B(n_604),
.Y(n_711)
);

NOR3xp33_ASAP7_75t_L g712 ( 
.A(n_675),
.B(n_500),
.C(n_498),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_649),
.A2(n_532),
.B(n_518),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_650),
.A2(n_532),
.B1(n_550),
.B2(n_518),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_667),
.B(n_542),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_636),
.Y(n_716)
);

O2A1O1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_691),
.A2(n_505),
.B(n_494),
.C(n_576),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_630),
.B(n_609),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_657),
.B(n_498),
.Y(n_719)
);

OAI22x1_ASAP7_75t_L g720 ( 
.A1(n_680),
.A2(n_574),
.B1(n_566),
.B2(n_389),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_685),
.A2(n_550),
.B1(n_577),
.B2(n_332),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_687),
.Y(n_722)
);

OAI321xp33_ASAP7_75t_L g723 ( 
.A1(n_680),
.A2(n_342),
.A3(n_336),
.B1(n_345),
.B2(n_339),
.C(n_322),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_676),
.A2(n_577),
.B(n_351),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_646),
.B(n_347),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_642),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_669),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_655),
.B(n_359),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_660),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_656),
.A2(n_653),
.B1(n_673),
.B2(n_670),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_662),
.B(n_361),
.Y(n_731)
);

CKINVDCx10_ASAP7_75t_R g732 ( 
.A(n_656),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_664),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_663),
.B(n_383),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_668),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_656),
.A2(n_577),
.B1(n_376),
.B2(n_379),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_641),
.A2(n_387),
.B(n_378),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_679),
.A2(n_396),
.B(n_395),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_688),
.A2(n_409),
.B(n_403),
.Y(n_739)
);

NOR2x1_ASAP7_75t_L g740 ( 
.A(n_644),
.B(n_665),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_635),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_690),
.A2(n_420),
.B(n_414),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_631),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_689),
.A2(n_424),
.B(n_421),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_631),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_671),
.A2(n_439),
.B(n_438),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_643),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_654),
.A2(n_577),
.B(n_446),
.Y(n_748)
);

OAI321xp33_ASAP7_75t_L g749 ( 
.A1(n_643),
.A2(n_471),
.A3(n_467),
.B1(n_472),
.B2(n_468),
.C(n_465),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_674),
.B(n_639),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_651),
.A2(n_479),
.B1(n_485),
.B2(n_477),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_682),
.B(n_400),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_674),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_682),
.B(n_500),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_654),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_661),
.A2(n_576),
.B(n_540),
.C(n_552),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_639),
.B(n_331),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_R g758 ( 
.A(n_639),
.B(n_337),
.Y(n_758)
);

AOI21x1_ASAP7_75t_L g759 ( 
.A1(n_637),
.A2(n_540),
.B(n_535),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_639),
.B(n_637),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_634),
.B(n_343),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_634),
.A2(n_344),
.B1(n_356),
.B2(n_349),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_638),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_648),
.B(n_552),
.Y(n_764)
);

OAI321xp33_ASAP7_75t_L g765 ( 
.A1(n_633),
.A2(n_557),
.A3(n_537),
.B1(n_538),
.B2(n_528),
.C(n_451),
.Y(n_765)
);

INVx11_ASAP7_75t_L g766 ( 
.A(n_647),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_638),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_683),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_672),
.A2(n_367),
.B(n_366),
.Y(n_769)
);

BUFx12f_ASAP7_75t_L g770 ( 
.A(n_647),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_634),
.A2(n_371),
.B(n_370),
.Y(n_771)
);

AOI22x1_ASAP7_75t_L g772 ( 
.A1(n_672),
.A2(n_563),
.B1(n_373),
.B2(n_374),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_634),
.B(n_381),
.Y(n_773)
);

A2O1A1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_634),
.A2(n_393),
.B(n_394),
.C(n_385),
.Y(n_774)
);

AO21x1_ASAP7_75t_L g775 ( 
.A1(n_633),
.A2(n_26),
.B(n_28),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_634),
.A2(n_398),
.B(n_397),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_672),
.A2(n_402),
.B(n_399),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_634),
.B(n_410),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_686),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_683),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_638),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_634),
.A2(n_426),
.B(n_425),
.Y(n_782)
);

O2A1O1Ixp5_ASAP7_75t_L g783 ( 
.A1(n_672),
.A2(n_429),
.B(n_434),
.C(n_427),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_640),
.A2(n_441),
.B(n_447),
.C(n_437),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_694),
.A2(n_463),
.B(n_460),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_692),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_692),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_743),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_713),
.A2(n_478),
.B(n_475),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_754),
.B(n_480),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_708),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_719),
.B(n_483),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_764),
.B(n_528),
.Y(n_793)
);

OAI21x1_ASAP7_75t_SL g794 ( 
.A1(n_775),
.A2(n_124),
.B(n_123),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_722),
.B(n_537),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_705),
.B(n_537),
.Y(n_796)
);

O2A1O1Ixp5_ASAP7_75t_L g797 ( 
.A1(n_783),
.A2(n_724),
.B(n_695),
.C(n_761),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_698),
.B(n_538),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_718),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_727),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_699),
.A2(n_419),
.B(n_443),
.C(n_405),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_757),
.A2(n_760),
.B(n_706),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_701),
.A2(n_473),
.B(n_464),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_763),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_700),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_767),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_704),
.B(n_538),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_693),
.A2(n_557),
.B1(n_491),
.B2(n_129),
.Y(n_808)
);

OA22x2_ASAP7_75t_L g809 ( 
.A1(n_720),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_809)
);

INVx5_ASAP7_75t_L g810 ( 
.A(n_692),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_716),
.Y(n_811)
);

AO31x2_ASAP7_75t_L g812 ( 
.A1(n_730),
.A2(n_34),
.A3(n_32),
.B(n_33),
.Y(n_812)
);

INVxp67_ASAP7_75t_SL g813 ( 
.A(n_745),
.Y(n_813)
);

INVx5_ASAP7_75t_L g814 ( 
.A(n_745),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_SL g815 ( 
.A1(n_745),
.A2(n_133),
.B(n_132),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_770),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_781),
.Y(n_817)
);

NAND2x1p5_ASAP7_75t_L g818 ( 
.A(n_703),
.B(n_709),
.Y(n_818)
);

BUFx12f_ASAP7_75t_L g819 ( 
.A(n_766),
.Y(n_819)
);

AOI22x1_ASAP7_75t_L g820 ( 
.A1(n_771),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_820)
);

NOR2xp67_ASAP7_75t_L g821 ( 
.A(n_762),
.B(n_141),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_714),
.B(n_35),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_714),
.B(n_36),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_SL g824 ( 
.A1(n_710),
.A2(n_734),
.B1(n_732),
.B2(n_696),
.Y(n_824)
);

OAI21xp33_ASAP7_75t_L g825 ( 
.A1(n_762),
.A2(n_36),
.B(n_37),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_784),
.A2(n_41),
.B(n_37),
.C(n_40),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_774),
.A2(n_778),
.B(n_773),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_729),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_702),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_697),
.B(n_42),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_768),
.B(n_42),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_748),
.A2(n_143),
.B(n_142),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_780),
.B(n_43),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_779),
.B(n_145),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_702),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_733),
.B(n_147),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_741),
.Y(n_837)
);

NOR2x1_ASAP7_75t_SL g838 ( 
.A(n_759),
.B(n_149),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_707),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_SL g840 ( 
.A(n_715),
.B(n_150),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_747),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_765),
.A2(n_782),
.B(n_776),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_736),
.B(n_44),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_725),
.B(n_712),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_726),
.B(n_46),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_753),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_723),
.B(n_153),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_726),
.B(n_46),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_740),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_755),
.B(n_47),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_735),
.B(n_47),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_SL g852 ( 
.A1(n_751),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_728),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_756),
.B(n_48),
.Y(n_854)
);

AOI22x1_ASAP7_75t_SL g855 ( 
.A1(n_749),
.A2(n_54),
.B1(n_49),
.B2(n_52),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_721),
.A2(n_160),
.B1(n_161),
.B2(n_158),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_731),
.B(n_52),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_772),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_769),
.A2(n_165),
.B(n_164),
.Y(n_859)
);

NAND3x1_ASAP7_75t_L g860 ( 
.A(n_721),
.B(n_54),
.C(n_55),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_717),
.B(n_55),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_737),
.B(n_56),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_777),
.A2(n_170),
.B1(n_171),
.B2(n_169),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_744),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_746),
.A2(n_60),
.B(n_57),
.C(n_58),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_738),
.A2(n_173),
.B(n_172),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_758),
.B(n_60),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_739),
.B(n_61),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_742),
.A2(n_177),
.B(n_175),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_754),
.B(n_62),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_L g871 ( 
.A(n_695),
.B(n_178),
.Y(n_871)
);

NOR2xp67_ASAP7_75t_L g872 ( 
.A(n_752),
.B(n_184),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_700),
.Y(n_873)
);

AO21x1_ASAP7_75t_L g874 ( 
.A1(n_784),
.A2(n_62),
.B(n_63),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_699),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_708),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_754),
.B(n_65),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_704),
.A2(n_235),
.B1(n_317),
.B2(n_316),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_766),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_708),
.Y(n_880)
);

INVx6_ASAP7_75t_L g881 ( 
.A(n_770),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_711),
.A2(n_189),
.B(n_187),
.Y(n_882)
);

AOI21x1_ASAP7_75t_L g883 ( 
.A1(n_757),
.A2(n_197),
.B(n_193),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_719),
.B(n_66),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_703),
.B(n_201),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_704),
.B(n_67),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_719),
.B(n_68),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_694),
.A2(n_203),
.B(n_202),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_719),
.B(n_68),
.Y(n_889)
);

NOR4xp25_ASAP7_75t_L g890 ( 
.A(n_723),
.B(n_69),
.C(n_70),
.D(n_71),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_754),
.B(n_204),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_719),
.B(n_69),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_754),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_704),
.B(n_71),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_754),
.B(n_213),
.Y(n_895)
);

AOI21xp33_ASAP7_75t_L g896 ( 
.A1(n_734),
.A2(n_72),
.B(n_73),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_708),
.Y(n_897)
);

NOR2x1_ASAP7_75t_SL g898 ( 
.A(n_692),
.B(n_215),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_754),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_711),
.A2(n_219),
.B(n_218),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_703),
.B(n_220),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_711),
.A2(n_222),
.B(n_221),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_708),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_708),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_SL g905 ( 
.A(n_704),
.B(n_74),
.C(n_75),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_708),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_698),
.B(n_74),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_829),
.Y(n_908)
);

NOR2x1_ASAP7_75t_SL g909 ( 
.A(n_810),
.B(n_223),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_907),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_787),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_885),
.B(n_225),
.Y(n_912)
);

OR3x4_ASAP7_75t_SL g913 ( 
.A(n_824),
.B(n_77),
.C(n_78),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_837),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_893),
.B(n_78),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_842),
.A2(n_844),
.B1(n_903),
.B2(n_880),
.Y(n_916)
);

NAND2x1p5_ASAP7_75t_L g917 ( 
.A(n_810),
.B(n_228),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_810),
.A2(n_814),
.B(n_882),
.Y(n_918)
);

OAI21x1_ASAP7_75t_SL g919 ( 
.A1(n_898),
.A2(n_262),
.B(n_310),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_837),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_885),
.B(n_901),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_880),
.Y(n_922)
);

NAND2x1p5_ASAP7_75t_L g923 ( 
.A(n_814),
.B(n_230),
.Y(n_923)
);

AO21x1_ASAP7_75t_L g924 ( 
.A1(n_900),
.A2(n_902),
.B(n_823),
.Y(n_924)
);

BUFx8_ASAP7_75t_SL g925 ( 
.A(n_819),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_817),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_899),
.B(n_79),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_804),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_825),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_929)
);

NAND2x1p5_ASAP7_75t_L g930 ( 
.A(n_814),
.B(n_231),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_806),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_789),
.A2(n_256),
.B(n_305),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_799),
.B(n_81),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_793),
.B(n_82),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_870),
.B(n_83),
.Y(n_935)
);

CKINVDCx6p67_ASAP7_75t_R g936 ( 
.A(n_816),
.Y(n_936)
);

NOR2xp67_ASAP7_75t_L g937 ( 
.A(n_879),
.B(n_232),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_904),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_800),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_905),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_805),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_877),
.Y(n_942)
);

NOR2x1_ASAP7_75t_SL g943 ( 
.A(n_858),
.B(n_234),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_822),
.A2(n_265),
.B(n_304),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_904),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_811),
.Y(n_946)
);

OR2x6_ASAP7_75t_SL g947 ( 
.A(n_835),
.B(n_839),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_807),
.B(n_85),
.Y(n_948)
);

OAI222xp33_ASAP7_75t_L g949 ( 
.A1(n_886),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.C1(n_89),
.C2(n_90),
.Y(n_949)
);

AO31x2_ASAP7_75t_L g950 ( 
.A1(n_874),
.A2(n_858),
.A3(n_838),
.B(n_826),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_818),
.Y(n_951)
);

AO31x2_ASAP7_75t_L g952 ( 
.A1(n_856),
.A2(n_87),
.A3(n_88),
.B(n_89),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_791),
.B(n_90),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_894),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_954)
);

BUFx2_ASAP7_75t_R g955 ( 
.A(n_843),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_828),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_850),
.Y(n_957)
);

INVx5_ASAP7_75t_L g958 ( 
.A(n_787),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_873),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_792),
.B(n_92),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_795),
.B(n_884),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_901),
.B(n_236),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_876),
.A2(n_267),
.B1(n_301),
.B2(n_300),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_834),
.B(n_94),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_788),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_897),
.A2(n_264),
.B1(n_297),
.B2(n_295),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_788),
.Y(n_967)
);

AOI31xp33_ASAP7_75t_L g968 ( 
.A1(n_852),
.A2(n_95),
.A3(n_96),
.B(n_97),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_906),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_821),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_SL g971 ( 
.A1(n_896),
.A2(n_99),
.B(n_100),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_834),
.B(n_836),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_846),
.Y(n_973)
);

INVx4_ASAP7_75t_SL g974 ( 
.A(n_881),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_853),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_887),
.B(n_889),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_881),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_841),
.Y(n_978)
);

AO21x2_ASAP7_75t_L g979 ( 
.A1(n_803),
.A2(n_246),
.B(n_286),
.Y(n_979)
);

NAND3xp33_ASAP7_75t_L g980 ( 
.A(n_854),
.B(n_101),
.C(n_102),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_872),
.A2(n_245),
.B1(n_285),
.B2(n_283),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_787),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_836),
.Y(n_983)
);

AO32x2_ASAP7_75t_L g984 ( 
.A1(n_890),
.A2(n_101),
.A3(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_841),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_892),
.B(n_105),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_820),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_849),
.B(n_107),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_841),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_790),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_809),
.B(n_867),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_796),
.B(n_108),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_891),
.A2(n_242),
.B1(n_279),
.B2(n_278),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_786),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_SL g995 ( 
.A1(n_855),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_860),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_801),
.A2(n_273),
.B(n_276),
.Y(n_997)
);

NOR2x1_ASAP7_75t_L g998 ( 
.A(n_786),
.B(n_110),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_830),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_861),
.A2(n_111),
.B1(n_113),
.B2(n_895),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_808),
.A2(n_813),
.B1(n_878),
.B2(n_847),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_831),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_851),
.A2(n_871),
.B(n_869),
.C(n_785),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_833),
.Y(n_1004)
);

CKINVDCx16_ASAP7_75t_R g1005 ( 
.A(n_855),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_815),
.B(n_888),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_845),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_848),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_857),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_812),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_862),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_812),
.Y(n_1012)
);

AO31x2_ASAP7_75t_L g1013 ( 
.A1(n_875),
.A2(n_864),
.A3(n_865),
.B(n_832),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_868),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_798),
.Y(n_1015)
);

BUFx2_ASAP7_75t_SL g1016 ( 
.A(n_863),
.Y(n_1016)
);

OA21x2_ASAP7_75t_L g1017 ( 
.A1(n_883),
.A2(n_859),
.B(n_866),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_840),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_837),
.Y(n_1019)
);

AOI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_839),
.A2(n_588),
.B1(n_704),
.B2(n_633),
.C(n_650),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_SL g1021 ( 
.A1(n_898),
.A2(n_775),
.B(n_794),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_802),
.A2(n_750),
.B(n_658),
.Y(n_1022)
);

OA21x2_ASAP7_75t_L g1023 ( 
.A1(n_797),
.A2(n_827),
.B(n_842),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_893),
.B(n_899),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_817),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_817),
.Y(n_1026)
);

AOI221xp5_ASAP7_75t_L g1027 ( 
.A1(n_839),
.A2(n_588),
.B1(n_704),
.B2(n_633),
.C(n_650),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_907),
.A2(n_842),
.B1(n_634),
.B2(n_825),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_907),
.A2(n_842),
.B1(n_634),
.B2(n_825),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_787),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_837),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_837),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_907),
.A2(n_842),
.B1(n_634),
.B2(n_825),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_837),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_SL g1035 ( 
.A1(n_824),
.A2(n_663),
.B1(n_839),
.B2(n_704),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_804),
.B(n_806),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_817),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_893),
.B(n_899),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_1024),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_1036),
.B(n_928),
.Y(n_1040)
);

AOI222xp33_ASAP7_75t_L g1041 ( 
.A1(n_1020),
.A2(n_1027),
.B1(n_949),
.B2(n_929),
.C1(n_954),
.C2(n_940),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_926),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_921),
.B(n_972),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_908),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_1026),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_920),
.Y(n_1046)
);

OA21x2_ASAP7_75t_L g1047 ( 
.A1(n_924),
.A2(n_1022),
.B(n_1003),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_958),
.Y(n_1048)
);

AO21x2_ASAP7_75t_L g1049 ( 
.A1(n_932),
.A2(n_1021),
.B(n_918),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_921),
.B(n_912),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_920),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_942),
.B(n_957),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_983),
.B(n_912),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_1038),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_922),
.B(n_938),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_962),
.B(n_977),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1035),
.A2(n_990),
.B1(n_1011),
.B2(n_1018),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_989),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1019),
.Y(n_1059)
);

INVxp33_ASAP7_75t_SL g1060 ( 
.A(n_1037),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_962),
.B(n_939),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_991),
.B(n_927),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1031),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_946),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_916),
.B(n_976),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_951),
.B(n_1025),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_945),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_935),
.B(n_964),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_910),
.A2(n_980),
.B1(n_1033),
.B2(n_1029),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_914),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1032),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1034),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_988),
.B(n_996),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1009),
.B(n_995),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_931),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_975),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_915),
.B(n_1004),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_956),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_969),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_974),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_999),
.B(n_1002),
.Y(n_1081)
);

OR2x6_ASAP7_75t_L g1082 ( 
.A(n_1018),
.B(n_917),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_960),
.B(n_961),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_958),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_941),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1007),
.B(n_1014),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_958),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_925),
.Y(n_1088)
);

AO31x2_ASAP7_75t_L g1089 ( 
.A1(n_1001),
.A2(n_1007),
.A3(n_943),
.B(n_1008),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_959),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_973),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_974),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_986),
.B(n_1005),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_911),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_955),
.B(n_948),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_1030),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_933),
.B(n_953),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_936),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_1030),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_934),
.B(n_1015),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_965),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1028),
.A2(n_1023),
.B(n_944),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_967),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_947),
.B(n_998),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_982),
.Y(n_1105)
);

AO21x2_ASAP7_75t_L g1106 ( 
.A1(n_997),
.A2(n_979),
.B(n_1012),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_992),
.B(n_978),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_982),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_985),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_971),
.B(n_1000),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_923),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_994),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_937),
.B(n_1006),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1010),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_SL g1115 ( 
.A(n_1016),
.B(n_930),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_952),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_919),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_970),
.B(n_984),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_984),
.B(n_987),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_984),
.B(n_952),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1013),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1013),
.B(n_950),
.Y(n_1122)
);

INVx5_ASAP7_75t_L g1123 ( 
.A(n_909),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_952),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_909),
.B(n_943),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_968),
.B(n_993),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_963),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_966),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_981),
.B(n_913),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1017),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1062),
.B(n_1068),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1121),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_1039),
.B(n_1040),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1086),
.B(n_1097),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_1066),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1041),
.A2(n_1126),
.B1(n_1110),
.B2(n_1069),
.Y(n_1136)
);

INVx5_ASAP7_75t_L g1137 ( 
.A(n_1048),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1086),
.B(n_1097),
.Y(n_1138)
);

INVx4_ASAP7_75t_R g1139 ( 
.A(n_1084),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1074),
.B(n_1077),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1076),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1079),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1083),
.B(n_1073),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1055),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1048),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1042),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_1053),
.B(n_1050),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1083),
.B(n_1052),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1054),
.B(n_1057),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1100),
.B(n_1054),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_1081),
.B(n_1107),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_1075),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1093),
.B(n_1053),
.Y(n_1153)
);

CKINVDCx6p67_ASAP7_75t_R g1154 ( 
.A(n_1088),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1044),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1050),
.B(n_1056),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1050),
.B(n_1056),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1045),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1043),
.B(n_1095),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1126),
.B(n_1129),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1067),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1061),
.B(n_1056),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_1048),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1078),
.B(n_1070),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1104),
.B(n_1090),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1066),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1064),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1101),
.B(n_1103),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1075),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1087),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1085),
.B(n_1070),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1046),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1071),
.B(n_1072),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1041),
.A2(n_1069),
.B1(n_1118),
.B2(n_1065),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1051),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1059),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1065),
.B(n_1063),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1096),
.B(n_1099),
.Y(n_1178)
);

AND2x4_ASAP7_75t_SL g1179 ( 
.A(n_1087),
.B(n_1044),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_1109),
.B(n_1112),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1105),
.B(n_1108),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1091),
.B(n_1058),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1127),
.B(n_1128),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1114),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1099),
.B(n_1084),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1119),
.B(n_1089),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1089),
.B(n_1113),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1116),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1060),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1089),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1089),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1060),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1172),
.Y(n_1193)
);

INVxp67_ASAP7_75t_SL g1194 ( 
.A(n_1144),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1140),
.B(n_1094),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1175),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_1137),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1148),
.B(n_1082),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1136),
.A2(n_1160),
.B1(n_1174),
.B2(n_1149),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1176),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1186),
.B(n_1120),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1186),
.B(n_1122),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1133),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1188),
.B(n_1124),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1135),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1134),
.B(n_1138),
.Y(n_1206)
);

NOR2xp67_ASAP7_75t_L g1207 ( 
.A(n_1152),
.B(n_1098),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1135),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1141),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1142),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1151),
.B(n_1047),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1134),
.B(n_1115),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1138),
.B(n_1115),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1167),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1156),
.B(n_1117),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1143),
.B(n_1047),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1131),
.B(n_1111),
.Y(n_1217)
);

NOR2xp67_ASAP7_75t_L g1218 ( 
.A(n_1152),
.B(n_1098),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1150),
.B(n_1049),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1157),
.B(n_1117),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1132),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_1164),
.B(n_1080),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1136),
.B(n_1111),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1144),
.B(n_1111),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1160),
.B(n_1049),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1171),
.B(n_1102),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1173),
.B(n_1102),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_1146),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1165),
.B(n_1125),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1182),
.B(n_1153),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1161),
.B(n_1123),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1147),
.B(n_1106),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1147),
.B(n_1162),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1232),
.B(n_1187),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1203),
.B(n_1183),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1206),
.B(n_1183),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1221),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1201),
.B(n_1190),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1201),
.B(n_1190),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1193),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1231),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1196),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1202),
.B(n_1191),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1202),
.B(n_1191),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1219),
.B(n_1187),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1215),
.B(n_1184),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1228),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1212),
.B(n_1181),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1213),
.B(n_1169),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1194),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1204),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1230),
.B(n_1155),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1225),
.B(n_1216),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1211),
.B(n_1177),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1233),
.B(n_1166),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1217),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1200),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1197),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1224),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1209),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1204),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1194),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1226),
.B(n_1177),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1210),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1214),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1240),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1240),
.Y(n_1267)
);

AND2x2_ASAP7_75t_SL g1268 ( 
.A(n_1250),
.B(n_1199),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1256),
.B(n_1259),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1242),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1257),
.Y(n_1271)
);

NAND2xp33_ASAP7_75t_SL g1272 ( 
.A(n_1247),
.B(n_1199),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1253),
.B(n_1198),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1260),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1246),
.A2(n_1223),
.B1(n_1220),
.B2(n_1215),
.Y(n_1275)
);

NOR2x1p5_ASAP7_75t_SL g1276 ( 
.A(n_1254),
.B(n_1130),
.Y(n_1276)
);

NAND2x1_ASAP7_75t_SL g1277 ( 
.A(n_1262),
.B(n_1253),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1236),
.B(n_1215),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1264),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1264),
.Y(n_1280)
);

NAND4xp25_ASAP7_75t_L g1281 ( 
.A(n_1249),
.B(n_1218),
.C(n_1207),
.D(n_1222),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1265),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1234),
.B(n_1229),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1254),
.B(n_1227),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1246),
.Y(n_1285)
);

NAND2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1258),
.B(n_1197),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1268),
.A2(n_1220),
.B1(n_1246),
.B2(n_1245),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1266),
.Y(n_1288)
);

AOI322xp5_ASAP7_75t_L g1289 ( 
.A1(n_1272),
.A2(n_1238),
.A3(n_1239),
.B1(n_1235),
.B2(n_1252),
.C1(n_1248),
.C2(n_1159),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1275),
.A2(n_1245),
.B1(n_1263),
.B2(n_1258),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1267),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1270),
.Y(n_1292)
);

AO221x1_ASAP7_75t_L g1293 ( 
.A1(n_1271),
.A2(n_1241),
.B1(n_1237),
.B2(n_1261),
.C(n_1251),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_1269),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1274),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1279),
.Y(n_1296)
);

OAI32xp33_ASAP7_75t_L g1297 ( 
.A1(n_1272),
.A2(n_1278),
.A3(n_1284),
.B1(n_1285),
.B2(n_1281),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1280),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1268),
.B(n_1278),
.C(n_1284),
.Y(n_1299)
);

NAND2xp33_ASAP7_75t_SL g1300 ( 
.A(n_1277),
.B(n_1088),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1273),
.B(n_1234),
.Y(n_1301)
);

NOR3xp33_ASAP7_75t_L g1302 ( 
.A(n_1297),
.B(n_1208),
.C(n_1205),
.Y(n_1302)
);

NOR2xp67_ASAP7_75t_L g1303 ( 
.A(n_1299),
.B(n_1282),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1300),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1294),
.B(n_1283),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1287),
.A2(n_1285),
.B1(n_1220),
.B2(n_1286),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1288),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1301),
.B(n_1234),
.Y(n_1308)
);

AOI221xp5_ASAP7_75t_L g1309 ( 
.A1(n_1302),
.A2(n_1290),
.B1(n_1293),
.B2(n_1296),
.C(n_1295),
.Y(n_1309)
);

NAND4xp25_ASAP7_75t_L g1310 ( 
.A(n_1303),
.B(n_1289),
.C(n_1255),
.D(n_1195),
.Y(n_1310)
);

AOI322xp5_ASAP7_75t_L g1311 ( 
.A1(n_1304),
.A2(n_1289),
.A3(n_1239),
.B1(n_1238),
.B2(n_1244),
.C1(n_1243),
.C2(n_1292),
.Y(n_1311)
);

OAI21xp33_ASAP7_75t_L g1312 ( 
.A1(n_1304),
.A2(n_1276),
.B(n_1263),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1306),
.B(n_1286),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1310),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1312),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1313),
.B(n_1308),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1309),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1311),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1313),
.A2(n_1307),
.B(n_1305),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1316),
.B(n_1189),
.Y(n_1320)
);

NOR3x1_ASAP7_75t_L g1321 ( 
.A(n_1317),
.B(n_1158),
.C(n_1092),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1318),
.B(n_1291),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_SL g1323 ( 
.A1(n_1322),
.A2(n_1315),
.B(n_1319),
.Y(n_1323)
);

NOR2x1_ASAP7_75t_L g1324 ( 
.A(n_1320),
.B(n_1189),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1323),
.B(n_1314),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1325),
.B(n_1321),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1326),
.B(n_1324),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1326),
.B(n_1314),
.Y(n_1328)
);

XNOR2xp5_ASAP7_75t_L g1329 ( 
.A(n_1327),
.B(n_1179),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1328),
.A2(n_1154),
.B1(n_1192),
.B2(n_1179),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1329),
.A2(n_1139),
.B(n_1180),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1330),
.A2(n_1192),
.B(n_1185),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1332),
.A2(n_1185),
.B(n_1168),
.Y(n_1333)
);

AOI21xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1331),
.A2(n_1170),
.B(n_1145),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1334),
.A2(n_1178),
.B(n_1298),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1335),
.B(n_1333),
.Y(n_1336)
);

AOI21xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1336),
.A2(n_1163),
.B(n_1145),
.Y(n_1337)
);


endmodule