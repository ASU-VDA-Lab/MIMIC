module fake_jpeg_6592_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR3xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.C(n_1),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_24),
.Y(n_45)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_24),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_17),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_23),
.B1(n_29),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_49),
.B1(n_52),
.B2(n_17),
.Y(n_72)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_51),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_19),
.B1(n_28),
.B2(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_19),
.B1(n_28),
.B2(n_29),
.Y(n_52)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_19),
.B1(n_23),
.B2(n_34),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_60),
.Y(n_112)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_65),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_35),
.Y(n_60)
);

FAx1_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_39),
.CI(n_34),
.CON(n_61),
.SN(n_61)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_61),
.B(n_63),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_22),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_39),
.B(n_36),
.C(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_68),
.Y(n_95)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_36),
.CI(n_37),
.CON(n_68),
.SN(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_83),
.B(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_16),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_22),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_16),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_77),
.Y(n_94)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_79),
.Y(n_99)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_82),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_33),
.B1(n_21),
.B2(n_20),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_36),
.B(n_26),
.C(n_31),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_68),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_36),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_109),
.C(n_104),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_37),
.C(n_50),
.Y(n_109)
);

AOI32xp33_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_37),
.A3(n_50),
.B1(n_33),
.B2(n_40),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_94),
.B(n_89),
.C(n_78),
.D(n_37),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_121),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_99),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_68),
.B1(n_59),
.B2(n_87),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_116),
.A2(n_124),
.B(n_126),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_58),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_125),
.B(n_27),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_122),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_65),
.B1(n_83),
.B2(n_60),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_127),
.B1(n_131),
.B2(n_133),
.Y(n_150)
);

OAI221xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_71),
.B1(n_77),
.B2(n_64),
.C(n_67),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_74),
.B(n_86),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_81),
.B(n_84),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_80),
.B1(n_66),
.B2(n_40),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_129),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_37),
.B(n_40),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_132),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_40),
.B1(n_20),
.B2(n_30),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_16),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_104),
.B1(n_102),
.B2(n_112),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_136),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_50),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_137),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_32),
.B1(n_27),
.B2(n_18),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_108),
.B1(n_105),
.B2(n_62),
.Y(n_155)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_140),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_103),
.B1(n_91),
.B2(n_93),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_117),
.B1(n_123),
.B2(n_125),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_144),
.B(n_148),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_118),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_147),
.C(n_153),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

HB1xp67_ASAP7_75t_SL g175 ( 
.A(n_151),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_116),
.B(n_13),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_155),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_108),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_160),
.C(n_161),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_32),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_88),
.C(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_32),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_166),
.A2(n_140),
.B(n_32),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_129),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_179),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_129),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_156),
.C(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_143),
.B(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_0),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_141),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_27),
.B1(n_18),
.B2(n_88),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_188),
.A2(n_144),
.B1(n_142),
.B2(n_158),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_182),
.A2(n_158),
.B(n_161),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_203),
.B(n_180),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_200),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_201),
.C(n_185),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_146),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_195),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_153),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_171),
.B(n_179),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_197),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_172),
.C(n_176),
.Y(n_201)
);

NAND2x1p5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_151),
.Y(n_203)
);

BUFx4f_ASAP7_75t_SL g204 ( 
.A(n_178),
.Y(n_204)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_154),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_183),
.B1(n_168),
.B2(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_193),
.C(n_195),
.Y(n_230)
);

XOR2x2_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_166),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_190),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_170),
.B1(n_181),
.B2(n_187),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_203),
.B(n_202),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_150),
.B1(n_169),
.B2(n_188),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_150),
.B1(n_186),
.B2(n_177),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_200),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_88),
.B1(n_27),
.B2(n_5),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_221),
.Y(n_231)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_204),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_225),
.B(n_226),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_204),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_201),
.B(n_191),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_212),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_214),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_207),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_210),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_236),
.B1(n_206),
.B2(n_208),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_234),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_216),
.B1(n_228),
.B2(n_224),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_13),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_1),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_230),
.B1(n_209),
.B2(n_15),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_242),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_237),
.A2(n_209),
.B1(n_15),
.B2(n_14),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_2),
.B(n_5),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_231),
.C(n_233),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_2),
.B(n_5),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_246),
.B(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_2),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_244),
.A3(n_7),
.B1(n_9),
.B2(n_10),
.C1(n_6),
.C2(n_12),
.Y(n_250)
);

OA21x2_ASAP7_75t_SL g253 ( 
.A1(n_250),
.A2(n_252),
.B(n_11),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_240),
.C(n_10),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_254),
.Y(n_255)
);

OA21x2_ASAP7_75t_SL g254 ( 
.A1(n_251),
.A2(n_6),
.B(n_10),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_6),
.B(n_11),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_11),
.Y(n_257)
);


endmodule