module fake_jpeg_14379_n_435 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_435);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_435;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_6),
.B(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_13),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_47),
.B(n_56),
.Y(n_120)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_51),
.Y(n_136)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_13),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_57),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_91),
.Y(n_96)
);

INVx2_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_83),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_24),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_26),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_88),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_24),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_92),
.Y(n_130)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_31),
.B1(n_44),
.B2(n_36),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_98),
.A2(n_102),
.B1(n_113),
.B2(n_126),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_29),
.B1(n_44),
.B2(n_36),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_25),
.B1(n_27),
.B2(n_45),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_40),
.B1(n_45),
.B2(n_42),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_116),
.A2(n_62),
.A3(n_22),
.B1(n_26),
.B2(n_37),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_27),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_54),
.B(n_25),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_0),
.C(n_1),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_48),
.A2(n_91),
.B1(n_50),
.B2(n_51),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_57),
.A2(n_40),
.B1(n_35),
.B2(n_46),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_134),
.B1(n_140),
.B2(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_55),
.B(n_42),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_133),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_61),
.A2(n_78),
.B1(n_86),
.B2(n_82),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_32),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_141),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_66),
.A2(n_46),
.B1(n_44),
.B2(n_36),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_75),
.B(n_32),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_65),
.A2(n_29),
.B1(n_30),
.B2(n_22),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_64),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_161),
.C(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_30),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_168),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_53),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_149),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_108),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_151),
.B(n_153),
.Y(n_223)
);

OR2x4_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_22),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_152),
.B(n_171),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_154),
.B(n_169),
.Y(n_198)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_67),
.B1(n_80),
.B2(n_71),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_159),
.A2(n_189),
.B1(n_146),
.B2(n_144),
.Y(n_196)
);

BUFx24_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_160),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_70),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_95),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_60),
.B1(n_68),
.B2(n_90),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_97),
.B1(n_101),
.B2(n_103),
.Y(n_197)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_167),
.B(n_170),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_0),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_37),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_99),
.B(n_107),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_106),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_104),
.B(n_74),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_0),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_110),
.B(n_125),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_176),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_114),
.B(n_37),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_177),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_34),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_34),
.C(n_16),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_100),
.B(n_1),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_186),
.Y(n_204)
);

INVx4_ASAP7_75t_SL g181 ( 
.A(n_95),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

AO22x2_ASAP7_75t_L g186 ( 
.A1(n_97),
.A2(n_16),
.B1(n_34),
.B2(n_3),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_187),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_222)
);

NAND2x1_ASAP7_75t_L g188 ( 
.A(n_122),
.B(n_112),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_188),
.A2(n_34),
.B(n_16),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_128),
.A2(n_126),
.B1(n_140),
.B2(n_138),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_196),
.A2(n_212),
.B1(n_219),
.B2(n_158),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_197),
.A2(n_216),
.B1(n_165),
.B2(n_173),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_149),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_208),
.C(n_221),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_124),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_148),
.B(n_129),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_218),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_192),
.A2(n_147),
.B1(n_183),
.B2(n_152),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_158),
.A2(n_135),
.B1(n_101),
.B2(n_103),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_SL g248 ( 
.A1(n_214),
.A2(n_179),
.B(n_184),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_147),
.A2(n_146),
.B1(n_121),
.B2(n_142),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_121),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_160),
.A2(n_144),
.B1(n_142),
.B2(n_94),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_160),
.A2(n_1),
.B(n_2),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_220),
.A2(n_188),
.B(n_172),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_161),
.B(n_34),
.C(n_16),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_172),
.C(n_188),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_228),
.A2(n_205),
.B(n_194),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_174),
.B(n_2),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_2),
.Y(n_246)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_232),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_221),
.C(n_225),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_156),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_234),
.B(n_237),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_223),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_238),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_219),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_247),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_199),
.B(n_156),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_240),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_166),
.B1(n_164),
.B2(n_160),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_241),
.A2(n_255),
.B1(n_193),
.B2(n_217),
.Y(n_294)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_200),
.A2(n_164),
.B1(n_175),
.B2(n_150),
.Y(n_245)
);

AOI22x1_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_253),
.B1(n_196),
.B2(n_209),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_246),
.B(n_254),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_248),
.A2(n_197),
.B1(n_209),
.B2(n_222),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_199),
.B(n_229),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_251),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_250),
.A2(n_263),
.B(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_161),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_200),
.A2(n_186),
.B1(n_157),
.B2(n_185),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_211),
.B(n_151),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_204),
.A2(n_186),
.B1(n_190),
.B2(n_187),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_215),
.B(n_153),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_259),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_258),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_201),
.B(n_186),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_155),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_204),
.B(n_227),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_205),
.B(n_208),
.Y(n_264)
);

OAI32xp33_ASAP7_75t_L g265 ( 
.A1(n_194),
.A2(n_186),
.A3(n_162),
.B1(n_181),
.B2(n_191),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_216),
.B1(n_206),
.B2(n_228),
.Y(n_280)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_271),
.A2(n_294),
.B1(n_261),
.B2(n_257),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_247),
.A2(n_207),
.B(n_209),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_273),
.A2(n_286),
.B(n_265),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_237),
.A2(n_207),
.B(n_230),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_279),
.A2(n_291),
.B(n_292),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_233),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_284),
.C(n_285),
.Y(n_308)
);

AO22x1_ASAP7_75t_SL g283 ( 
.A1(n_253),
.A2(n_210),
.B1(n_226),
.B2(n_213),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_294),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_264),
.C(n_263),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_195),
.C(n_224),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_241),
.B(n_255),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_195),
.C(n_224),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_243),
.C(n_252),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_250),
.A2(n_231),
.B(n_210),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_236),
.A2(n_203),
.B(n_193),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_245),
.B(n_262),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_298),
.B(n_310),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_306),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_249),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_311),
.C(n_314),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_256),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_301),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_267),
.B(n_234),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_305),
.Y(n_327)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_304),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_SL g305 ( 
.A(n_266),
.B(n_254),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_269),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_286),
.A2(n_239),
.B1(n_238),
.B2(n_235),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_307),
.A2(n_266),
.B1(n_270),
.B2(n_280),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_287),
.A2(n_240),
.B1(n_235),
.B2(n_251),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_309),
.A2(n_319),
.B1(n_321),
.B2(n_272),
.Y(n_325)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_268),
.Y(n_312)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_282),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_315),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_246),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_296),
.B(n_232),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_232),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_318),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_260),
.C(n_258),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_324),
.C(n_279),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_296),
.B(n_257),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_217),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_320),
.Y(n_328)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_248),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_280),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_181),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_325),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_333),
.B1(n_334),
.B2(n_343),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_307),
.A2(n_266),
.B1(n_270),
.B2(n_280),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_302),
.A2(n_322),
.B1(n_298),
.B2(n_310),
.Y(n_334)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_321),
.A2(n_268),
.B1(n_278),
.B2(n_283),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_278),
.Y(n_338)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_283),
.Y(n_341)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_341),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_323),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_299),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_302),
.A2(n_289),
.B1(n_281),
.B2(n_274),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_347),
.C(n_311),
.Y(n_355)
);

MAJx2_ASAP7_75t_L g347 ( 
.A(n_308),
.B(n_291),
.C(n_274),
.Y(n_347)
);

XNOR2x1_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_290),
.Y(n_348)
);

XOR2x2_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_324),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_290),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_349),
.B(n_308),
.Y(n_351)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_355),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_317),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_354),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_304),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_330),
.B(n_319),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_359),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_314),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_343),
.C(n_347),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_368),
.C(n_345),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_305),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_366),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_277),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_364),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_342),
.B(n_277),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_297),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_367),
.A2(n_370),
.B1(n_346),
.B2(n_334),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_297),
.C(n_191),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_327),
.B(n_2),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_352),
.A2(n_329),
.B1(n_363),
.B2(n_357),
.Y(n_373)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

NOR3xp33_ASAP7_75t_SL g375 ( 
.A(n_361),
.B(n_344),
.C(n_335),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_375),
.B(n_377),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_358),
.A2(n_344),
.B(n_340),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_378),
.A2(n_379),
.B(n_383),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_348),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_360),
.C(n_362),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g382 ( 
.A(n_355),
.B(n_344),
.CI(n_333),
.CON(n_382),
.SN(n_382)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_182),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_350),
.A2(n_340),
.B(n_331),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_332),
.C(n_339),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_386),
.B(n_339),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_383),
.A2(n_369),
.B1(n_356),
.B2(n_365),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_389),
.A2(n_379),
.B1(n_382),
.B2(n_191),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_397),
.C(n_380),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_366),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_395),
.Y(n_401)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_396),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_372),
.A2(n_365),
.B1(n_356),
.B2(n_369),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_394),
.A2(n_384),
.B1(n_385),
.B2(n_375),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_381),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_354),
.C(n_364),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_378),
.A2(n_370),
.B(n_332),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_398),
.A2(n_399),
.B(n_3),
.Y(n_408)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_400),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_403),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_371),
.C(n_376),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_R g404 ( 
.A(n_397),
.B(n_376),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_404),
.B(n_410),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_393),
.Y(n_405)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_405),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_408),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_388),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_409),
.B(n_398),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_387),
.A2(n_4),
.B(n_7),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_392),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_390),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_412),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_407),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_414),
.B(n_418),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_401),
.B(n_394),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_415),
.B(n_403),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_422),
.A2(n_413),
.B1(n_409),
.B2(n_411),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_424),
.C(n_425),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_419),
.B(n_392),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_406),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_419),
.C(n_417),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_428),
.C(n_429),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_421),
.B(n_389),
.C(n_16),
.Y(n_429)
);

O2A1O1Ixp33_ASAP7_75t_SL g431 ( 
.A1(n_426),
.A2(n_420),
.B(n_8),
.C(n_9),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_431),
.A2(n_4),
.B(n_8),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_430),
.C(n_9),
.Y(n_433)
);

O2A1O1Ixp33_ASAP7_75t_L g434 ( 
.A1(n_433),
.A2(n_12),
.B(n_4),
.C(n_9),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_12),
.Y(n_435)
);


endmodule