module fake_jpeg_17703_n_89 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_89);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_89;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_0),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_0),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_53),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_35),
.C(n_32),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_1),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_16),
.B1(n_26),
.B2(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_2),
.Y(n_64)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_64),
.B1(n_63),
.B2(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_72),
.Y(n_77)
);

AOI32xp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_15),
.A3(n_24),
.B1(n_5),
.B2(n_6),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_76),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_18),
.B1(n_23),
.B2(n_8),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_3),
.B(n_4),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_73),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_3),
.Y(n_76)
);

OAI21x1_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_12),
.B(n_13),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_69),
.B(n_75),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_82),
.Y(n_83)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_78),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_76),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_80),
.B(n_67),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_70),
.B(n_74),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_14),
.B(n_19),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_20),
.Y(n_89)
);


endmodule