module fake_ariane_724_n_2877 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_39, n_155, n_127, n_2877);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_2877;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_416;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_524;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_520;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_338;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_559;
wire n_2233;
wire n_2663;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_2782;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_334;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_533;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_355;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_2703;
wire n_696;
wire n_1442;
wire n_482;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_555;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_436;
wire n_2871;
wire n_2745;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_2628;
wire n_619;
wire n_337;
wire n_967;
wire n_1083;
wire n_437;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_470;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_2294;
wire n_489;
wire n_2274;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_397;
wire n_2467;
wire n_2768;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_404;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_347;
wire n_2434;
wire n_1042;
wire n_2311;
wire n_1234;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_552;
wire n_348;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_379;
wire n_2834;
wire n_2483;
wire n_441;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1609;
wire n_1053;
wire n_481;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_529;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_590;
wire n_699;
wire n_727;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_545;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_2853;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_390;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2861;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_388;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_342;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_358;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_463;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_374;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_586;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_354;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_335;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_1958;
wire n_2747;
wire n_467;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2431;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_413;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_361;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_453;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_540;
wire n_2624;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_493;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2809;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_353;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_385;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_399;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2580;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_1459;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_369;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_550;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_459;
wire n_2515;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_2869;
wire n_450;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_1946;
wire n_774;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_537;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_389;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_719;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1252;
wire n_2239;
wire n_1129;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_1299;
wire n_457;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_431;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_357;
wire n_1251;
wire n_412;
wire n_1989;
wire n_1421;
wire n_447;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_2851;
wire n_2823;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_43),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_63),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_290),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_142),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_72),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_14),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_3),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_131),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_184),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_82),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_244),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_177),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_322),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_333),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_140),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_69),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_294),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_36),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_180),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_223),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_225),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_291),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_40),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_89),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_281),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_222),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_36),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_293),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_68),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_318),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_232),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_241),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_148),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_320),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_198),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_134),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_48),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_111),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_75),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_9),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_288),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_4),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_224),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_330),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_29),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_297),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_195),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_193),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_199),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_243),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_121),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_300),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_90),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_249),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_33),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_30),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_113),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_177),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_85),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_236),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_68),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_26),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_155),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_271),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_136),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_161),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_287),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_150),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_39),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_258),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_135),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_26),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_207),
.Y(n_408)
);

INVxp33_ASAP7_75t_L g409 ( 
.A(n_143),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_323),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_0),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_219),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_192),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_158),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_16),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_217),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_101),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_136),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_125),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_313),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_211),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_201),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_254),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_168),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_265),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_310),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_218),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_128),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_66),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_306),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_103),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_256),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_327),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_273),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_105),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_74),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_298),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_99),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_127),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_140),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_280),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_148),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_18),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_174),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_189),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_233),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_174),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_179),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_71),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_67),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_19),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_123),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_117),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_81),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_29),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_49),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_30),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_9),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_166),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_175),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_234),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_277),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_314),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_8),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_206),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_186),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_131),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_79),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_53),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_235),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_215),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_315),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_261),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_109),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_302),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_106),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_286),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_226),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_104),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_231),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_146),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_13),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_156),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_214),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_110),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_130),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_182),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_245),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_7),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_252),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_228),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_316),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_301),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_138),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_309),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_59),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_331),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_187),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_269),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_73),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_283),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_35),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_100),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_305),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_73),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_6),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_16),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_299),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_91),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_135),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_325),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_146),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_79),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_171),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_329),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_62),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_35),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_292),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_197),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_200),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_170),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_122),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_38),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_141),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_312),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_103),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_10),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_319),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_278),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_53),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_257),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_161),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_77),
.Y(n_534)
);

BUFx8_ASAP7_75t_SL g535 ( 
.A(n_154),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_181),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_101),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_12),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_60),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_183),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_106),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_25),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_112),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_94),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_296),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_200),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_109),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_75),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_151),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_48),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_227),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_321),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_98),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_328),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_196),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_170),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_133),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_230),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_28),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_239),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_279),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_188),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_172),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_14),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_63),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_204),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_162),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_96),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_94),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_212),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_267),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_49),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_179),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_197),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_262),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_229),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_132),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_107),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_70),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_164),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_295),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_33),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_282),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_311),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_144),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_188),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_81),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_82),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_176),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_111),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_317),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_108),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_43),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_97),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_274),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_308),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_41),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_260),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_120),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_206),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_180),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_93),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_8),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_88),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_4),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_187),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_102),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_112),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_192),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_88),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_87),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_121),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_97),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_124),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_326),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_194),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_250),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_147),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_5),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_208),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_46),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_126),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_17),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_157),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_307),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_198),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_62),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_145),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_50),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_345),
.Y(n_630)
);

INVxp33_ASAP7_75t_L g631 ( 
.A(n_535),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_340),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_340),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_354),
.Y(n_634)
);

INVxp33_ASAP7_75t_SL g635 ( 
.A(n_352),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_386),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_354),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g638 ( 
.A(n_352),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_366),
.Y(n_639)
);

INVxp67_ASAP7_75t_SL g640 ( 
.A(n_391),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_562),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_366),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_374),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_390),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_562),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_390),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_405),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_440),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_391),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_391),
.B(n_0),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_345),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_395),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_423),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_395),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_374),
.Y(n_655)
);

BUFx2_ASAP7_75t_SL g656 ( 
.A(n_473),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_334),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_462),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_491),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_399),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_526),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_399),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_414),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_414),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_374),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_427),
.Y(n_666)
);

BUFx5_ASAP7_75t_L g667 ( 
.A(n_427),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_428),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_428),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_423),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_435),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_374),
.Y(n_672)
);

INVxp33_ASAP7_75t_SL g673 ( 
.A(n_335),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_409),
.Y(n_674)
);

INVxp33_ASAP7_75t_L g675 ( 
.A(n_343),
.Y(n_675)
);

INVxp33_ASAP7_75t_L g676 ( 
.A(n_343),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_431),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_431),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_438),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_346),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_438),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_406),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_464),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_346),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_349),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_464),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_374),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_479),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_479),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_485),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_485),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_374),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_423),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_337),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_557),
.Y(n_695)
);

INVxp33_ASAP7_75t_SL g696 ( 
.A(n_338),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_339),
.Y(n_697)
);

INVxp33_ASAP7_75t_SL g698 ( 
.A(n_341),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_557),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_416),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_557),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_574),
.Y(n_702)
);

INVxp33_ASAP7_75t_SL g703 ( 
.A(n_342),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_574),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_494),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_344),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_350),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_494),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_345),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_574),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_353),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_532),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_358),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_415),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_523),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_616),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_616),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_616),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_556),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_590),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_361),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_363),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_568),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_614),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_532),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_552),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_552),
.Y(n_727)
);

INVxp33_ASAP7_75t_SL g728 ( 
.A(n_369),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_561),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_561),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_571),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_571),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_584),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_370),
.Y(n_734)
);

CKINVDCx16_ASAP7_75t_R g735 ( 
.A(n_375),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_558),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_568),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_584),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_618),
.Y(n_739)
);

CKINVDCx16_ASAP7_75t_R g740 ( 
.A(n_375),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_595),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_595),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_572),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_572),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_572),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_371),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_619),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_601),
.Y(n_748)
);

INVxp33_ASAP7_75t_SL g749 ( 
.A(n_372),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_601),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_415),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_601),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_373),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_415),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_415),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_415),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_415),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_507),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_379),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_507),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_421),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_507),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_507),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_507),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_507),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_514),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_656),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_643),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_656),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_636),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_643),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_647),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_635),
.A2(n_425),
.B1(n_610),
.B2(n_477),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_671),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_SL g775 ( 
.A(n_735),
.B(n_421),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_655),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_655),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_665),
.Y(n_778)
);

OA21x2_ASAP7_75t_L g779 ( 
.A1(n_754),
.A2(n_498),
.B(n_380),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_650),
.B(n_630),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_671),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_665),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_630),
.B(n_474),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_672),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_651),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_651),
.B(n_709),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_674),
.A2(n_477),
.B1(n_610),
.B2(n_425),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_709),
.B(n_474),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_687),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_754),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_671),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_755),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_761),
.A2(n_629),
.B1(n_451),
.B2(n_576),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_687),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_736),
.B(n_496),
.Y(n_795)
);

CKINVDCx11_ASAP7_75t_R g796 ( 
.A(n_700),
.Y(n_796)
);

OA21x2_ASAP7_75t_L g797 ( 
.A1(n_755),
.A2(n_498),
.B(n_380),
.Y(n_797)
);

BUFx12f_ASAP7_75t_L g798 ( 
.A(n_694),
.Y(n_798)
);

AND2x6_ASAP7_75t_L g799 ( 
.A(n_650),
.B(n_380),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_756),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_650),
.B(n_514),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_641),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_653),
.B(n_496),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_673),
.B(n_576),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_650),
.B(n_514),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_692),
.Y(n_806)
);

INVxp33_ASAP7_75t_SL g807 ( 
.A(n_658),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_671),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_756),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_736),
.B(n_471),
.Y(n_810)
);

INVx6_ASAP7_75t_L g811 ( 
.A(n_667),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_632),
.B(n_633),
.Y(n_812)
);

NOR2x1_ASAP7_75t_L g813 ( 
.A(n_632),
.B(n_558),
.Y(n_813)
);

BUFx8_ASAP7_75t_L g814 ( 
.A(n_645),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_638),
.A2(n_629),
.B1(n_381),
.B2(n_385),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_692),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_645),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_682),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_675),
.A2(n_461),
.B1(n_499),
.B2(n_452),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_633),
.B(n_512),
.Y(n_820)
);

AOI22x1_ASAP7_75t_L g821 ( 
.A1(n_634),
.A2(n_357),
.B1(n_376),
.B2(n_349),
.Y(n_821)
);

CKINVDCx6p67_ASAP7_75t_R g822 ( 
.A(n_740),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_757),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_693),
.Y(n_824)
);

OA21x2_ASAP7_75t_L g825 ( 
.A1(n_757),
.A2(n_760),
.B(n_758),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_758),
.Y(n_826)
);

OA21x2_ASAP7_75t_L g827 ( 
.A1(n_760),
.A2(n_598),
.B(n_498),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_653),
.B(n_367),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_714),
.Y(n_829)
);

CKINVDCx6p67_ASAP7_75t_R g830 ( 
.A(n_648),
.Y(n_830)
);

OA21x2_ASAP7_75t_L g831 ( 
.A1(n_762),
.A2(n_598),
.B(n_376),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_714),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_695),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_751),
.A2(n_598),
.B(n_383),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_762),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_751),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_763),
.Y(n_837)
);

INVxp33_ASAP7_75t_L g838 ( 
.A(n_657),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_699),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_763),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_764),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_670),
.B(n_367),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_671),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_667),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_764),
.A2(n_383),
.B(n_357),
.Y(n_845)
);

OA21x2_ASAP7_75t_L g846 ( 
.A1(n_765),
.A2(n_394),
.B(n_389),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_634),
.B(n_472),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_706),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_765),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_766),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_766),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_L g852 ( 
.A(n_707),
.B(n_514),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_637),
.B(n_639),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_667),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_743),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_743),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_667),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_637),
.B(n_741),
.Y(n_858)
);

AND2x2_ASAP7_75t_SL g859 ( 
.A(n_639),
.B(n_435),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_642),
.B(n_472),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_744),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_SL g862 ( 
.A1(n_715),
.A2(n_382),
.B1(n_392),
.B2(n_387),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_667),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_642),
.B(n_514),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_744),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_667),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_667),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_745),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_745),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_667),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_644),
.B(n_519),
.Y(n_871)
);

OA21x2_ASAP7_75t_L g872 ( 
.A1(n_644),
.A2(n_394),
.B(n_389),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_646),
.B(n_336),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_701),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_748),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_670),
.B(n_367),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_646),
.A2(n_397),
.B(n_396),
.Y(n_877)
);

OA21x2_ASAP7_75t_L g878 ( 
.A1(n_652),
.A2(n_397),
.B(n_396),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_748),
.Y(n_879)
);

BUFx8_ASAP7_75t_L g880 ( 
.A(n_631),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_652),
.B(n_347),
.Y(n_881)
);

OA21x2_ASAP7_75t_L g882 ( 
.A1(n_654),
.A2(n_411),
.B(n_400),
.Y(n_882)
);

OA21x2_ASAP7_75t_L g883 ( 
.A1(n_654),
.A2(n_411),
.B(n_400),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_750),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_702),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_750),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_660),
.B(n_514),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_697),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_676),
.B(n_367),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_752),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_861),
.Y(n_891)
);

NOR2xp67_ASAP7_75t_L g892 ( 
.A(n_798),
.B(n_711),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_796),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_861),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_818),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_818),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_798),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_798),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_861),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_825),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_780),
.B(n_640),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_861),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_848),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_785),
.B(n_649),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_770),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_804),
.A2(n_769),
.B1(n_767),
.B2(n_803),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_814),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_861),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_772),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_R g910 ( 
.A(n_822),
.B(n_661),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_R g911 ( 
.A(n_822),
.B(n_659),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_R g912 ( 
.A(n_822),
.B(n_713),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_824),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_807),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_825),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_830),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_861),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_824),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_830),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_817),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_848),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_830),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_814),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_814),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_814),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_880),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_880),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_824),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_817),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_880),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_833),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_880),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_862),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_793),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_865),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_793),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_862),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_802),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_833),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_802),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_888),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_812),
.B(n_710),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_767),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_865),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_888),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_833),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_839),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_R g948 ( 
.A(n_775),
.B(n_721),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_769),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_785),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_815),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_815),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_839),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_839),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_865),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_874),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_874),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_825),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_874),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_885),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_785),
.B(n_717),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_885),
.Y(n_962)
);

CKINVDCx16_ASAP7_75t_R g963 ( 
.A(n_775),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_R g964 ( 
.A(n_852),
.B(n_722),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_885),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_810),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_810),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_773),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_855),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_773),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_889),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_803),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_811),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_825),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_889),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_787),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_786),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_787),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_865),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_855),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_865),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_828),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_819),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_819),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_783),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_783),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_825),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_R g988 ( 
.A(n_788),
.B(n_734),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_856),
.Y(n_989)
);

BUFx10_ASAP7_75t_L g990 ( 
.A(n_780),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_851),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_788),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_856),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_869),
.Y(n_994)
);

NOR2x1p5_ASAP7_75t_L g995 ( 
.A(n_828),
.B(n_746),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_869),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_884),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_R g998 ( 
.A(n_795),
.B(n_753),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_842),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_L g1000 ( 
.A(n_799),
.B(n_547),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_851),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_795),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_842),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_851),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_812),
.B(n_858),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_876),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_876),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_780),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_780),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_859),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_820),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_768),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_786),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_884),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_873),
.B(n_696),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_820),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_847),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_847),
.Y(n_1018)
);

AOI21x1_ASAP7_75t_L g1019 ( 
.A1(n_845),
.A2(n_662),
.B(n_660),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_865),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_860),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_860),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_812),
.B(n_759),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_871),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_871),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_873),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_881),
.Y(n_1027)
);

NOR2xp67_ASAP7_75t_L g1028 ( 
.A(n_853),
.B(n_680),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_881),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_868),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_868),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_886),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_868),
.Y(n_1033)
);

AND2x6_ASAP7_75t_L g1034 ( 
.A(n_801),
.B(n_558),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_859),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_768),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_811),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_859),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_886),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_812),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_768),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_858),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_858),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_858),
.Y(n_1044)
);

NAND2xp33_ASAP7_75t_R g1045 ( 
.A(n_846),
.B(n_698),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_799),
.B(n_737),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_890),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_771),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_811),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_821),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_821),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_771),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_811),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_771),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_799),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_853),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_811),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_799),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_799),
.Y(n_1059)
);

INVxp67_ASAP7_75t_SL g1060 ( 
.A(n_854),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_838),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1017),
.B(n_799),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_990),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_990),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1005),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1005),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1012),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_1055),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_969),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_980),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_989),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_1055),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1018),
.B(n_799),
.Y(n_1073)
);

AND2x6_ASAP7_75t_L g1074 ( 
.A(n_900),
.B(n_801),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1021),
.B(n_1016),
.Y(n_1075)
);

INVxp67_ASAP7_75t_L g1076 ( 
.A(n_941),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_993),
.Y(n_1077)
);

INVx6_ASAP7_75t_L g1078 ( 
.A(n_990),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_994),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_902),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_996),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_903),
.B(n_921),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_997),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1024),
.B(n_684),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1012),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_966),
.B(n_799),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_985),
.B(n_703),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_985),
.B(n_728),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_967),
.B(n_799),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_902),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_902),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1022),
.B(n_801),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_895),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1014),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_902),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_905),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_1058),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1032),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_905),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_909),
.Y(n_1100)
);

INVx4_ASAP7_75t_L g1101 ( 
.A(n_1058),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_909),
.Y(n_1102)
);

OR2x2_ASAP7_75t_SL g1103 ( 
.A(n_963),
.B(n_719),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_902),
.Y(n_1104)
);

NOR2x1p5_ASAP7_75t_L g1105 ( 
.A(n_897),
.B(n_404),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1026),
.B(n_844),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_986),
.B(n_801),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1040),
.A2(n_805),
.B1(n_749),
.B2(n_401),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_1061),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_986),
.B(n_805),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1039),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_992),
.B(n_805),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1047),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_992),
.B(n_805),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_901),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_1002),
.B(n_844),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1002),
.B(n_813),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_901),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_SL g1119 ( 
.A1(n_983),
.A2(n_720),
.B1(n_739),
.B2(n_724),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_942),
.B(n_864),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_901),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_942),
.B(n_864),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1036),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1027),
.B(n_1029),
.Y(n_1124)
);

INVx4_ASAP7_75t_L g1125 ( 
.A(n_1059),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1003),
.B(n_685),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1040),
.A2(n_813),
.B1(n_887),
.B2(n_864),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_945),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_955),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_913),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_995),
.B(n_864),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_938),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1003),
.B(n_747),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_914),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_918),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_977),
.B(n_844),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1015),
.B(n_887),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1006),
.B(n_704),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_955),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_1059),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_896),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1036),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1041),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_906),
.B(n_1050),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_928),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_931),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1034),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1013),
.B(n_887),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1050),
.B(n_844),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1041),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1028),
.B(n_887),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_940),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1006),
.B(n_718),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1042),
.B(n_716),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1007),
.B(n_971),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1034),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_943),
.B(n_890),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1008),
.B(n_854),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_939),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_949),
.B(n_854),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_946),
.Y(n_1161)
);

OAI221xp5_ASAP7_75t_L g1162 ( 
.A1(n_983),
.A2(n_430),
.B1(n_439),
.B2(n_419),
.C(n_418),
.Y(n_1162)
);

OR2x6_ASAP7_75t_L g1163 ( 
.A(n_892),
.B(n_872),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1048),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_904),
.B(n_857),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_947),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1048),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1008),
.B(n_857),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_953),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1034),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_960),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1009),
.B(n_857),
.Y(n_1172)
);

BUFx4f_ASAP7_75t_L g1173 ( 
.A(n_1034),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_950),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_920),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1007),
.B(n_666),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_961),
.B(n_863),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_965),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_991),
.Y(n_1179)
);

OAI22xp33_ASAP7_75t_SL g1180 ( 
.A1(n_976),
.A2(n_403),
.B1(n_407),
.B2(n_393),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1051),
.B(n_863),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1009),
.B(n_1042),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_L g1183 ( 
.A(n_1043),
.B(n_863),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_914),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_897),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_973),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1043),
.B(n_662),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_955),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_955),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1051),
.B(n_866),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_991),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1052),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1044),
.B(n_663),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1001),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1054),
.Y(n_1195)
);

CKINVDCx16_ASAP7_75t_R g1196 ( 
.A(n_910),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1001),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_893),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_975),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1054),
.Y(n_1200)
);

BUFx4f_ASAP7_75t_L g1201 ( 
.A(n_1034),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_954),
.B(n_866),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1004),
.Y(n_1203)
);

INVx8_ASAP7_75t_L g1204 ( 
.A(n_1034),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1044),
.B(n_866),
.Y(n_1205)
);

BUFx10_ASAP7_75t_L g1206 ( 
.A(n_898),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_956),
.B(n_867),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_984),
.A2(n_878),
.B1(n_882),
.B2(n_872),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_929),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_957),
.B(n_870),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1004),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_959),
.B(n_870),
.Y(n_1212)
);

INVx5_ASAP7_75t_L g1213 ( 
.A(n_981),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1023),
.B(n_663),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1046),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1025),
.B(n_679),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_915),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_958),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_948),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_898),
.Y(n_1220)
);

NAND2xp33_ASAP7_75t_SL g1221 ( 
.A(n_988),
.B(n_664),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1011),
.B(n_679),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_962),
.B(n_870),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_891),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_981),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_981),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1010),
.B(n_664),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_982),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1010),
.B(n_408),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_1056),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1035),
.B(n_666),
.Y(n_1231)
);

AO22x2_ASAP7_75t_L g1232 ( 
.A1(n_968),
.A2(n_970),
.B1(n_978),
.B2(n_976),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_891),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_981),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1035),
.B(n_668),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_891),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_894),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1038),
.B(n_413),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_894),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1037),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_894),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_972),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_951),
.B(n_668),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_998),
.B(n_877),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_899),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1038),
.B(n_669),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_952),
.B(n_669),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_950),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1063),
.B(n_981),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1243),
.B(n_978),
.Y(n_1250)
);

NAND2x1p5_ASAP7_75t_L g1251 ( 
.A(n_1147),
.B(n_899),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1227),
.B(n_999),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1124),
.B(n_933),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1115),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1231),
.B(n_1031),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1152),
.B(n_924),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1124),
.A2(n_1045),
.B1(n_937),
.B2(n_1033),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1067),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1235),
.B(n_1060),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1246),
.B(n_964),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1137),
.B(n_987),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1118),
.B(n_987),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1121),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1147),
.B(n_916),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1156),
.B(n_1170),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1069),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1106),
.A2(n_1053),
.B(n_1049),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1067),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1082),
.Y(n_1269)
);

INVxp33_ASAP7_75t_L g1270 ( 
.A(n_1132),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1063),
.B(n_1020),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1063),
.B(n_1020),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1247),
.B(n_974),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1144),
.A2(n_936),
.B1(n_934),
.B2(n_911),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1116),
.B(n_912),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1116),
.B(n_899),
.Y(n_1276)
);

AND3x1_ASAP7_75t_L g1277 ( 
.A(n_1133),
.B(n_430),
.C(n_419),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1176),
.B(n_908),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1078),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1187),
.B(n_908),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1187),
.B(n_908),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1085),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1187),
.B(n_917),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1085),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1075),
.B(n_924),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1144),
.B(n_925),
.Y(n_1286)
);

NOR2x1p5_ASAP7_75t_L g1287 ( 
.A(n_1102),
.B(n_1096),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1063),
.B(n_1030),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1070),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1071),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_1078),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1077),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1123),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1079),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1106),
.A2(n_1053),
.B(n_1049),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1229),
.A2(n_916),
.B1(n_922),
.B2(n_919),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1064),
.B(n_1020),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1193),
.B(n_917),
.Y(n_1298)
);

NOR3xp33_ASAP7_75t_L g1299 ( 
.A(n_1087),
.B(n_1088),
.C(n_1182),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1123),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_SL g1301 ( 
.A(n_1196),
.B(n_919),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1096),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1204),
.Y(n_1303)
);

NOR3xp33_ASAP7_75t_L g1304 ( 
.A(n_1087),
.B(n_439),
.C(n_418),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1182),
.B(n_922),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1084),
.B(n_926),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1064),
.B(n_1020),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1193),
.B(n_917),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1088),
.B(n_1107),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1193),
.B(n_935),
.Y(n_1310)
);

AND2x6_ASAP7_75t_SL g1311 ( 
.A(n_1155),
.B(n_446),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1126),
.B(n_927),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1110),
.B(n_935),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1093),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1112),
.B(n_935),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1114),
.B(n_944),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1120),
.B(n_944),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1120),
.B(n_944),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1081),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1156),
.B(n_930),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1120),
.B(n_979),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1204),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1117),
.B(n_979),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1083),
.Y(n_1324)
);

NOR2xp67_ASAP7_75t_L g1325 ( 
.A(n_1219),
.B(n_932),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1064),
.B(n_1020),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1216),
.B(n_907),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1229),
.B(n_979),
.Y(n_1328)
);

NOR2xp67_ASAP7_75t_L g1329 ( 
.A(n_1220),
.B(n_879),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1142),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1122),
.B(n_677),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1141),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1142),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1122),
.B(n_677),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1221),
.A2(n_1000),
.B1(n_1030),
.B2(n_1057),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1122),
.B(n_678),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1143),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_SL g1338 ( 
.A(n_1206),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1094),
.Y(n_1339)
);

NAND2xp33_ASAP7_75t_L g1340 ( 
.A(n_1064),
.B(n_1030),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1143),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1238),
.B(n_1065),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_1170),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1158),
.A2(n_1057),
.B1(n_1030),
.B2(n_429),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1150),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1150),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1136),
.B(n_678),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1102),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1164),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1164),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1136),
.B(n_681),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1092),
.B(n_681),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1238),
.B(n_1030),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1173),
.B(n_1019),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1098),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1232),
.A2(n_923),
.B1(n_482),
.B2(n_398),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1214),
.B(n_683),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1173),
.B(n_877),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1111),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1214),
.B(n_1066),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1157),
.B(n_420),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1222),
.B(n_1138),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1186),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1113),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1153),
.B(n_872),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1167),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1062),
.B(n_432),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1201),
.B(n_1174),
.Y(n_1368)
);

AND2x6_ASAP7_75t_SL g1369 ( 
.A(n_1198),
.B(n_449),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_SL g1370 ( 
.A(n_1206),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1232),
.A2(n_482),
.B1(n_398),
.B2(n_473),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1130),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1073),
.B(n_436),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1201),
.B(n_877),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1214),
.B(n_683),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1158),
.B(n_686),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1168),
.B(n_686),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1076),
.B(n_872),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1109),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1174),
.B(n_868),
.Y(n_1380)
);

AND2x2_ASAP7_75t_SL g1381 ( 
.A(n_1183),
.B(n_878),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1186),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1221),
.A2(n_882),
.B1(n_883),
.B2(n_878),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1168),
.B(n_688),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1068),
.B(n_868),
.Y(n_1385)
);

NAND2x1_ASAP7_75t_L g1386 ( 
.A(n_1078),
.B(n_878),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1198),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1185),
.B(n_473),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1135),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1080),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1086),
.B(n_437),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1149),
.A2(n_845),
.B(n_882),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1145),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_1248),
.Y(n_1394)
);

INVxp33_ASAP7_75t_SL g1395 ( 
.A(n_1134),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1146),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1068),
.B(n_868),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1080),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1167),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1390),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1309),
.A2(n_1162),
.B(n_1172),
.C(n_1244),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1250),
.B(n_1230),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1347),
.A2(n_1183),
.B(n_1244),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1362),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1309),
.B(n_1199),
.Y(n_1405)
);

AOI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1354),
.A2(n_1190),
.B(n_1149),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1351),
.A2(n_1377),
.B(n_1376),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1252),
.B(n_1099),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1384),
.A2(n_1212),
.B(n_1202),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1279),
.Y(n_1410)
);

AO22x1_ASAP7_75t_L g1411 ( 
.A1(n_1253),
.A2(n_1185),
.B1(n_1184),
.B2(n_1134),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1266),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1342),
.B(n_1154),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1342),
.B(n_1099),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1299),
.B(n_1154),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1253),
.B(n_1154),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1304),
.A2(n_1108),
.B(n_1209),
.C(n_1175),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1390),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1265),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1353),
.B(n_1248),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1348),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1361),
.A2(n_1100),
.B(n_1180),
.C(n_1242),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1258),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1361),
.A2(n_1275),
.B(n_1305),
.C(n_1285),
.Y(n_1424)
);

O2A1O1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1305),
.A2(n_1100),
.B(n_1160),
.C(n_1205),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1390),
.Y(n_1426)
);

OAI21xp33_ASAP7_75t_L g1427 ( 
.A1(n_1388),
.A2(n_1184),
.B(n_1172),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1273),
.B(n_1232),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1264),
.B(n_1131),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1258),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1257),
.B(n_1357),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1269),
.B(n_1228),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1306),
.A2(n_1119),
.B1(n_1109),
.B2(n_1131),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1323),
.A2(n_1208),
.B(n_1207),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1276),
.A2(n_1210),
.B(n_1207),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1375),
.B(n_1285),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1312),
.B(n_1089),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1289),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1360),
.B(n_1148),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1290),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1292),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1387),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1302),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1268),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1327),
.B(n_1128),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1268),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1282),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1353),
.A2(n_1223),
.B(n_1210),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1379),
.B(n_1103),
.Y(n_1449)
);

AO21x1_ASAP7_75t_L g1450 ( 
.A1(n_1328),
.A2(n_1190),
.B(n_1223),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1282),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1328),
.A2(n_1177),
.B(n_1165),
.Y(n_1452)
);

A2O1A1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1367),
.A2(n_689),
.B(n_690),
.C(n_688),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1264),
.B(n_1131),
.Y(n_1454)
);

BUFx4f_ASAP7_75t_L g1455 ( 
.A(n_1264),
.Y(n_1455)
);

A2O1A1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1367),
.A2(n_690),
.B(n_691),
.C(n_689),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1314),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1331),
.B(n_1215),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1390),
.Y(n_1459)
);

NOR3xp33_ASAP7_75t_L g1460 ( 
.A(n_1260),
.B(n_1205),
.C(n_445),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1395),
.A2(n_1105),
.B1(n_1206),
.B2(n_1074),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1381),
.B(n_1080),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1398),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1354),
.A2(n_1181),
.B(n_1104),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1358),
.A2(n_1226),
.B(n_1104),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1381),
.B(n_1080),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1334),
.B(n_1151),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1294),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1323),
.A2(n_1074),
.B(n_1159),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1265),
.B(n_1068),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1286),
.B(n_1161),
.Y(n_1471)
);

AOI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1249),
.A2(n_1191),
.B(n_1179),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1319),
.Y(n_1473)
);

OAI21xp33_ASAP7_75t_L g1474 ( 
.A1(n_1278),
.A2(n_444),
.B(n_441),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1286),
.A2(n_1163),
.B1(n_1127),
.B2(n_1166),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1373),
.A2(n_1171),
.B(n_1178),
.C(n_1169),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1358),
.A2(n_1104),
.B(n_1095),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1265),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1336),
.B(n_1217),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1332),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1256),
.B(n_1163),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1255),
.B(n_1217),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1284),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1352),
.B(n_1218),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1302),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1301),
.A2(n_1074),
.B1(n_1097),
.B2(n_1072),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1284),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1424),
.A2(n_1373),
.B(n_1391),
.C(n_1329),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1423),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1452),
.A2(n_1374),
.B(n_1340),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1430),
.Y(n_1491)
);

O2A1O1Ixp5_ASAP7_75t_L g1492 ( 
.A1(n_1401),
.A2(n_1385),
.B(n_1397),
.C(n_1368),
.Y(n_1492)
);

BUFx4f_ASAP7_75t_L g1493 ( 
.A(n_1470),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1405),
.B(n_1296),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1414),
.B(n_1277),
.Y(n_1495)
);

AOI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1403),
.A2(n_1374),
.B(n_1392),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1401),
.A2(n_1339),
.B1(n_1355),
.B2(n_1324),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1407),
.A2(n_1261),
.B(n_1385),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1444),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1455),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1413),
.A2(n_1414),
.B1(n_1436),
.B2(n_1415),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1458),
.B(n_1365),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1400),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1431),
.B(n_1259),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1405),
.B(n_1274),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1409),
.A2(n_1397),
.B(n_1368),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1471),
.B(n_1359),
.Y(n_1507)
);

AO31x2_ASAP7_75t_L g1508 ( 
.A1(n_1450),
.A2(n_1300),
.A3(n_1330),
.B(n_1293),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1427),
.A2(n_1372),
.B(n_1393),
.C(n_1389),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1446),
.Y(n_1510)
);

NOR3xp33_ASAP7_75t_SL g1511 ( 
.A(n_1442),
.B(n_450),
.C(n_448),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1435),
.A2(n_1386),
.B(n_1271),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1464),
.A2(n_1271),
.B(n_1249),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1471),
.B(n_1364),
.Y(n_1514)
);

INVx4_ASAP7_75t_L g1515 ( 
.A(n_1455),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1447),
.Y(n_1516)
);

INVx3_ASAP7_75t_SL g1517 ( 
.A(n_1429),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1404),
.B(n_1378),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1400),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1400),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1428),
.A2(n_1371),
.B1(n_1356),
.B2(n_1391),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1469),
.A2(n_1288),
.B(n_1272),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1481),
.B(n_1254),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1400),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1448),
.A2(n_1288),
.B(n_1272),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1404),
.B(n_1263),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1406),
.A2(n_834),
.B(n_1267),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1429),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1419),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1451),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1416),
.B(n_1425),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1483),
.Y(n_1532)
);

O2A1O1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1453),
.A2(n_1396),
.B(n_1281),
.C(n_1283),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1408),
.B(n_1411),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1408),
.B(n_1270),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1432),
.B(n_1320),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1432),
.B(n_1320),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1419),
.B(n_1398),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1418),
.Y(n_1539)
);

O2A1O1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1453),
.A2(n_1298),
.B(n_1308),
.C(n_1280),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1490),
.A2(n_1466),
.B(n_1462),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1488),
.A2(n_1498),
.B(n_1507),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1499),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1496),
.A2(n_1477),
.B(n_1465),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1514),
.B(n_1412),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1501),
.B(n_1535),
.Y(n_1546)
);

AOI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1496),
.A2(n_1472),
.B(n_1466),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1527),
.A2(n_1462),
.B(n_1434),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1508),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1527),
.A2(n_1512),
.B(n_1513),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1501),
.A2(n_1420),
.B(n_1456),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1494),
.A2(n_1495),
.B1(n_1534),
.B2(n_1505),
.Y(n_1552)
);

AOI21x1_ASAP7_75t_SL g1553 ( 
.A1(n_1518),
.A2(n_1402),
.B(n_1445),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1519),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1504),
.A2(n_1420),
.B(n_1456),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1508),
.Y(n_1556)
);

O2A1O1Ixp33_ASAP7_75t_SL g1557 ( 
.A1(n_1531),
.A2(n_1476),
.B(n_1461),
.C(n_1437),
.Y(n_1557)
);

NOR4xp25_ASAP7_75t_L g1558 ( 
.A(n_1521),
.B(n_1422),
.C(n_443),
.D(n_446),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1504),
.A2(n_1307),
.B(n_1297),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1525),
.A2(n_834),
.B(n_1295),
.Y(n_1560)
);

OA21x2_ASAP7_75t_L g1561 ( 
.A1(n_1522),
.A2(n_834),
.B(n_1482),
.Y(n_1561)
);

AOI211x1_ASAP7_75t_L g1562 ( 
.A1(n_1526),
.A2(n_443),
.B(n_449),
.C(n_445),
.Y(n_1562)
);

NAND2x1_ASAP7_75t_L g1563 ( 
.A(n_1503),
.B(n_1418),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1536),
.A2(n_1437),
.B1(n_1433),
.B2(n_1417),
.Y(n_1564)
);

AO31x2_ASAP7_75t_L g1565 ( 
.A1(n_1497),
.A2(n_1484),
.A3(n_1487),
.B(n_1479),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1508),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1492),
.A2(n_1460),
.B(n_1506),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1537),
.B(n_1311),
.Y(n_1568)
);

AO31x2_ASAP7_75t_L g1569 ( 
.A1(n_1497),
.A2(n_1293),
.A3(n_1330),
.B(n_1300),
.Y(n_1569)
);

AO31x2_ASAP7_75t_L g1570 ( 
.A1(n_1489),
.A2(n_1337),
.A3(n_1341),
.B(n_1333),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1503),
.A2(n_1307),
.B(n_1297),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1502),
.A2(n_1326),
.B(n_1467),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1523),
.B(n_1438),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1503),
.A2(n_1326),
.B(n_1380),
.Y(n_1574)
);

AO31x2_ASAP7_75t_L g1575 ( 
.A1(n_1489),
.A2(n_1510),
.A3(n_1516),
.B(n_1491),
.Y(n_1575)
);

BUFx12f_ASAP7_75t_L g1576 ( 
.A(n_1500),
.Y(n_1576)
);

OAI21x1_ASAP7_75t_L g1577 ( 
.A1(n_1524),
.A2(n_1380),
.B(n_845),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1529),
.B(n_1440),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1508),
.Y(n_1579)
);

BUFx8_ASAP7_75t_L g1580 ( 
.A(n_1500),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1529),
.B(n_1441),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1523),
.B(n_1468),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1519),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1538),
.B(n_1478),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1493),
.B(n_1475),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1528),
.B(n_1421),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1519),
.Y(n_1587)
);

OA21x2_ASAP7_75t_L g1588 ( 
.A1(n_1502),
.A2(n_1383),
.B(n_1315),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1511),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1509),
.A2(n_1460),
.B(n_1344),
.Y(n_1590)
);

AOI21xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1546),
.A2(n_1517),
.B(n_456),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1576),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1554),
.B(n_1524),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1578),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1568),
.A2(n_1449),
.B1(n_1499),
.B2(n_1491),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1557),
.A2(n_1564),
.B(n_1552),
.C(n_1590),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1550),
.A2(n_1544),
.B(n_1542),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1554),
.B(n_1524),
.Y(n_1598)
);

INVx6_ASAP7_75t_L g1599 ( 
.A(n_1580),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1554),
.B(n_1519),
.Y(n_1600)
);

INVx5_ASAP7_75t_L g1601 ( 
.A(n_1576),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_SL g1602 ( 
.A1(n_1586),
.A2(n_456),
.B(n_480),
.C(n_459),
.Y(n_1602)
);

AO31x2_ASAP7_75t_L g1603 ( 
.A1(n_1549),
.A2(n_1516),
.A3(n_1530),
.B(n_1510),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1578),
.B(n_1508),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1575),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1550),
.A2(n_1532),
.B(n_1530),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1589),
.A2(n_1517),
.B1(n_1485),
.B2(n_453),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1544),
.A2(n_1540),
.B(n_1533),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1581),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1575),
.Y(n_1610)
);

AOI21xp33_ASAP7_75t_L g1611 ( 
.A1(n_1585),
.A2(n_1163),
.B(n_1474),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1547),
.A2(n_1532),
.B(n_1470),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1551),
.A2(n_1493),
.B(n_1519),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1581),
.B(n_1520),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1583),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1547),
.A2(n_1560),
.B(n_1548),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1575),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1575),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1543),
.A2(n_1439),
.B1(n_1454),
.B2(n_1457),
.Y(n_1619)
);

INVx4_ASAP7_75t_L g1620 ( 
.A(n_1583),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1556),
.B(n_1520),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1556),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1575),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1570),
.Y(n_1624)
);

OA21x2_ASAP7_75t_L g1625 ( 
.A1(n_1548),
.A2(n_752),
.B(n_705),
.Y(n_1625)
);

INVx2_ASAP7_75t_SL g1626 ( 
.A(n_1583),
.Y(n_1626)
);

CKINVDCx6p67_ASAP7_75t_R g1627 ( 
.A(n_1545),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_SL g1628 ( 
.A1(n_1567),
.A2(n_1515),
.B(n_1486),
.Y(n_1628)
);

AND2x4_ASAP7_75t_SL g1629 ( 
.A(n_1584),
.B(n_1500),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1566),
.A2(n_1316),
.B(n_1313),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1570),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1573),
.B(n_1480),
.Y(n_1632)
);

OR2x6_ASAP7_75t_L g1633 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1633)
);

AOI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1558),
.A2(n_475),
.B1(n_480),
.B2(n_459),
.C(n_453),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1589),
.B(n_1443),
.Y(n_1635)
);

INVx4_ASAP7_75t_SL g1636 ( 
.A(n_1569),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1587),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_SL g1638 ( 
.A1(n_1572),
.A2(n_1515),
.B(n_1528),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1566),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1555),
.A2(n_1325),
.B(n_1493),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1560),
.A2(n_1337),
.B(n_1333),
.Y(n_1641)
);

O2A1O1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1559),
.A2(n_475),
.B(n_501),
.C(n_483),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1562),
.A2(n_1517),
.B1(n_1528),
.B2(n_1287),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_L g1644 ( 
.A(n_1582),
.B(n_1480),
.C(n_536),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1584),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1579),
.A2(n_705),
.B(n_691),
.Y(n_1646)
);

BUFx12f_ASAP7_75t_L g1647 ( 
.A(n_1580),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1584),
.A2(n_1454),
.B1(n_1500),
.B2(n_1320),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1574),
.A2(n_1345),
.B(n_1341),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1580),
.Y(n_1650)
);

OAI222xp33_ASAP7_75t_L g1651 ( 
.A1(n_1579),
.A2(n_1473),
.B1(n_522),
.B2(n_501),
.C1(n_524),
.C2(n_511),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1565),
.B(n_1520),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1587),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_SL g1654 ( 
.A1(n_1541),
.A2(n_1410),
.B(n_1310),
.Y(n_1654)
);

AOI22x1_ASAP7_75t_L g1655 ( 
.A1(n_1587),
.A2(n_1410),
.B1(n_511),
.B2(n_522),
.Y(n_1655)
);

O2A1O1Ixp33_ASAP7_75t_SL g1656 ( 
.A1(n_1563),
.A2(n_524),
.B(n_525),
.C(n_483),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1574),
.A2(n_1346),
.B(n_1345),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1571),
.A2(n_1349),
.B(n_1346),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1588),
.A2(n_1457),
.B1(n_1350),
.B2(n_1366),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1571),
.A2(n_1350),
.B(n_1349),
.Y(n_1660)
);

NOR2x1_ASAP7_75t_SL g1661 ( 
.A(n_1553),
.B(n_1500),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1565),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1577),
.A2(n_1394),
.B(n_712),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1563),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1570),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_R g1666 ( 
.A(n_1565),
.B(n_1279),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1577),
.A2(n_1399),
.B(n_1366),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1570),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1565),
.B(n_1538),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1569),
.B(n_1520),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1569),
.Y(n_1671)
);

A2O1A1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1588),
.A2(n_712),
.B(n_725),
.C(n_708),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1588),
.B(n_1538),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1561),
.A2(n_1399),
.B1(n_473),
.B2(n_596),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1569),
.B(n_1539),
.Y(n_1675)
);

AO31x2_ASAP7_75t_L g1676 ( 
.A1(n_1671),
.A2(n_1569),
.A3(n_879),
.B(n_1570),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1596),
.A2(n_1561),
.B(n_1539),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_SL g1678 ( 
.A1(n_1646),
.A2(n_1369),
.B1(n_482),
.B2(n_398),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1597),
.A2(n_1561),
.B(n_1188),
.Y(n_1679)
);

OR2x6_ASAP7_75t_L g1680 ( 
.A(n_1633),
.B(n_1539),
.Y(n_1680)
);

A2O1A1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1591),
.A2(n_528),
.B(n_531),
.C(n_525),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1622),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1613),
.A2(n_1539),
.B(n_1398),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1632),
.B(n_528),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1622),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1639),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1666),
.A2(n_1539),
.B(n_1398),
.Y(n_1687)
);

AND2x6_ASAP7_75t_L g1688 ( 
.A(n_1652),
.B(n_1670),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1627),
.B(n_531),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1597),
.A2(n_1188),
.B(n_1095),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1639),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1616),
.A2(n_1188),
.B(n_1095),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1594),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1594),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1591),
.A2(n_622),
.B(n_549),
.Y(n_1695)
);

OAI21x1_ASAP7_75t_SL g1696 ( 
.A1(n_1661),
.A2(n_549),
.B(n_536),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1627),
.B(n_567),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1666),
.A2(n_1343),
.B(n_1418),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1616),
.A2(n_1226),
.B(n_1189),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1605),
.Y(n_1700)
);

AO21x2_ASAP7_75t_L g1701 ( 
.A1(n_1671),
.A2(n_723),
.B(n_879),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1614),
.B(n_1538),
.Y(n_1702)
);

INVxp67_ASAP7_75t_SL g1703 ( 
.A(n_1662),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1609),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1614),
.B(n_567),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1609),
.B(n_1418),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1604),
.B(n_577),
.Y(n_1707)
);

OAI21x1_ASAP7_75t_L g1708 ( 
.A1(n_1608),
.A2(n_1226),
.B(n_1189),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1604),
.Y(n_1709)
);

NAND2x1p5_ASAP7_75t_L g1710 ( 
.A(n_1601),
.B(n_1426),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1645),
.B(n_1593),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1593),
.B(n_577),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1652),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1593),
.B(n_582),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1637),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1654),
.A2(n_1459),
.B(n_1426),
.Y(n_1716)
);

AO31x2_ASAP7_75t_L g1717 ( 
.A1(n_1662),
.A2(n_1631),
.A3(n_1668),
.B(n_1624),
.Y(n_1717)
);

OAI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1608),
.A2(n_1189),
.B(n_1363),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1654),
.A2(n_1459),
.B(n_1426),
.Y(n_1719)
);

AO31x2_ASAP7_75t_L g1720 ( 
.A1(n_1624),
.A2(n_792),
.A3(n_800),
.B(n_790),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1628),
.A2(n_1459),
.B(n_1426),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1655),
.A2(n_1370),
.B1(n_1338),
.B2(n_582),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1605),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1669),
.B(n_708),
.Y(n_1724)
);

AO21x2_ASAP7_75t_L g1725 ( 
.A1(n_1630),
.A2(n_1668),
.B(n_1631),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1673),
.B(n_725),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1640),
.B(n_585),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1621),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1621),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1603),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1647),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1603),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1637),
.B(n_585),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1603),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1675),
.B(n_726),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1653),
.B(n_593),
.Y(n_1736)
);

BUFx5_ASAP7_75t_L g1737 ( 
.A(n_1670),
.Y(n_1737)
);

AOI21x1_ASAP7_75t_L g1738 ( 
.A1(n_1646),
.A2(n_727),
.B(n_726),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1603),
.Y(n_1739)
);

AO31x2_ASAP7_75t_L g1740 ( 
.A1(n_1610),
.A2(n_792),
.A3(n_800),
.B(n_790),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1603),
.Y(n_1741)
);

OAI21x1_ASAP7_75t_L g1742 ( 
.A1(n_1628),
.A2(n_1382),
.B(n_1363),
.Y(n_1742)
);

AO31x2_ASAP7_75t_L g1743 ( 
.A1(n_1610),
.A2(n_823),
.A3(n_826),
.B(n_809),
.Y(n_1743)
);

BUFx12f_ASAP7_75t_L g1744 ( 
.A(n_1647),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1606),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1638),
.A2(n_1463),
.B(n_1459),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1606),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1598),
.B(n_593),
.Y(n_1748)
);

CKINVDCx8_ASAP7_75t_R g1749 ( 
.A(n_1635),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1653),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1598),
.B(n_605),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1598),
.B(n_605),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1661),
.B(n_612),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1664),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1664),
.Y(n_1755)
);

INVx4_ASAP7_75t_L g1756 ( 
.A(n_1599),
.Y(n_1756)
);

OAI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1641),
.A2(n_1382),
.B(n_1262),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1617),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1606),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1606),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1617),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1618),
.Y(n_1762)
);

OAI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1642),
.A2(n_613),
.B(n_612),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1675),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1646),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1626),
.B(n_727),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1623),
.Y(n_1767)
);

A2O1A1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1634),
.A2(n_621),
.B(n_622),
.C(n_613),
.Y(n_1768)
);

BUFx2_ASAP7_75t_R g1769 ( 
.A(n_1650),
.Y(n_1769)
);

AOI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1646),
.A2(n_730),
.B(n_729),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1650),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1625),
.Y(n_1772)
);

AO21x2_ASAP7_75t_L g1773 ( 
.A1(n_1630),
.A2(n_730),
.B(n_729),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1623),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1620),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1625),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1670),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1626),
.Y(n_1778)
);

INVx6_ASAP7_75t_L g1779 ( 
.A(n_1601),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1615),
.Y(n_1780)
);

OAI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1602),
.A2(n_621),
.B(n_731),
.Y(n_1781)
);

OAI21x1_ASAP7_75t_L g1782 ( 
.A1(n_1641),
.A2(n_1478),
.B(n_1203),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1615),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1665),
.Y(n_1784)
);

AO21x2_ASAP7_75t_L g1785 ( 
.A1(n_1630),
.A2(n_732),
.B(n_731),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1643),
.B(n_1),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1615),
.B(n_1463),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1665),
.Y(n_1788)
);

OA21x2_ASAP7_75t_L g1789 ( 
.A1(n_1612),
.A2(n_733),
.B(n_732),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1644),
.B(n_1),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1600),
.B(n_1463),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1620),
.B(n_2),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1612),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1633),
.B(n_1463),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1633),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1600),
.B(n_733),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1633),
.Y(n_1797)
);

OA21x2_ASAP7_75t_L g1798 ( 
.A1(n_1658),
.A2(n_741),
.B(n_738),
.Y(n_1798)
);

OAI21x1_ASAP7_75t_L g1799 ( 
.A1(n_1667),
.A2(n_1203),
.B(n_1197),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1651),
.A2(n_454),
.B1(n_458),
.B2(n_457),
.C(n_455),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1620),
.Y(n_1801)
);

AO21x2_ASAP7_75t_L g1802 ( 
.A1(n_1611),
.A2(n_742),
.B(n_738),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1636),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1638),
.A2(n_1213),
.B(n_1097),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1600),
.B(n_742),
.Y(n_1805)
);

OAI21x1_ASAP7_75t_L g1806 ( 
.A1(n_1667),
.A2(n_1211),
.B(n_1194),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1636),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1672),
.A2(n_465),
.B(n_460),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1592),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1656),
.A2(n_467),
.B(n_466),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1592),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1636),
.Y(n_1812)
);

INVx6_ASAP7_75t_L g1813 ( 
.A(n_1601),
.Y(n_1813)
);

OAI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1649),
.A2(n_1251),
.B(n_1192),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1663),
.A2(n_1213),
.B(n_1097),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1636),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1629),
.B(n_547),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1658),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1649),
.A2(n_1251),
.B(n_1192),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1625),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1625),
.A2(n_1213),
.B(n_1101),
.Y(n_1821)
);

AO21x2_ASAP7_75t_L g1822 ( 
.A1(n_1660),
.A2(n_823),
.B(n_809),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1660),
.Y(n_1823)
);

AOI21x1_ASAP7_75t_L g1824 ( 
.A1(n_1657),
.A2(n_835),
.B(n_826),
.Y(n_1824)
);

AOI21x1_ASAP7_75t_L g1825 ( 
.A1(n_1745),
.A2(n_1657),
.B(n_841),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1713),
.B(n_1601),
.Y(n_1826)
);

HB1xp67_ASAP7_75t_L g1827 ( 
.A(n_1704),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1755),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1700),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1713),
.B(n_1601),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1700),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1723),
.Y(n_1832)
);

AOI21x1_ASAP7_75t_L g1833 ( 
.A1(n_1745),
.A2(n_841),
.B(n_835),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1682),
.Y(n_1834)
);

NAND3xp33_ASAP7_75t_L g1835 ( 
.A(n_1727),
.B(n_1595),
.C(n_1674),
.Y(n_1835)
);

AO21x2_ASAP7_75t_L g1836 ( 
.A1(n_1747),
.A2(n_1648),
.B(n_778),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1728),
.B(n_1599),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1682),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1685),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1723),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1705),
.B(n_1659),
.Y(n_1841)
);

OR2x6_ASAP7_75t_L g1842 ( 
.A(n_1680),
.B(n_1599),
.Y(n_1842)
);

NOR2x1p5_ASAP7_75t_L g1843 ( 
.A(n_1744),
.B(n_1592),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1758),
.Y(n_1844)
);

OAI222xp33_ASAP7_75t_L g1845 ( 
.A1(n_1678),
.A2(n_1619),
.B1(n_1655),
.B2(n_484),
.C1(n_469),
.C2(n_486),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1704),
.Y(n_1846)
);

AO21x2_ASAP7_75t_L g1847 ( 
.A1(n_1759),
.A2(n_778),
.B(n_777),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1686),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1758),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1709),
.B(n_1592),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1769),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1761),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1733),
.B(n_1592),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1761),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1715),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1691),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1762),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1764),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1729),
.B(n_1599),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1755),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1703),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1762),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1703),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1688),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1715),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1693),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1702),
.B(n_1629),
.Y(n_1867)
);

OR2x2_ASAP7_75t_SL g1868 ( 
.A(n_1707),
.B(n_1724),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1688),
.B(n_547),
.Y(n_1869)
);

INVx1_ASAP7_75t_SL g1870 ( 
.A(n_1731),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1694),
.Y(n_1871)
);

INVx1_ASAP7_75t_SL g1872 ( 
.A(n_1771),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1727),
.A2(n_470),
.B(n_468),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1774),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1750),
.B(n_547),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1736),
.Y(n_1876)
);

BUFx2_ASAP7_75t_L g1877 ( 
.A(n_1754),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1767),
.Y(n_1878)
);

OA21x2_ASAP7_75t_L g1879 ( 
.A1(n_1760),
.A2(n_1732),
.B(n_1730),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1780),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1783),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1778),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1740),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1717),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1740),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1688),
.B(n_547),
.Y(n_1886)
);

BUFx3_ASAP7_75t_L g1887 ( 
.A(n_1749),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1712),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1714),
.Y(n_1889)
);

INVx3_ASAP7_75t_L g1890 ( 
.A(n_1688),
.Y(n_1890)
);

INVx4_ASAP7_75t_L g1891 ( 
.A(n_1811),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1711),
.B(n_547),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1809),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1748),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1775),
.Y(n_1895)
);

INVx2_ASAP7_75t_SL g1896 ( 
.A(n_1779),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1717),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1751),
.Y(n_1898)
);

OR2x6_ASAP7_75t_L g1899 ( 
.A(n_1680),
.B(n_1607),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1735),
.B(n_2),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1752),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1717),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1689),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1726),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1777),
.B(n_1688),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1777),
.B(n_3),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1795),
.B(n_5),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1737),
.B(n_6),
.Y(n_1908)
);

OR2x6_ASAP7_75t_L g1909 ( 
.A(n_1680),
.B(n_1291),
.Y(n_1909)
);

OAI21x1_ASAP7_75t_L g1910 ( 
.A1(n_1708),
.A2(n_1200),
.B(n_1195),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1801),
.Y(n_1911)
);

INVx2_ASAP7_75t_SL g1912 ( 
.A(n_1779),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1797),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1740),
.Y(n_1914)
);

OAI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1681),
.A2(n_488),
.B(n_487),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1740),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1743),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1765),
.B(n_7),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1737),
.B(n_10),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1743),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1743),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1756),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1717),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1734),
.Y(n_1924)
);

OAI21x1_ASAP7_75t_L g1925 ( 
.A1(n_1679),
.A2(n_1718),
.B(n_1677),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1684),
.B(n_11),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1739),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1805),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1741),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1743),
.Y(n_1930)
);

OA21x2_ASAP7_75t_L g1931 ( 
.A1(n_1677),
.A2(n_778),
.B(n_777),
.Y(n_1931)
);

INVx8_ASAP7_75t_L g1932 ( 
.A(n_1794),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1720),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1725),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1725),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1737),
.Y(n_1936)
);

OR2x6_ASAP7_75t_L g1937 ( 
.A(n_1698),
.B(n_1291),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1720),
.Y(n_1938)
);

INVxp67_ASAP7_75t_L g1939 ( 
.A(n_1697),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1737),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1720),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1737),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1737),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1784),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1807),
.B(n_11),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1720),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1676),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1676),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1796),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1772),
.B(n_1776),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1792),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1676),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1676),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1772),
.B(n_12),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1784),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1773),
.Y(n_1956)
);

NAND3xp33_ASAP7_75t_L g1957 ( 
.A(n_1753),
.B(n_875),
.C(n_495),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1788),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1793),
.Y(n_1959)
);

AO21x2_ASAP7_75t_L g1960 ( 
.A1(n_1773),
.A2(n_784),
.B(n_777),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1756),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1785),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1785),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1776),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1820),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1706),
.B(n_13),
.Y(n_1966)
);

NAND2x1_ASAP7_75t_L g1967 ( 
.A(n_1779),
.B(n_435),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1818),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1823),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1812),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1706),
.B(n_15),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1816),
.Y(n_1972)
);

BUFx2_ASAP7_75t_L g1973 ( 
.A(n_1813),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1766),
.B(n_15),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1792),
.B(n_490),
.Y(n_1975)
);

OAI21x1_ASAP7_75t_L g1976 ( 
.A1(n_1698),
.A2(n_1200),
.B(n_1195),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1789),
.Y(n_1977)
);

INVx2_ASAP7_75t_SL g1978 ( 
.A(n_1813),
.Y(n_1978)
);

AOI21x1_ASAP7_75t_L g1979 ( 
.A1(n_1967),
.A2(n_1770),
.B(n_1738),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1951),
.A2(n_1786),
.B1(n_1681),
.B2(n_1678),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1967),
.Y(n_1981)
);

OA21x2_ASAP7_75t_L g1982 ( 
.A1(n_1964),
.A2(n_1803),
.B(n_1687),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1835),
.A2(n_1841),
.B1(n_1903),
.B2(n_1802),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1877),
.B(n_1787),
.Y(n_1984)
);

INVx3_ASAP7_75t_L g1985 ( 
.A(n_1864),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1839),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1864),
.B(n_1794),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1950),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1869),
.A2(n_1802),
.B1(n_1786),
.B2(n_1790),
.Y(n_1989)
);

AOI211xp5_ASAP7_75t_L g1990 ( 
.A1(n_1954),
.A2(n_1790),
.B(n_1753),
.C(n_1695),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1944),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1950),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1861),
.Y(n_1993)
);

AOI222xp33_ASAP7_75t_L g1994 ( 
.A1(n_1873),
.A2(n_1763),
.B1(n_1800),
.B2(n_1808),
.C1(n_1768),
.C2(n_1810),
.Y(n_1994)
);

OAI22xp33_ASAP7_75t_SL g1995 ( 
.A1(n_1954),
.A2(n_1813),
.B1(n_1687),
.B2(n_1722),
.Y(n_1995)
);

INVx2_ASAP7_75t_SL g1996 ( 
.A(n_1887),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1839),
.Y(n_1997)
);

OA21x2_ASAP7_75t_L g1998 ( 
.A1(n_1964),
.A2(n_1683),
.B(n_1692),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1944),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1869),
.A2(n_1701),
.B1(n_1696),
.B2(n_1817),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1955),
.Y(n_2001)
);

INVx4_ASAP7_75t_L g2002 ( 
.A(n_1887),
.Y(n_2002)
);

OAI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1899),
.A2(n_1815),
.B1(n_1683),
.B2(n_1781),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1949),
.B(n_1791),
.Y(n_2004)
);

INVxp67_ASAP7_75t_L g2005 ( 
.A(n_1877),
.Y(n_2005)
);

AOI21xp33_ASAP7_75t_L g2006 ( 
.A1(n_1918),
.A2(n_1789),
.B(n_1768),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1864),
.B(n_1710),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1869),
.A2(n_1789),
.B1(n_1798),
.B2(n_1822),
.Y(n_2008)
);

OAI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1899),
.A2(n_1815),
.B1(n_1721),
.B2(n_1821),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1890),
.B(n_1721),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1892),
.B(n_1716),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1890),
.B(n_1710),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1955),
.Y(n_2013)
);

AOI221xp5_ASAP7_75t_L g2014 ( 
.A1(n_1975),
.A2(n_497),
.B1(n_506),
.B2(n_504),
.C(n_503),
.Y(n_2014)
);

AOI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1886),
.A2(n_1798),
.B1(n_1822),
.B2(n_596),
.Y(n_2015)
);

OAI221xp5_ASAP7_75t_L g2016 ( 
.A1(n_1926),
.A2(n_508),
.B1(n_515),
.B2(n_513),
.C(n_510),
.Y(n_2016)
);

AOI22xp33_ASAP7_75t_SL g2017 ( 
.A1(n_1908),
.A2(n_1798),
.B1(n_482),
.B2(n_398),
.Y(n_2017)
);

OA21x2_ASAP7_75t_L g2018 ( 
.A1(n_1884),
.A2(n_1699),
.B(n_1690),
.Y(n_2018)
);

BUFx12f_ASAP7_75t_L g2019 ( 
.A(n_1926),
.Y(n_2019)
);

AOI22xp33_ASAP7_75t_SL g2020 ( 
.A1(n_1908),
.A2(n_1821),
.B1(n_1370),
.B2(n_1338),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1858),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1937),
.A2(n_1719),
.B(n_1716),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1958),
.Y(n_2023)
);

AOI31xp33_ASAP7_75t_L g2024 ( 
.A1(n_1851),
.A2(n_1746),
.A3(n_1719),
.B(n_1804),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_1886),
.A2(n_596),
.B1(n_875),
.B2(n_794),
.Y(n_2025)
);

OAI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1899),
.A2(n_1868),
.B1(n_1945),
.B2(n_1918),
.Y(n_2026)
);

OAI221xp5_ASAP7_75t_L g2027 ( 
.A1(n_1915),
.A2(n_517),
.B1(n_521),
.B2(n_520),
.C(n_518),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1858),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1892),
.B(n_1746),
.Y(n_2029)
);

AOI221xp5_ASAP7_75t_SL g2030 ( 
.A1(n_1872),
.A2(n_1804),
.B1(n_19),
.B2(n_17),
.C(n_18),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1870),
.Y(n_2031)
);

OA21x2_ASAP7_75t_L g2032 ( 
.A1(n_1884),
.A2(n_1757),
.B(n_1782),
.Y(n_2032)
);

AOI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1937),
.A2(n_1742),
.B(n_1806),
.Y(n_2033)
);

AOI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_1886),
.A2(n_596),
.B1(n_875),
.B2(n_794),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1961),
.Y(n_2035)
);

INVxp67_ASAP7_75t_L g2036 ( 
.A(n_1875),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1958),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1834),
.Y(n_2038)
);

AOI21xp33_ASAP7_75t_L g2039 ( 
.A1(n_1970),
.A2(n_533),
.B(n_527),
.Y(n_2039)
);

OAI221xp5_ASAP7_75t_L g2040 ( 
.A1(n_1900),
.A2(n_534),
.B1(n_539),
.B2(n_538),
.C(n_537),
.Y(n_2040)
);

NAND3xp33_ASAP7_75t_L g2041 ( 
.A(n_1970),
.B(n_1972),
.C(n_1838),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1904),
.A2(n_1939),
.B1(n_1888),
.B2(n_1894),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_1889),
.A2(n_875),
.B1(n_794),
.B2(n_806),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1875),
.Y(n_2044)
);

OAI211xp5_ASAP7_75t_L g2045 ( 
.A1(n_1919),
.A2(n_541),
.B(n_542),
.C(n_540),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1890),
.B(n_1824),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1834),
.Y(n_2047)
);

OR2x6_ASAP7_75t_L g2048 ( 
.A(n_1937),
.B(n_1909),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_SL g2049 ( 
.A1(n_1919),
.A2(n_544),
.B1(n_546),
.B2(n_543),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1838),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1848),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1876),
.B(n_1799),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1898),
.B(n_548),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1826),
.Y(n_2054)
);

AOI211xp5_ASAP7_75t_L g2055 ( 
.A1(n_1845),
.A2(n_553),
.B(n_555),
.C(n_550),
.Y(n_2055)
);

AOI221xp5_ASAP7_75t_L g2056 ( 
.A1(n_1901),
.A2(n_559),
.B1(n_565),
.B2(n_564),
.C(n_563),
.Y(n_2056)
);

AOI222xp33_ASAP7_75t_L g2057 ( 
.A1(n_1957),
.A2(n_569),
.B1(n_573),
.B2(n_579),
.C1(n_578),
.C2(n_566),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1956),
.A2(n_875),
.B1(n_806),
.B2(n_816),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1856),
.Y(n_2059)
);

AOI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_1956),
.A2(n_875),
.B1(n_806),
.B2(n_816),
.Y(n_2060)
);

OR2x6_ASAP7_75t_L g2061 ( 
.A(n_1937),
.B(n_1814),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_SL g2062 ( 
.A1(n_1900),
.A2(n_586),
.B1(n_587),
.B2(n_580),
.Y(n_2062)
);

OAI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1899),
.A2(n_589),
.B1(n_592),
.B2(n_588),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1962),
.A2(n_1963),
.B1(n_1972),
.B2(n_1836),
.Y(n_2064)
);

AOI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_1945),
.A2(n_883),
.B1(n_882),
.B2(n_597),
.Y(n_2065)
);

NAND3xp33_ASAP7_75t_L g2066 ( 
.A(n_1882),
.B(n_599),
.C(n_594),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1895),
.B(n_1819),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1880),
.Y(n_2068)
);

OAI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1974),
.A2(n_602),
.B1(n_603),
.B2(n_600),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_1962),
.A2(n_816),
.B1(n_829),
.B2(n_789),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1829),
.Y(n_2071)
);

AO21x2_ASAP7_75t_L g2072 ( 
.A1(n_1934),
.A2(n_832),
.B(n_829),
.Y(n_2072)
);

OAI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_1868),
.A2(n_606),
.B1(n_607),
.B2(n_604),
.Y(n_2073)
);

OR2x6_ASAP7_75t_L g2074 ( 
.A(n_1909),
.B(n_1303),
.Y(n_2074)
);

OA21x2_ASAP7_75t_L g2075 ( 
.A1(n_1897),
.A2(n_609),
.B(n_608),
.Y(n_2075)
);

OAI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_1974),
.A2(n_620),
.B1(n_623),
.B2(n_611),
.Y(n_2076)
);

AOI22xp33_ASAP7_75t_L g2077 ( 
.A1(n_1963),
.A2(n_1836),
.B1(n_1913),
.B2(n_1914),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_1861),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_1836),
.A2(n_1917),
.B1(n_1920),
.B2(n_1916),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1880),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_1843),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_1921),
.A2(n_832),
.B1(n_836),
.B2(n_829),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1881),
.Y(n_2083)
);

OAI22xp33_ASAP7_75t_L g2084 ( 
.A1(n_1907),
.A2(n_626),
.B1(n_627),
.B2(n_624),
.Y(n_2084)
);

AOI222xp33_ASAP7_75t_L g2085 ( 
.A1(n_1906),
.A2(n_628),
.B1(n_442),
.B2(n_435),
.C1(n_836),
.C2(n_832),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1829),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1866),
.B(n_1882),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1895),
.B(n_20),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1866),
.B(n_20),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1837),
.B(n_21),
.Y(n_2090)
);

OAI22xp33_ASAP7_75t_L g2091 ( 
.A1(n_1907),
.A2(n_442),
.B1(n_435),
.B2(n_1335),
.Y(n_2091)
);

OAI222xp33_ASAP7_75t_L g2092 ( 
.A1(n_1928),
.A2(n_356),
.B1(n_351),
.B2(n_359),
.C1(n_355),
.C2(n_348),
.Y(n_2092)
);

INVx3_ASAP7_75t_L g2093 ( 
.A(n_1826),
.Y(n_2093)
);

OAI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_1945),
.A2(n_1317),
.B1(n_1321),
.B2(n_1318),
.Y(n_2094)
);

OAI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1961),
.A2(n_883),
.B1(n_442),
.B2(n_435),
.Y(n_2095)
);

OAI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_1853),
.A2(n_883),
.B1(n_442),
.B2(n_1224),
.Y(n_2096)
);

AOI221xp5_ASAP7_75t_L g2097 ( 
.A1(n_1863),
.A2(n_442),
.B1(n_364),
.B2(n_365),
.C(n_362),
.Y(n_2097)
);

AOI22xp33_ASAP7_75t_L g2098 ( 
.A1(n_1930),
.A2(n_837),
.B1(n_840),
.B2(n_836),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_1827),
.B(n_21),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_SL g2100 ( 
.A1(n_1906),
.A2(n_442),
.B1(n_883),
.B2(n_368),
.Y(n_2100)
);

BUFx4f_ASAP7_75t_SL g2101 ( 
.A(n_1891),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_1905),
.A2(n_782),
.B1(n_776),
.B2(n_831),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_1933),
.A2(n_837),
.B1(n_840),
.B2(n_831),
.Y(n_2103)
);

INVx1_ASAP7_75t_SL g2104 ( 
.A(n_1893),
.Y(n_2104)
);

AOI221xp5_ASAP7_75t_L g2105 ( 
.A1(n_1863),
.A2(n_378),
.B1(n_384),
.B2(n_377),
.C(n_360),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1881),
.Y(n_2106)
);

INVx3_ASAP7_75t_L g2107 ( 
.A(n_1826),
.Y(n_2107)
);

OAI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_1893),
.A2(n_1236),
.B1(n_1237),
.B2(n_1233),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1871),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_1938),
.A2(n_837),
.B1(n_840),
.B2(n_831),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_1909),
.A2(n_1241),
.B1(n_1245),
.B2(n_1239),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_1931),
.A2(n_1213),
.B(n_1091),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1968),
.Y(n_2113)
);

INVx5_ASAP7_75t_SL g2114 ( 
.A(n_1909),
.Y(n_2114)
);

OAI22xp5_ASAP7_75t_L g2115 ( 
.A1(n_1830),
.A2(n_402),
.B1(n_410),
.B2(n_388),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1968),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_1941),
.A2(n_831),
.B1(n_850),
.B2(n_849),
.Y(n_2117)
);

OAI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_1966),
.A2(n_1971),
.B(n_1911),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_1846),
.B(n_22),
.Y(n_2119)
);

BUFx3_ASAP7_75t_L g2120 ( 
.A(n_1966),
.Y(n_2120)
);

BUFx2_ASAP7_75t_L g2121 ( 
.A(n_1891),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1837),
.B(n_22),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_1946),
.A2(n_831),
.B1(n_850),
.B2(n_849),
.Y(n_2123)
);

BUFx2_ASAP7_75t_L g2124 ( 
.A(n_1891),
.Y(n_2124)
);

OAI21xp33_ASAP7_75t_L g2125 ( 
.A1(n_1865),
.A2(n_782),
.B(n_776),
.Y(n_2125)
);

OAI21x1_ASAP7_75t_L g2126 ( 
.A1(n_1925),
.A2(n_782),
.B(n_776),
.Y(n_2126)
);

OAI22xp33_ASAP7_75t_L g2127 ( 
.A1(n_1842),
.A2(n_417),
.B1(n_422),
.B2(n_412),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1831),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_1883),
.A2(n_850),
.B1(n_849),
.B2(n_782),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1831),
.Y(n_2130)
);

AOI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_1931),
.A2(n_1091),
.B(n_1090),
.Y(n_2131)
);

AOI21xp33_ASAP7_75t_L g2132 ( 
.A1(n_1969),
.A2(n_23),
.B(n_24),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_1932),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1969),
.Y(n_2134)
);

HB1xp67_ASAP7_75t_L g2135 ( 
.A(n_1855),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1832),
.Y(n_2136)
);

OAI21x1_ASAP7_75t_L g2137 ( 
.A1(n_1925),
.A2(n_776),
.B(n_846),
.Y(n_2137)
);

AOI221xp5_ASAP7_75t_L g2138 ( 
.A1(n_1965),
.A2(n_433),
.B1(n_434),
.B2(n_426),
.C(n_424),
.Y(n_2138)
);

AOI221xp5_ASAP7_75t_L g2139 ( 
.A1(n_1965),
.A2(n_476),
.B1(n_478),
.B2(n_463),
.C(n_447),
.Y(n_2139)
);

NAND2x1_ASAP7_75t_L g2140 ( 
.A(n_1985),
.B(n_1830),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1986),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1997),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1982),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2036),
.B(n_1865),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2036),
.B(n_1850),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_2135),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2054),
.B(n_1828),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2109),
.B(n_1959),
.Y(n_2148)
);

HB1xp67_ASAP7_75t_L g2149 ( 
.A(n_2135),
.Y(n_2149)
);

INVxp67_ASAP7_75t_SL g2150 ( 
.A(n_1993),
.Y(n_2150)
);

BUFx2_ASAP7_75t_L g2151 ( 
.A(n_2002),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2087),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1984),
.B(n_1859),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1987),
.B(n_1859),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1987),
.B(n_1828),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2120),
.B(n_1828),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2031),
.B(n_1860),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2054),
.B(n_2093),
.Y(n_2158)
);

NOR2x1_ASAP7_75t_L g2159 ( 
.A(n_2002),
.B(n_1860),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2093),
.B(n_1860),
.Y(n_2160)
);

INVx4_ASAP7_75t_L g2161 ( 
.A(n_2101),
.Y(n_2161)
);

AND2x4_ASAP7_75t_L g2162 ( 
.A(n_2048),
.B(n_1830),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2021),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_1988),
.B(n_1850),
.Y(n_2164)
);

CKINVDCx14_ASAP7_75t_R g2165 ( 
.A(n_2063),
.Y(n_2165)
);

INVx2_ASAP7_75t_SL g2166 ( 
.A(n_1985),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2028),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2113),
.Y(n_2168)
);

OR2x2_ASAP7_75t_L g2169 ( 
.A(n_1988),
.B(n_1959),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2029),
.B(n_1971),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2107),
.B(n_1973),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_2044),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2011),
.B(n_1867),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2044),
.B(n_1867),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2107),
.B(n_1973),
.Y(n_2175)
);

OAI222xp33_ASAP7_75t_L g2176 ( 
.A1(n_1983),
.A2(n_2026),
.B1(n_2073),
.B2(n_1980),
.C1(n_1989),
.C2(n_2017),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_1992),
.B(n_1896),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1992),
.B(n_1922),
.Y(n_2178)
);

INVx5_ASAP7_75t_L g2179 ( 
.A(n_2048),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2044),
.B(n_1936),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1982),
.Y(n_2181)
);

OR2x2_ASAP7_75t_L g2182 ( 
.A(n_2004),
.B(n_1896),
.Y(n_2182)
);

OR2x2_ASAP7_75t_L g2183 ( 
.A(n_2005),
.B(n_1978),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2005),
.B(n_1936),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2121),
.B(n_1922),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2007),
.B(n_1922),
.Y(n_2186)
);

OAI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_2003),
.A2(n_1942),
.B(n_1940),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2051),
.B(n_1940),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2012),
.B(n_1912),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2038),
.B(n_2047),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2071),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2086),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2116),
.Y(n_2193)
);

AND2x4_ASAP7_75t_SL g2194 ( 
.A(n_2048),
.B(n_1842),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_1993),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2124),
.B(n_1912),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2134),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2081),
.B(n_1978),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2068),
.Y(n_2199)
);

AND2x4_ASAP7_75t_L g2200 ( 
.A(n_2010),
.B(n_2061),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_1996),
.B(n_1932),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2080),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2118),
.B(n_1905),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2128),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2067),
.B(n_1942),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2083),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2059),
.B(n_1943),
.Y(n_2207)
);

OAI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_2003),
.A2(n_1990),
.B1(n_2020),
.B2(n_2024),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2130),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2106),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2010),
.B(n_1943),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2136),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2050),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2089),
.B(n_1879),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2099),
.B(n_2119),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2041),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2078),
.B(n_1842),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1991),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2078),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2104),
.B(n_1842),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2052),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_2035),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1999),
.Y(n_2223)
);

AOI22xp33_ASAP7_75t_L g2224 ( 
.A1(n_1994),
.A2(n_1977),
.B1(n_1931),
.B2(n_1883),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_2061),
.B(n_1947),
.Y(n_2225)
);

INVxp67_ASAP7_75t_SL g2226 ( 
.A(n_1995),
.Y(n_2226)
);

OR2x2_ASAP7_75t_L g2227 ( 
.A(n_2042),
.B(n_1879),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2133),
.B(n_1932),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2090),
.B(n_1932),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_2061),
.B(n_1947),
.Y(n_2230)
);

INVx1_ASAP7_75t_SL g2231 ( 
.A(n_2019),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2001),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2013),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2023),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2088),
.B(n_2122),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_2114),
.B(n_1879),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2046),
.B(n_1924),
.Y(n_2237)
);

INVx5_ASAP7_75t_L g2238 ( 
.A(n_2074),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2030),
.B(n_1924),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2037),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2053),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2114),
.B(n_1998),
.Y(n_2242)
);

AND2x4_ASAP7_75t_L g2243 ( 
.A(n_2074),
.B(n_1948),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2009),
.B(n_1927),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1998),
.Y(n_2245)
);

OR2x2_ASAP7_75t_L g2246 ( 
.A(n_2114),
.B(n_1927),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2020),
.B(n_1929),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2075),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_2018),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2074),
.B(n_1929),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_SL g2251 ( 
.A1(n_2062),
.A2(n_1977),
.B1(n_1885),
.B2(n_1902),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2075),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2062),
.B(n_2069),
.Y(n_2253)
);

NAND2x1p5_ASAP7_75t_L g2254 ( 
.A(n_1981),
.B(n_1976),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_1981),
.Y(n_2255)
);

OR2x2_ASAP7_75t_L g2256 ( 
.A(n_2064),
.B(n_1885),
.Y(n_2256)
);

HB1xp67_ASAP7_75t_L g2257 ( 
.A(n_2018),
.Y(n_2257)
);

AND2x4_ASAP7_75t_L g2258 ( 
.A(n_2022),
.B(n_1948),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2032),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2076),
.B(n_1833),
.Y(n_2260)
);

BUFx2_ASAP7_75t_L g2261 ( 
.A(n_1981),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2022),
.B(n_1833),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2033),
.B(n_1825),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2032),
.Y(n_2264)
);

AO22x1_ASAP7_75t_L g2265 ( 
.A1(n_2094),
.A2(n_1953),
.B1(n_1952),
.B2(n_1902),
.Y(n_2265)
);

AND2x4_ASAP7_75t_SL g2266 ( 
.A(n_2220),
.B(n_2000),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2141),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2142),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2163),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2167),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2168),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2203),
.B(n_2049),
.Y(n_2272)
);

NAND2xp67_ASAP7_75t_L g2273 ( 
.A(n_2242),
.B(n_2033),
.Y(n_2273)
);

OAI21xp33_ASAP7_75t_L g2274 ( 
.A1(n_2226),
.A2(n_2049),
.B(n_2132),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2203),
.B(n_2039),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2143),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2198),
.B(n_2115),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2220),
.B(n_2126),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2193),
.Y(n_2279)
);

INVx2_ASAP7_75t_SL g2280 ( 
.A(n_2157),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2197),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2199),
.Y(n_2282)
);

OR2x2_ASAP7_75t_L g2283 ( 
.A(n_2144),
.B(n_2040),
.Y(n_2283)
);

INVx4_ASAP7_75t_L g2284 ( 
.A(n_2161),
.Y(n_2284)
);

OAI221xp5_ASAP7_75t_SL g2285 ( 
.A1(n_2226),
.A2(n_2045),
.B1(n_2016),
.B2(n_2040),
.C(n_2027),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2158),
.B(n_2077),
.Y(n_2286)
);

INVx4_ASAP7_75t_L g2287 ( 
.A(n_2161),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2216),
.B(n_2084),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_2238),
.B(n_2066),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2202),
.Y(n_2290)
);

AND2x4_ASAP7_75t_L g2291 ( 
.A(n_2238),
.B(n_2079),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_2208),
.B(n_2017),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2206),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2178),
.B(n_2008),
.Y(n_2294)
);

INVxp67_ASAP7_75t_L g2295 ( 
.A(n_2151),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2178),
.B(n_2006),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2210),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2143),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2171),
.B(n_2015),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2239),
.B(n_2125),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2171),
.B(n_2102),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2213),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2152),
.B(n_2016),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2190),
.Y(n_2304)
);

OR2x2_ASAP7_75t_L g2305 ( 
.A(n_2145),
.B(n_2096),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2175),
.B(n_2155),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2170),
.B(n_2127),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2181),
.Y(n_2308)
);

OA21x2_ASAP7_75t_L g2309 ( 
.A1(n_2245),
.A2(n_1935),
.B(n_1923),
.Y(n_2309)
);

NAND2x1p5_ASAP7_75t_L g2310 ( 
.A(n_2179),
.B(n_1976),
.Y(n_2310)
);

NAND2x1_ASAP7_75t_L g2311 ( 
.A(n_2159),
.B(n_1952),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2181),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2154),
.B(n_2196),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2259),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2264),
.Y(n_2315)
);

AND2x4_ASAP7_75t_SL g2316 ( 
.A(n_2229),
.B(n_2065),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2146),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2185),
.B(n_2108),
.Y(n_2318)
);

HB1xp67_ASAP7_75t_L g2319 ( 
.A(n_2195),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2146),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2241),
.B(n_2127),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2149),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2149),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2195),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2219),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2164),
.B(n_1953),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2185),
.B(n_2137),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2148),
.Y(n_2328)
);

AOI22xp33_ASAP7_75t_L g2329 ( 
.A1(n_2165),
.A2(n_2027),
.B1(n_2097),
.B2(n_2138),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2175),
.B(n_1825),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2147),
.B(n_2045),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2249),
.Y(n_2332)
);

AND2x4_ASAP7_75t_L g2333 ( 
.A(n_2238),
.B(n_1897),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2150),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2150),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_2238),
.B(n_1923),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2249),
.Y(n_2337)
);

AND2x4_ASAP7_75t_L g2338 ( 
.A(n_2162),
.B(n_1979),
.Y(n_2338)
);

INVxp67_ASAP7_75t_L g2339 ( 
.A(n_2260),
.Y(n_2339)
);

NAND3xp33_ASAP7_75t_L g2340 ( 
.A(n_2224),
.B(n_2056),
.C(n_2097),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_2156),
.B(n_2111),
.Y(n_2341)
);

NAND3xp33_ASAP7_75t_L g2342 ( 
.A(n_2224),
.B(n_2056),
.C(n_2014),
.Y(n_2342)
);

BUFx2_ASAP7_75t_L g2343 ( 
.A(n_2161),
.Y(n_2343)
);

OR2x2_ASAP7_75t_L g2344 ( 
.A(n_2173),
.B(n_1832),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2248),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2179),
.B(n_2138),
.Y(n_2346)
);

INVx4_ASAP7_75t_L g2347 ( 
.A(n_2222),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2214),
.B(n_2139),
.Y(n_2348)
);

HB1xp67_ASAP7_75t_L g2349 ( 
.A(n_2221),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2252),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2257),
.Y(n_2351)
);

OR2x2_ASAP7_75t_L g2352 ( 
.A(n_2215),
.B(n_1840),
.Y(n_2352)
);

AND2x4_ASAP7_75t_L g2353 ( 
.A(n_2162),
.B(n_1935),
.Y(n_2353)
);

OR2x2_ASAP7_75t_L g2354 ( 
.A(n_2177),
.B(n_1840),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2147),
.B(n_2129),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2257),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2160),
.B(n_2100),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2169),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2186),
.B(n_2100),
.Y(n_2359)
);

OR2x2_ASAP7_75t_L g2360 ( 
.A(n_2183),
.B(n_1844),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_2162),
.B(n_1844),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2237),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2189),
.B(n_1849),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2153),
.B(n_1849),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2188),
.Y(n_2365)
);

OR2x2_ASAP7_75t_L g2366 ( 
.A(n_2244),
.B(n_2182),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2207),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2262),
.B(n_2139),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2262),
.B(n_2085),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2217),
.B(n_2095),
.Y(n_2370)
);

BUFx2_ASAP7_75t_L g2371 ( 
.A(n_2222),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2232),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2233),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2217),
.B(n_1852),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2237),
.Y(n_2375)
);

HB1xp67_ASAP7_75t_L g2376 ( 
.A(n_2184),
.Y(n_2376)
);

INVx6_ASAP7_75t_L g2377 ( 
.A(n_2179),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2234),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2309),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2313),
.B(n_2228),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_SL g2381 ( 
.A1(n_2368),
.A2(n_2165),
.B1(n_2251),
.B2(n_2227),
.Y(n_2381)
);

INVx4_ASAP7_75t_L g2382 ( 
.A(n_2284),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2348),
.B(n_2272),
.Y(n_2383)
);

OAI33xp33_ASAP7_75t_L g2384 ( 
.A1(n_2292),
.A2(n_2253),
.A3(n_2256),
.B1(n_2235),
.B2(n_2176),
.B3(n_2236),
.Y(n_2384)
);

AND2x4_ASAP7_75t_L g2385 ( 
.A(n_2280),
.B(n_2200),
.Y(n_2385)
);

AOI221xp5_ASAP7_75t_L g2386 ( 
.A1(n_2339),
.A2(n_2014),
.B1(n_2263),
.B2(n_2258),
.C(n_2242),
.Y(n_2386)
);

AND2x4_ASAP7_75t_SL g2387 ( 
.A(n_2331),
.B(n_2201),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_2338),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2319),
.Y(n_2389)
);

OAI33xp33_ASAP7_75t_L g2390 ( 
.A1(n_2292),
.A2(n_2180),
.A3(n_2246),
.B1(n_2240),
.B2(n_2174),
.B3(n_2091),
.Y(n_2390)
);

AND2x4_ASAP7_75t_L g2391 ( 
.A(n_2280),
.B(n_2200),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2331),
.B(n_2201),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2318),
.B(n_2231),
.Y(n_2393)
);

NAND2x1p5_ASAP7_75t_L g2394 ( 
.A(n_2289),
.B(n_2179),
.Y(n_2394)
);

OAI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_2342),
.A2(n_2263),
.B(n_2258),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2332),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2309),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2347),
.B(n_2255),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2309),
.Y(n_2399)
);

AOI21xp5_ASAP7_75t_L g2400 ( 
.A1(n_2274),
.A2(n_2265),
.B(n_2247),
.Y(n_2400)
);

AOI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_2340),
.A2(n_2247),
.B1(n_2258),
.B2(n_2105),
.Y(n_2401)
);

AOI22xp33_ASAP7_75t_L g2402 ( 
.A1(n_2369),
.A2(n_2105),
.B1(n_2057),
.B2(n_2225),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2319),
.Y(n_2403)
);

INVx2_ASAP7_75t_SL g2404 ( 
.A(n_2371),
.Y(n_2404)
);

INVxp67_ASAP7_75t_SL g2405 ( 
.A(n_2321),
.Y(n_2405)
);

OAI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2307),
.A2(n_2172),
.B1(n_2261),
.B2(n_2200),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2345),
.Y(n_2407)
);

OAI221xp5_ASAP7_75t_L g2408 ( 
.A1(n_2339),
.A2(n_2187),
.B1(n_2055),
.B2(n_2250),
.C(n_2205),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2306),
.B(n_2166),
.Y(n_2409)
);

AOI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2283),
.A2(n_2230),
.B1(n_2225),
.B2(n_2243),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2306),
.B(n_2166),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2275),
.B(n_2250),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2296),
.B(n_2211),
.Y(n_2413)
);

INVx3_ASAP7_75t_L g2414 ( 
.A(n_2338),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2350),
.Y(n_2415)
);

NAND3xp33_ASAP7_75t_L g2416 ( 
.A(n_2329),
.B(n_2230),
.C(n_2243),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2267),
.Y(n_2417)
);

OAI33xp33_ASAP7_75t_L g2418 ( 
.A1(n_2295),
.A2(n_2204),
.A3(n_2191),
.B1(n_2212),
.B2(n_2209),
.B3(n_2192),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2362),
.Y(n_2419)
);

NAND3xp33_ASAP7_75t_L g2420 ( 
.A(n_2285),
.B(n_2230),
.C(n_2243),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2362),
.Y(n_2421)
);

INVx4_ASAP7_75t_L g2422 ( 
.A(n_2284),
.Y(n_2422)
);

AOI22xp33_ASAP7_75t_L g2423 ( 
.A1(n_2288),
.A2(n_2300),
.B1(n_2303),
.B2(n_2346),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2375),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2299),
.B(n_2205),
.Y(n_2425)
);

OAI33xp33_ASAP7_75t_L g2426 ( 
.A1(n_2295),
.A2(n_2204),
.A3(n_2191),
.B1(n_2212),
.B2(n_2209),
.B3(n_2192),
.Y(n_2426)
);

OAI221xp5_ASAP7_75t_L g2427 ( 
.A1(n_2346),
.A2(n_2370),
.B1(n_2351),
.B2(n_2356),
.C(n_2337),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2375),
.Y(n_2428)
);

OAI221xp5_ASAP7_75t_L g2429 ( 
.A1(n_2332),
.A2(n_2223),
.B1(n_2218),
.B2(n_2211),
.C(n_2254),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2268),
.Y(n_2430)
);

INVx5_ASAP7_75t_L g2431 ( 
.A(n_2284),
.Y(n_2431)
);

BUFx2_ASAP7_75t_L g2432 ( 
.A(n_2343),
.Y(n_2432)
);

OAI21x1_ASAP7_75t_L g2433 ( 
.A1(n_2276),
.A2(n_2140),
.B(n_2218),
.Y(n_2433)
);

NAND3xp33_ASAP7_75t_L g2434 ( 
.A(n_2317),
.B(n_2034),
.C(n_2025),
.Y(n_2434)
);

NAND4xp25_ASAP7_75t_L g2435 ( 
.A(n_2287),
.B(n_2043),
.C(n_2112),
.D(n_2060),
.Y(n_2435)
);

INVx1_ASAP7_75t_SL g2436 ( 
.A(n_2277),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_2347),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2299),
.B(n_2223),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2296),
.B(n_2194),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2269),
.Y(n_2440)
);

BUFx2_ASAP7_75t_L g2441 ( 
.A(n_2287),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2294),
.B(n_2194),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2304),
.B(n_2254),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2294),
.B(n_1852),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2270),
.Y(n_2445)
);

OR2x2_ASAP7_75t_L g2446 ( 
.A(n_2358),
.B(n_1854),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2337),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2271),
.Y(n_2448)
);

NOR2xp67_ASAP7_75t_SL g2449 ( 
.A(n_2287),
.B(n_2112),
.Y(n_2449)
);

OR2x2_ASAP7_75t_L g2450 ( 
.A(n_2328),
.B(n_1854),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2279),
.Y(n_2451)
);

OR2x2_ASAP7_75t_L g2452 ( 
.A(n_2366),
.B(n_1857),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2281),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2351),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2282),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2355),
.B(n_2376),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2356),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2290),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2276),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_2341),
.B(n_1857),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2355),
.B(n_1862),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2293),
.Y(n_2462)
);

AOI221xp5_ASAP7_75t_L g2463 ( 
.A1(n_2314),
.A2(n_2092),
.B1(n_2131),
.B2(n_2123),
.C(n_2117),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2297),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2376),
.B(n_1862),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2392),
.B(n_2330),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2436),
.B(n_2357),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2456),
.B(n_2357),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2396),
.Y(n_2469)
);

AOI211x1_ASAP7_75t_L g2470 ( 
.A1(n_2427),
.A2(n_2286),
.B(n_2322),
.C(n_2320),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2379),
.Y(n_2471)
);

OR2x2_ASAP7_75t_L g2472 ( 
.A(n_2425),
.B(n_2323),
.Y(n_2472)
);

OR2x2_ASAP7_75t_L g2473 ( 
.A(n_2456),
.B(n_2324),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2380),
.B(n_2330),
.Y(n_2474)
);

AOI31xp33_ASAP7_75t_SL g2475 ( 
.A1(n_2386),
.A2(n_2314),
.A3(n_2315),
.B(n_2305),
.Y(n_2475)
);

INVx3_ASAP7_75t_SL g2476 ( 
.A(n_2437),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2396),
.Y(n_2477)
);

NAND4xp25_ASAP7_75t_L g2478 ( 
.A(n_2398),
.B(n_2347),
.C(n_2335),
.D(n_2334),
.Y(n_2478)
);

OR2x2_ASAP7_75t_L g2479 ( 
.A(n_2419),
.B(n_2325),
.Y(n_2479)
);

INVx3_ASAP7_75t_L g2480 ( 
.A(n_2388),
.Y(n_2480)
);

AOI22xp33_ASAP7_75t_L g2481 ( 
.A1(n_2384),
.A2(n_2291),
.B1(n_2266),
.B2(n_2298),
.Y(n_2481)
);

BUFx3_ASAP7_75t_L g2482 ( 
.A(n_2437),
.Y(n_2482)
);

O2A1O1Ixp33_ASAP7_75t_L g2483 ( 
.A1(n_2395),
.A2(n_2289),
.B(n_2349),
.C(n_2291),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2447),
.Y(n_2484)
);

AND2x4_ASAP7_75t_L g2485 ( 
.A(n_2404),
.B(n_2289),
.Y(n_2485)
);

NOR2x1_ASAP7_75t_L g2486 ( 
.A(n_2382),
.B(n_2315),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2447),
.Y(n_2487)
);

BUFx2_ASAP7_75t_L g2488 ( 
.A(n_2393),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2401),
.B(n_2402),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2387),
.B(n_2338),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2454),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2387),
.B(n_2365),
.Y(n_2492)
);

AOI211xp5_ASAP7_75t_L g2493 ( 
.A1(n_2400),
.A2(n_2291),
.B(n_2349),
.C(n_2092),
.Y(n_2493)
);

AOI221xp5_ASAP7_75t_L g2494 ( 
.A1(n_2418),
.A2(n_2298),
.B1(n_2312),
.B2(n_2308),
.C(n_2286),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2379),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2454),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2397),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2457),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2401),
.B(n_2402),
.Y(n_2499)
);

AOI22xp33_ASAP7_75t_L g2500 ( 
.A1(n_2383),
.A2(n_2266),
.B1(n_2312),
.B2(n_2308),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2397),
.Y(n_2501)
);

OR2x6_ASAP7_75t_L g2502 ( 
.A(n_2394),
.B(n_2377),
.Y(n_2502)
);

NAND2xp33_ASAP7_75t_SL g2503 ( 
.A(n_2404),
.B(n_2302),
.Y(n_2503)
);

AND2x4_ASAP7_75t_L g2504 ( 
.A(n_2385),
.B(n_2367),
.Y(n_2504)
);

HB1xp67_ASAP7_75t_L g2505 ( 
.A(n_2432),
.Y(n_2505)
);

AND2x4_ASAP7_75t_L g2506 ( 
.A(n_2385),
.B(n_2278),
.Y(n_2506)
);

AOI22xp33_ASAP7_75t_L g2507 ( 
.A1(n_2381),
.A2(n_2423),
.B1(n_2390),
.B2(n_2426),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2457),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2407),
.Y(n_2509)
);

INVx6_ASAP7_75t_L g2510 ( 
.A(n_2437),
.Y(n_2510)
);

AOI221xp5_ASAP7_75t_L g2511 ( 
.A1(n_2423),
.A2(n_2359),
.B1(n_2373),
.B2(n_2378),
.C(n_2372),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2415),
.Y(n_2512)
);

INVxp67_ASAP7_75t_SL g2513 ( 
.A(n_2398),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2405),
.B(n_2301),
.Y(n_2514)
);

INVx1_ASAP7_75t_SL g2515 ( 
.A(n_2442),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2438),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2409),
.B(n_2327),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2412),
.B(n_2301),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2409),
.B(n_2311),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2411),
.B(n_2364),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2399),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2385),
.B(n_2361),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2413),
.B(n_2352),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2437),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2389),
.Y(n_2525)
);

INVx1_ASAP7_75t_SL g2526 ( 
.A(n_2442),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2403),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2391),
.B(n_2388),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2391),
.B(n_2361),
.Y(n_2529)
);

AOI21xp33_ASAP7_75t_L g2530 ( 
.A1(n_2419),
.A2(n_2424),
.B(n_2421),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2391),
.B(n_2361),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2388),
.B(n_2363),
.Y(n_2532)
);

BUFx2_ASAP7_75t_L g2533 ( 
.A(n_2441),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2414),
.B(n_2377),
.Y(n_2534)
);

INVx2_ASAP7_75t_SL g2535 ( 
.A(n_2431),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2414),
.B(n_2360),
.Y(n_2536)
);

BUFx3_ASAP7_75t_L g2537 ( 
.A(n_2431),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2421),
.B(n_2344),
.Y(n_2538)
);

HB1xp67_ASAP7_75t_L g2539 ( 
.A(n_2417),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2414),
.B(n_2374),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2399),
.Y(n_2541)
);

BUFx3_ASAP7_75t_L g2542 ( 
.A(n_2431),
.Y(n_2542)
);

OR2x2_ASAP7_75t_L g2543 ( 
.A(n_2424),
.B(n_2326),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2382),
.B(n_2273),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2444),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_L g2546 ( 
.A(n_2382),
.B(n_2354),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_2468),
.B(n_2430),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2471),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2488),
.B(n_2431),
.Y(n_2549)
);

HB1xp67_ASAP7_75t_L g2550 ( 
.A(n_2505),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2471),
.Y(n_2551)
);

OR2x2_ASAP7_75t_L g2552 ( 
.A(n_2473),
.B(n_2440),
.Y(n_2552)
);

OR2x2_ASAP7_75t_L g2553 ( 
.A(n_2473),
.B(n_2445),
.Y(n_2553)
);

OR2x2_ASAP7_75t_L g2554 ( 
.A(n_2467),
.B(n_2448),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2533),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_2470),
.B(n_2394),
.Y(n_2556)
);

HB1xp67_ASAP7_75t_L g2557 ( 
.A(n_2480),
.Y(n_2557)
);

BUFx6f_ASAP7_75t_L g2558 ( 
.A(n_2476),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2485),
.B(n_2422),
.Y(n_2559)
);

INVx1_ASAP7_75t_SL g2560 ( 
.A(n_2515),
.Y(n_2560)
);

AND2x2_ASAP7_75t_SL g2561 ( 
.A(n_2507),
.B(n_2422),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2485),
.B(n_2422),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2495),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2514),
.B(n_2428),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2480),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2495),
.Y(n_2566)
);

OR2x2_ASAP7_75t_L g2567 ( 
.A(n_2518),
.B(n_2451),
.Y(n_2567)
);

OR2x2_ASAP7_75t_L g2568 ( 
.A(n_2526),
.B(n_2472),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2480),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2497),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2497),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2485),
.B(n_2439),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2501),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2513),
.B(n_2428),
.Y(n_2574)
);

OR2x2_ASAP7_75t_L g2575 ( 
.A(n_2472),
.B(n_2453),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2528),
.B(n_2439),
.Y(n_2576)
);

INVx1_ASAP7_75t_SL g2577 ( 
.A(n_2528),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2504),
.B(n_2455),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2501),
.Y(n_2579)
);

NAND2x1_ASAP7_75t_SL g2580 ( 
.A(n_2476),
.B(n_2458),
.Y(n_2580)
);

NAND2x1_ASAP7_75t_L g2581 ( 
.A(n_2502),
.B(n_2406),
.Y(n_2581)
);

OR2x2_ASAP7_75t_L g2582 ( 
.A(n_2523),
.B(n_2462),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2540),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2510),
.B(n_2478),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2520),
.B(n_2464),
.Y(n_2585)
);

BUFx12f_ASAP7_75t_L g2586 ( 
.A(n_2510),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2521),
.Y(n_2587)
);

INVx1_ASAP7_75t_SL g2588 ( 
.A(n_2490),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2504),
.B(n_2460),
.Y(n_2589)
);

NAND2x1p5_ASAP7_75t_L g2590 ( 
.A(n_2482),
.B(n_2449),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2520),
.B(n_2443),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2521),
.Y(n_2592)
);

CKINVDCx16_ASAP7_75t_R g2593 ( 
.A(n_2482),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2522),
.B(n_2410),
.Y(n_2594)
);

NOR2x1_ASAP7_75t_L g2595 ( 
.A(n_2524),
.B(n_2537),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2541),
.Y(n_2596)
);

INVx1_ASAP7_75t_SL g2597 ( 
.A(n_2490),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_L g2598 ( 
.A(n_2510),
.B(n_2408),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2522),
.B(n_2410),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2541),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2540),
.Y(n_2601)
);

INVxp67_ASAP7_75t_L g2602 ( 
.A(n_2534),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2479),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2479),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2545),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2516),
.B(n_2434),
.Y(n_2606)
);

INVxp67_ASAP7_75t_SL g2607 ( 
.A(n_2493),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2550),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2550),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2557),
.Y(n_2610)
);

NAND2x2_ASAP7_75t_L g2611 ( 
.A(n_2581),
.B(n_2524),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2555),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2555),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2557),
.Y(n_2614)
);

OR2x2_ASAP7_75t_L g2615 ( 
.A(n_2568),
.B(n_2469),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2572),
.Y(n_2616)
);

NAND3xp33_ASAP7_75t_L g2617 ( 
.A(n_2556),
.B(n_2511),
.C(n_2499),
.Y(n_2617)
);

INVx2_ASAP7_75t_SL g2618 ( 
.A(n_2572),
.Y(n_2618)
);

OR2x6_ASAP7_75t_L g2619 ( 
.A(n_2558),
.B(n_2489),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2576),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2585),
.Y(n_2621)
);

OR2x2_ASAP7_75t_L g2622 ( 
.A(n_2560),
.B(n_2477),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2576),
.Y(n_2623)
);

INVx1_ASAP7_75t_SL g2624 ( 
.A(n_2580),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2558),
.Y(n_2625)
);

AOI21xp33_ASAP7_75t_L g2626 ( 
.A1(n_2607),
.A2(n_2483),
.B(n_2484),
.Y(n_2626)
);

A2O1A1Ixp33_ASAP7_75t_L g2627 ( 
.A1(n_2556),
.A2(n_2481),
.B(n_2494),
.C(n_2503),
.Y(n_2627)
);

AOI222xp33_ASAP7_75t_L g2628 ( 
.A1(n_2548),
.A2(n_2475),
.B1(n_2487),
.B2(n_2498),
.C1(n_2496),
.C2(n_2491),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_2593),
.B(n_2539),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2558),
.Y(n_2630)
);

OR2x2_ASAP7_75t_L g2631 ( 
.A(n_2577),
.B(n_2525),
.Y(n_2631)
);

AND2x4_ASAP7_75t_L g2632 ( 
.A(n_2559),
.B(n_2529),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2585),
.Y(n_2633)
);

O2A1O1Ixp33_ASAP7_75t_L g2634 ( 
.A1(n_2606),
.A2(n_2527),
.B(n_2530),
.C(n_2508),
.Y(n_2634)
);

OAI21xp33_ASAP7_75t_SL g2635 ( 
.A1(n_2561),
.A2(n_2486),
.B(n_2519),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2605),
.B(n_2603),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2583),
.Y(n_2637)
);

NOR2x1p5_ASAP7_75t_L g2638 ( 
.A(n_2586),
.B(n_2537),
.Y(n_2638)
);

OAI21xp33_ASAP7_75t_L g2639 ( 
.A1(n_2598),
.A2(n_2531),
.B(n_2529),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2558),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2588),
.B(n_2492),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2549),
.Y(n_2642)
);

OAI21xp5_ASAP7_75t_L g2643 ( 
.A1(n_2561),
.A2(n_2598),
.B(n_2503),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2583),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2601),
.Y(n_2645)
);

AOI221xp5_ASAP7_75t_L g2646 ( 
.A1(n_2564),
.A2(n_2512),
.B1(n_2509),
.B2(n_2500),
.C(n_2544),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2605),
.B(n_2504),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2601),
.Y(n_2648)
);

INVx1_ASAP7_75t_SL g2649 ( 
.A(n_2594),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2604),
.B(n_2551),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2597),
.B(n_2492),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2552),
.Y(n_2652)
);

OAI22xp33_ASAP7_75t_L g2653 ( 
.A1(n_2574),
.A2(n_2420),
.B1(n_2416),
.B2(n_2502),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2641),
.B(n_2602),
.Y(n_2654)
);

OAI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2611),
.A2(n_2617),
.B1(n_2627),
.B2(n_2649),
.Y(n_2655)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2656 ( 
.A1(n_2627),
.A2(n_2626),
.B(n_2643),
.C(n_2628),
.D(n_2629),
.Y(n_2656)
);

OAI21xp5_ASAP7_75t_L g2657 ( 
.A1(n_2634),
.A2(n_2566),
.B(n_2563),
.Y(n_2657)
);

OAI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2653),
.A2(n_2590),
.B1(n_2584),
.B2(n_2575),
.Y(n_2658)
);

AOI211xp5_ASAP7_75t_L g2659 ( 
.A1(n_2653),
.A2(n_2544),
.B(n_2599),
.C(n_2594),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2651),
.B(n_2599),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2619),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2620),
.B(n_2549),
.Y(n_2662)
);

OAI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2624),
.A2(n_2502),
.B1(n_2589),
.B2(n_2506),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2619),
.B(n_2559),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2618),
.B(n_2591),
.Y(n_2665)
);

OR2x2_ASAP7_75t_L g2666 ( 
.A(n_2623),
.B(n_2547),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2610),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2610),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2614),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2619),
.B(n_2591),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2626),
.A2(n_2570),
.B1(n_2573),
.B2(n_2571),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2629),
.B(n_2553),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2621),
.Y(n_2673)
);

O2A1O1Ixp33_ASAP7_75t_L g2674 ( 
.A1(n_2643),
.A2(n_2587),
.B(n_2592),
.C(n_2579),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2616),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2633),
.Y(n_2676)
);

NAND2x1_ASAP7_75t_L g2677 ( 
.A(n_2632),
.B(n_2502),
.Y(n_2677)
);

NOR2xp33_ASAP7_75t_L g2678 ( 
.A(n_2635),
.B(n_2562),
.Y(n_2678)
);

OAI32xp33_ASAP7_75t_L g2679 ( 
.A1(n_2615),
.A2(n_2590),
.A3(n_2584),
.B1(n_2554),
.B2(n_2567),
.Y(n_2679)
);

AOI21xp5_ASAP7_75t_L g2680 ( 
.A1(n_2634),
.A2(n_2578),
.B(n_2596),
.Y(n_2680)
);

AOI221xp5_ASAP7_75t_L g2681 ( 
.A1(n_2646),
.A2(n_2600),
.B1(n_2538),
.B2(n_2569),
.C(n_2565),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2625),
.B(n_2565),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2632),
.B(n_2562),
.Y(n_2683)
);

OR2x2_ASAP7_75t_L g2684 ( 
.A(n_2622),
.B(n_2582),
.Y(n_2684)
);

NAND3xp33_ASAP7_75t_L g2685 ( 
.A(n_2647),
.B(n_2595),
.C(n_2569),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2636),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2630),
.B(n_2466),
.Y(n_2687)
);

OAI221xp5_ASAP7_75t_L g2688 ( 
.A1(n_2646),
.A2(n_2429),
.B1(n_2543),
.B2(n_2545),
.C(n_2546),
.Y(n_2688)
);

OAI21xp5_ASAP7_75t_L g2689 ( 
.A1(n_2636),
.A2(n_2534),
.B(n_2535),
.Y(n_2689)
);

OAI22xp5_ASAP7_75t_L g2690 ( 
.A1(n_2652),
.A2(n_2506),
.B1(n_2519),
.B2(n_2531),
.Y(n_2690)
);

NOR2x1_ASAP7_75t_L g2691 ( 
.A(n_2670),
.B(n_2638),
.Y(n_2691)
);

XNOR2x2_ASAP7_75t_L g2692 ( 
.A(n_2655),
.B(n_2658),
.Y(n_2692)
);

AOI32xp33_ASAP7_75t_L g2693 ( 
.A1(n_2655),
.A2(n_2647),
.A3(n_2650),
.B1(n_2645),
.B2(n_2644),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2660),
.B(n_2640),
.Y(n_2694)
);

AOI221xp5_ASAP7_75t_L g2695 ( 
.A1(n_2657),
.A2(n_2650),
.B1(n_2648),
.B2(n_2637),
.C(n_2609),
.Y(n_2695)
);

AOI21xp33_ASAP7_75t_SL g2696 ( 
.A1(n_2658),
.A2(n_2631),
.B(n_2613),
.Y(n_2696)
);

NAND2x1_ASAP7_75t_SL g2697 ( 
.A(n_2654),
.B(n_2612),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2662),
.B(n_2661),
.Y(n_2698)
);

INVx1_ASAP7_75t_SL g2699 ( 
.A(n_2684),
.Y(n_2699)
);

BUFx2_ASAP7_75t_L g2700 ( 
.A(n_2689),
.Y(n_2700)
);

O2A1O1Ixp33_ASAP7_75t_L g2701 ( 
.A1(n_2656),
.A2(n_2608),
.B(n_2642),
.C(n_2639),
.Y(n_2701)
);

NAND2x1_ASAP7_75t_L g2702 ( 
.A(n_2683),
.B(n_2664),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2675),
.B(n_2466),
.Y(n_2703)
);

CKINVDCx6p67_ASAP7_75t_R g2704 ( 
.A(n_2672),
.Y(n_2704)
);

INVxp67_ASAP7_75t_L g2705 ( 
.A(n_2678),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2659),
.B(n_2474),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2686),
.B(n_2474),
.Y(n_2707)
);

OR2x2_ASAP7_75t_L g2708 ( 
.A(n_2665),
.B(n_2532),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2677),
.B(n_2517),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2666),
.Y(n_2710)
);

AOI21xp33_ASAP7_75t_SL g2711 ( 
.A1(n_2663),
.A2(n_2535),
.B(n_2546),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2680),
.B(n_2532),
.Y(n_2712)
);

OAI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_2671),
.A2(n_2543),
.B1(n_2459),
.B2(n_2536),
.Y(n_2713)
);

NOR2xp33_ASAP7_75t_SL g2714 ( 
.A(n_2657),
.B(n_2542),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2689),
.B(n_2536),
.Y(n_2715)
);

OAI221xp5_ASAP7_75t_SL g2716 ( 
.A1(n_2688),
.A2(n_2542),
.B1(n_2517),
.B2(n_2459),
.C(n_2463),
.Y(n_2716)
);

OAI22xp5_ASAP7_75t_L g2717 ( 
.A1(n_2685),
.A2(n_2452),
.B1(n_2444),
.B2(n_2461),
.Y(n_2717)
);

AOI321xp33_ASAP7_75t_SL g2718 ( 
.A1(n_2679),
.A2(n_2433),
.A3(n_2316),
.B1(n_2435),
.B2(n_2461),
.C(n_2465),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2681),
.B(n_2374),
.Y(n_2719)
);

OAI22xp33_ASAP7_75t_L g2720 ( 
.A1(n_2687),
.A2(n_2446),
.B1(n_2450),
.B2(n_2310),
.Y(n_2720)
);

AOI21xp33_ASAP7_75t_L g2721 ( 
.A1(n_2674),
.A2(n_2433),
.B(n_2353),
.Y(n_2721)
);

AOI322xp5_ASAP7_75t_L g2722 ( 
.A1(n_2713),
.A2(n_2668),
.A3(n_2667),
.B1(n_2669),
.B2(n_2673),
.C1(n_2676),
.C2(n_2682),
.Y(n_2722)
);

OAI31xp33_ASAP7_75t_L g2723 ( 
.A1(n_2716),
.A2(n_2690),
.A3(n_2316),
.B(n_2336),
.Y(n_2723)
);

NOR2x1_ASAP7_75t_L g2724 ( 
.A(n_2694),
.B(n_2690),
.Y(n_2724)
);

AOI322xp5_ASAP7_75t_L g2725 ( 
.A1(n_2719),
.A2(n_2712),
.A3(n_2695),
.B1(n_2706),
.B2(n_2699),
.C1(n_2700),
.C2(n_2705),
.Y(n_2725)
);

NAND3xp33_ASAP7_75t_L g2726 ( 
.A(n_2693),
.B(n_2353),
.C(n_2336),
.Y(n_2726)
);

OAI221xp5_ASAP7_75t_L g2727 ( 
.A1(n_2714),
.A2(n_2310),
.B1(n_2058),
.B2(n_2131),
.C(n_2333),
.Y(n_2727)
);

NOR2x1_ASAP7_75t_L g2728 ( 
.A(n_2702),
.B(n_2353),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2699),
.B(n_2697),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2704),
.Y(n_2730)
);

AOI221xp5_ASAP7_75t_L g2731 ( 
.A1(n_2696),
.A2(n_2336),
.B1(n_2333),
.B2(n_492),
.C(n_493),
.Y(n_2731)
);

OAI21xp5_ASAP7_75t_SL g2732 ( 
.A1(n_2709),
.A2(n_2333),
.B(n_23),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2703),
.Y(n_2733)
);

NAND4xp25_ASAP7_75t_SL g2734 ( 
.A(n_2701),
.B(n_27),
.C(n_24),
.D(n_25),
.Y(n_2734)
);

OAI221xp5_ASAP7_75t_L g2735 ( 
.A1(n_2721),
.A2(n_2070),
.B1(n_2098),
.B2(n_2082),
.C(n_2103),
.Y(n_2735)
);

NOR4xp25_ASAP7_75t_L g2736 ( 
.A(n_2710),
.B(n_32),
.C(n_28),
.D(n_31),
.Y(n_2736)
);

AOI21xp33_ASAP7_75t_L g2737 ( 
.A1(n_2715),
.A2(n_489),
.B(n_481),
.Y(n_2737)
);

OAI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2708),
.A2(n_2691),
.B1(n_2707),
.B2(n_2698),
.Y(n_2738)
);

OAI221xp5_ASAP7_75t_L g2739 ( 
.A1(n_2717),
.A2(n_2110),
.B1(n_1125),
.B2(n_1140),
.C(n_1101),
.Y(n_2739)
);

OAI211xp5_ASAP7_75t_L g2740 ( 
.A1(n_2711),
.A2(n_34),
.B(n_31),
.C(n_32),
.Y(n_2740)
);

NOR3xp33_ASAP7_75t_SL g2741 ( 
.A(n_2692),
.B(n_34),
.C(n_37),
.Y(n_2741)
);

OAI32xp33_ASAP7_75t_L g2742 ( 
.A1(n_2718),
.A2(n_39),
.A3(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_2717),
.B(n_41),
.Y(n_2743)
);

NAND3xp33_ASAP7_75t_SL g2744 ( 
.A(n_2720),
.B(n_502),
.C(n_500),
.Y(n_2744)
);

AND2x2_ASAP7_75t_L g2745 ( 
.A(n_2724),
.B(n_42),
.Y(n_2745)
);

AOI21xp5_ASAP7_75t_L g2746 ( 
.A1(n_2729),
.A2(n_42),
.B(n_44),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2734),
.A2(n_2728),
.B1(n_2726),
.B2(n_2727),
.Y(n_2747)
);

AOI22xp5_ASAP7_75t_L g2748 ( 
.A1(n_2738),
.A2(n_1847),
.B1(n_1960),
.B2(n_2072),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2733),
.Y(n_2749)
);

AOI211xp5_ASAP7_75t_L g2750 ( 
.A1(n_2742),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_2750)
);

O2A1O1Ixp33_ASAP7_75t_L g2751 ( 
.A1(n_2741),
.A2(n_50),
.B(n_45),
.C(n_47),
.Y(n_2751)
);

OAI221xp5_ASAP7_75t_L g2752 ( 
.A1(n_2732),
.A2(n_1125),
.B1(n_1140),
.B2(n_1101),
.C(n_1072),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2736),
.B(n_47),
.Y(n_2753)
);

AOI21xp5_ASAP7_75t_L g2754 ( 
.A1(n_2740),
.A2(n_51),
.B(n_52),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2730),
.Y(n_2755)
);

NOR3xp33_ASAP7_75t_L g2756 ( 
.A(n_2743),
.B(n_1125),
.C(n_1072),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2739),
.Y(n_2757)
);

AOI21xp33_ASAP7_75t_L g2758 ( 
.A1(n_2723),
.A2(n_509),
.B(n_505),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2737),
.B(n_2744),
.Y(n_2759)
);

OAI22xp5_ASAP7_75t_L g2760 ( 
.A1(n_2731),
.A2(n_1874),
.B1(n_1878),
.B2(n_529),
.Y(n_2760)
);

AOI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_2745),
.A2(n_2750),
.B1(n_2759),
.B2(n_2756),
.Y(n_2761)
);

AOI22xp5_ASAP7_75t_L g2762 ( 
.A1(n_2753),
.A2(n_2735),
.B1(n_2725),
.B2(n_2722),
.Y(n_2762)
);

AOI322xp5_ASAP7_75t_L g2763 ( 
.A1(n_2747),
.A2(n_2749),
.A3(n_2757),
.B1(n_2755),
.B2(n_2758),
.C1(n_2751),
.C2(n_2748),
.Y(n_2763)
);

AOI31xp33_ASAP7_75t_L g2764 ( 
.A1(n_2746),
.A2(n_56),
.A3(n_54),
.B(n_55),
.Y(n_2764)
);

OAI21xp33_ASAP7_75t_L g2765 ( 
.A1(n_2754),
.A2(n_1910),
.B(n_530),
.Y(n_2765)
);

AOI221xp5_ASAP7_75t_L g2766 ( 
.A1(n_2760),
.A2(n_551),
.B1(n_554),
.B2(n_545),
.C(n_516),
.Y(n_2766)
);

NOR2x1_ASAP7_75t_L g2767 ( 
.A(n_2752),
.B(n_55),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2745),
.B(n_57),
.Y(n_2768)
);

OAI311xp33_ASAP7_75t_L g2769 ( 
.A1(n_2762),
.A2(n_2761),
.A3(n_2763),
.B1(n_2765),
.C1(n_2768),
.Y(n_2769)
);

NAND3x1_ASAP7_75t_SL g2770 ( 
.A(n_2767),
.B(n_58),
.C(n_61),
.Y(n_2770)
);

AOI21xp5_ASAP7_75t_SL g2771 ( 
.A1(n_2764),
.A2(n_2766),
.B(n_61),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2762),
.B(n_64),
.Y(n_2772)
);

AOI211xp5_ASAP7_75t_SL g2773 ( 
.A1(n_2762),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_2773)
);

INVxp33_ASAP7_75t_SL g2774 ( 
.A(n_2762),
.Y(n_2774)
);

OAI211xp5_ASAP7_75t_L g2775 ( 
.A1(n_2762),
.A2(n_69),
.B(n_65),
.C(n_67),
.Y(n_2775)
);

NOR4xp25_ASAP7_75t_L g2776 ( 
.A(n_2769),
.B(n_77),
.C(n_74),
.D(n_76),
.Y(n_2776)
);

OR2x6_ASAP7_75t_L g2777 ( 
.A(n_2771),
.B(n_846),
.Y(n_2777)
);

NAND4xp25_ASAP7_75t_L g2778 ( 
.A(n_2773),
.B(n_80),
.C(n_76),
.D(n_78),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2772),
.B(n_78),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2770),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2775),
.Y(n_2781)
);

INVxp67_ASAP7_75t_SL g2782 ( 
.A(n_2774),
.Y(n_2782)
);

NOR2xp67_ASAP7_75t_L g2783 ( 
.A(n_2775),
.B(n_83),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2770),
.Y(n_2784)
);

NOR3xp33_ASAP7_75t_L g2785 ( 
.A(n_2775),
.B(n_570),
.C(n_560),
.Y(n_2785)
);

HB1xp67_ASAP7_75t_L g2786 ( 
.A(n_2782),
.Y(n_2786)
);

XOR2xp5_ASAP7_75t_L g2787 ( 
.A(n_2778),
.B(n_84),
.Y(n_2787)
);

NOR2x1_ASAP7_75t_L g2788 ( 
.A(n_2780),
.B(n_84),
.Y(n_2788)
);

NOR2xp67_ASAP7_75t_L g2789 ( 
.A(n_2784),
.B(n_85),
.Y(n_2789)
);

NOR3x2_ASAP7_75t_L g2790 ( 
.A(n_2776),
.B(n_2785),
.C(n_2783),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_2781),
.B(n_86),
.Y(n_2791)
);

INVx2_ASAP7_75t_SL g2792 ( 
.A(n_2779),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2777),
.Y(n_2793)
);

AND2x4_ASAP7_75t_L g2794 ( 
.A(n_2780),
.B(n_92),
.Y(n_2794)
);

AOI221xp5_ASAP7_75t_L g2795 ( 
.A1(n_2786),
.A2(n_575),
.B1(n_581),
.B2(n_583),
.C(n_591),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2788),
.Y(n_2796)
);

NAND4xp25_ASAP7_75t_L g2797 ( 
.A(n_2791),
.B(n_98),
.C(n_95),
.D(n_96),
.Y(n_2797)
);

AOI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2792),
.A2(n_617),
.B1(n_625),
.B2(n_615),
.Y(n_2798)
);

OAI22xp5_ASAP7_75t_SL g2799 ( 
.A1(n_2787),
.A2(n_102),
.B1(n_99),
.B2(n_100),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2789),
.Y(n_2800)
);

OAI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2794),
.A2(n_1874),
.B1(n_1878),
.B2(n_1322),
.Y(n_2801)
);

INVx2_ASAP7_75t_SL g2802 ( 
.A(n_2796),
.Y(n_2802)
);

NAND4xp75_ASAP7_75t_L g2803 ( 
.A(n_2800),
.B(n_2793),
.C(n_2790),
.D(n_2794),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2799),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2798),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2797),
.B(n_105),
.Y(n_2806)
);

AOI22x1_ASAP7_75t_L g2807 ( 
.A1(n_2795),
.A2(n_2801),
.B1(n_110),
.B2(n_107),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2796),
.B(n_108),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2799),
.Y(n_2809)
);

OAI22x1_ASAP7_75t_L g2810 ( 
.A1(n_2807),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2806),
.Y(n_2811)
);

AND2x2_ASAP7_75t_SL g2812 ( 
.A(n_2804),
.B(n_2809),
.Y(n_2812)
);

BUFx3_ASAP7_75t_L g2813 ( 
.A(n_2805),
.Y(n_2813)
);

NAND3x1_ASAP7_75t_L g2814 ( 
.A(n_2808),
.B(n_116),
.C(n_117),
.Y(n_2814)
);

AOI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2802),
.A2(n_118),
.B(n_119),
.Y(n_2815)
);

XNOR2xp5_ASAP7_75t_L g2816 ( 
.A(n_2803),
.B(n_118),
.Y(n_2816)
);

OAI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2814),
.A2(n_797),
.B(n_779),
.Y(n_2817)
);

AOI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2812),
.A2(n_1074),
.B1(n_797),
.B2(n_827),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2810),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2816),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2813),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2821),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2819),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2820),
.Y(n_2824)
);

OAI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2817),
.A2(n_2811),
.B(n_2815),
.Y(n_2825)
);

BUFx2_ASAP7_75t_L g2826 ( 
.A(n_2818),
.Y(n_2826)
);

INVxp67_ASAP7_75t_SL g2827 ( 
.A(n_2821),
.Y(n_2827)
);

INVx1_ASAP7_75t_SL g2828 ( 
.A(n_2821),
.Y(n_2828)
);

AOI21x1_ASAP7_75t_L g2829 ( 
.A1(n_2821),
.A2(n_129),
.B(n_130),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2827),
.Y(n_2830)
);

OAI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2828),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2823),
.B(n_139),
.Y(n_2832)
);

CKINVDCx20_ASAP7_75t_R g2833 ( 
.A(n_2824),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2829),
.Y(n_2834)
);

AOI22x1_ASAP7_75t_L g2835 ( 
.A1(n_2826),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_2835)
);

OAI22xp5_ASAP7_75t_L g2836 ( 
.A1(n_2825),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_2836)
);

INVx4_ASAP7_75t_L g2837 ( 
.A(n_2822),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2827),
.A2(n_159),
.B(n_160),
.Y(n_2838)
);

OAI211xp5_ASAP7_75t_L g2839 ( 
.A1(n_2827),
.A2(n_163),
.B(n_164),
.C(n_165),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2827),
.Y(n_2840)
);

OAI211xp5_ASAP7_75t_L g2841 ( 
.A1(n_2827),
.A2(n_167),
.B(n_168),
.C(n_169),
.Y(n_2841)
);

OA22x2_ASAP7_75t_L g2842 ( 
.A1(n_2840),
.A2(n_2837),
.B1(n_2841),
.B2(n_2839),
.Y(n_2842)
);

OAI22xp33_ASAP7_75t_L g2843 ( 
.A1(n_2836),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_2843)
);

AOI21xp5_ASAP7_75t_L g2844 ( 
.A1(n_2832),
.A2(n_827),
.B(n_178),
.Y(n_2844)
);

OAI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2835),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_2845)
);

OAI21x1_ASAP7_75t_L g2846 ( 
.A1(n_2838),
.A2(n_185),
.B(n_186),
.Y(n_2846)
);

AOI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2831),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.Y(n_2847)
);

OA21x2_ASAP7_75t_L g2848 ( 
.A1(n_2830),
.A2(n_202),
.B(n_203),
.Y(n_2848)
);

AO22x2_ASAP7_75t_L g2849 ( 
.A1(n_2834),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2837),
.B(n_205),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2833),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2833),
.Y(n_2852)
);

OAI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2851),
.A2(n_843),
.B(n_1240),
.Y(n_2853)
);

OAI21x1_ASAP7_75t_L g2854 ( 
.A1(n_2842),
.A2(n_209),
.B(n_210),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2852),
.Y(n_2855)
);

OAI21xp5_ASAP7_75t_L g2856 ( 
.A1(n_2846),
.A2(n_213),
.B(n_216),
.Y(n_2856)
);

AOI21xp5_ASAP7_75t_L g2857 ( 
.A1(n_2850),
.A2(n_808),
.B(n_791),
.Y(n_2857)
);

OAI22xp33_ASAP7_75t_L g2858 ( 
.A1(n_2847),
.A2(n_1129),
.B1(n_1090),
.B2(n_1091),
.Y(n_2858)
);

OAI22xp33_ASAP7_75t_L g2859 ( 
.A1(n_2845),
.A2(n_1139),
.B1(n_1090),
.B2(n_1129),
.Y(n_2859)
);

AOI21xp33_ASAP7_75t_L g2860 ( 
.A1(n_2848),
.A2(n_220),
.B(n_221),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2849),
.Y(n_2861)
);

AOI22x1_ASAP7_75t_L g2862 ( 
.A1(n_2855),
.A2(n_2849),
.B1(n_2844),
.B2(n_2843),
.Y(n_2862)
);

AOI222xp33_ASAP7_75t_SL g2863 ( 
.A1(n_2861),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.C1(n_242),
.C2(n_246),
.Y(n_2863)
);

OAI222xp33_ASAP7_75t_L g2864 ( 
.A1(n_2859),
.A2(n_247),
.B1(n_248),
.B2(n_251),
.C1(n_253),
.C2(n_255),
.Y(n_2864)
);

AOI22xp5_ASAP7_75t_L g2865 ( 
.A1(n_2858),
.A2(n_2856),
.B1(n_2860),
.B2(n_2853),
.Y(n_2865)
);

AOI222xp33_ASAP7_75t_L g2866 ( 
.A1(n_2854),
.A2(n_2857),
.B1(n_808),
.B2(n_791),
.C1(n_774),
.C2(n_781),
.Y(n_2866)
);

OAI21xp5_ASAP7_75t_L g2867 ( 
.A1(n_2855),
.A2(n_259),
.B(n_263),
.Y(n_2867)
);

AOI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2865),
.A2(n_774),
.B1(n_791),
.B2(n_808),
.Y(n_2868)
);

AOI222xp33_ASAP7_75t_L g2869 ( 
.A1(n_2864),
.A2(n_808),
.B1(n_791),
.B2(n_774),
.C1(n_781),
.C2(n_270),
.Y(n_2869)
);

AOI22xp5_ASAP7_75t_SL g2870 ( 
.A1(n_2867),
.A2(n_264),
.B1(n_266),
.B2(n_268),
.Y(n_2870)
);

AOI22xp5_ASAP7_75t_L g2871 ( 
.A1(n_2863),
.A2(n_774),
.B1(n_791),
.B2(n_808),
.Y(n_2871)
);

AOI222xp33_ASAP7_75t_L g2872 ( 
.A1(n_2862),
.A2(n_774),
.B1(n_781),
.B2(n_272),
.C1(n_275),
.C2(n_276),
.Y(n_2872)
);

AOI22xp5_ASAP7_75t_L g2873 ( 
.A1(n_2866),
.A2(n_781),
.B1(n_1225),
.B2(n_1234),
.Y(n_2873)
);

OAI21xp5_ASAP7_75t_L g2874 ( 
.A1(n_2870),
.A2(n_2869),
.B(n_2872),
.Y(n_2874)
);

AO21x2_ASAP7_75t_L g2875 ( 
.A1(n_2868),
.A2(n_285),
.B(n_289),
.Y(n_2875)
);

AOI21xp5_ASAP7_75t_L g2876 ( 
.A1(n_2874),
.A2(n_2873),
.B(n_2871),
.Y(n_2876)
);

AOI211xp5_ASAP7_75t_L g2877 ( 
.A1(n_2876),
.A2(n_2875),
.B(n_303),
.C(n_304),
.Y(n_2877)
);


endmodule