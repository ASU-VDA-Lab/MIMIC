module fake_netlist_6_3608_n_1835 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1835);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1835;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_155),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_82),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_109),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_20),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_16),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_15),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_4),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_27),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_21),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_56),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_189),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_58),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_156),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_157),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_50),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_38),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_25),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_104),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_9),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_111),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_70),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_0),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_4),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_69),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_127),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_161),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_179),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_89),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_67),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_20),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_113),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_16),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_81),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_78),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_169),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_99),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_90),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_56),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_50),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_57),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_154),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_43),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_160),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_48),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_94),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_141),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_153),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_107),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_6),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_138),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_100),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_164),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_49),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_181),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_148),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_27),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_114),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_9),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_133),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_130),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_85),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_19),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_10),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_15),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_39),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_57),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_172),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_47),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_33),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_143),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_188),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_174),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_13),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_43),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_183),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_121),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_58),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_77),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_61),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_134),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_42),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_19),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_103),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_31),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_117),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_110),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_72),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_86),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_73),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_135),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_71),
.Y(n_293)
);

INVxp33_ASAP7_75t_SL g294 ( 
.A(n_34),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_12),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_125),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_23),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_25),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_62),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_3),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_29),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_18),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_80),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_53),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_41),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_144),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_39),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_55),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_35),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_118),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_129),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_122),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_21),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_178),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_131),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_126),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_29),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_46),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_45),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_1),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_140),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_3),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_75),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_177),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_96),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_102),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_23),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_88),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_152),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_14),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_139),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_112),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_48),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_51),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_33),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_68),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_32),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_12),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_63),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_147),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_44),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_173),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_146),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_92),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_65),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_10),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_182),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_175),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_0),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_93),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_91),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_185),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_76),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_165),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_123),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_7),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_159),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_116),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_128),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_51),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_35),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_13),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_132),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_171),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_2),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_24),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_54),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_24),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_28),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_59),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_167),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_59),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_108),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_150),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_97),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_22),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_6),
.Y(n_377)
);

INVx4_ASAP7_75t_R g378 ( 
.A(n_26),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_87),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_346),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_272),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_196),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_233),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_270),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_196),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_196),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_196),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_235),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_196),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_369),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_240),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_308),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_308),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_308),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_291),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_296),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_308),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_234),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_308),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_207),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_234),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_263),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_207),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_228),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_228),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_263),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_239),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_299),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_365),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_365),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_361),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_209),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_366),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_366),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_237),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_247),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_330),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_249),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_193),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_199),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_263),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_236),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_328),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_253),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_260),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_194),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_311),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_253),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_271),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_283),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_250),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_284),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_286),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_297),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_305),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_327),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_333),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_353),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_361),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_334),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_335),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_263),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_341),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_195),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_202),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_360),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_343),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_218),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_368),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_204),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_204),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_220),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_211),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_351),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_224),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_231),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_211),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_254),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_243),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_213),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_361),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_213),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_241),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_241),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_256),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_257),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_262),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_195),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_273),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_263),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_277),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_382),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_381),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_446),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_393),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_413),
.A2(n_238),
.B1(n_309),
.B2(n_294),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_383),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_395),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_447),
.B(n_244),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_244),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_428),
.A2(n_201),
.B1(n_377),
.B2(n_376),
.Y(n_486)
);

AND2x2_ASAP7_75t_SL g487 ( 
.A(n_440),
.B(n_256),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_382),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_385),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_454),
.B(n_269),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_398),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_452),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_403),
.B(n_261),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_461),
.B(n_269),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_407),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_423),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_388),
.B(n_252),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_386),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_401),
.B(n_285),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_423),
.B(n_245),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_408),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_386),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_425),
.B(n_398),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_285),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_387),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_387),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_458),
.B(n_190),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_402),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_389),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_415),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_419),
.B(n_336),
.Y(n_515)
);

AND2x2_ASAP7_75t_SL g516 ( 
.A(n_384),
.B(n_336),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_418),
.B(n_274),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_420),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_441),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_389),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_463),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_392),
.B(n_190),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_392),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_394),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_394),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_390),
.B(n_275),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_470),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_397),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_419),
.B(n_375),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_397),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_452),
.B(n_453),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_399),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_444),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_399),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_444),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_453),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_396),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_409),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_455),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_472),
.Y(n_541)
);

OA21x2_ASAP7_75t_L g542 ( 
.A1(n_459),
.A2(n_375),
.B(n_259),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_472),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_384),
.Y(n_544)
);

OA21x2_ASAP7_75t_L g545 ( 
.A1(n_459),
.A2(n_290),
.B(n_248),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_462),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_462),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_464),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_464),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_465),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_412),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_465),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_481),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_477),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_533),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_481),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_506),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_477),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_477),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_533),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_551),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_480),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_502),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_551),
.Y(n_565)
);

BUFx4f_ASAP7_75t_L g566 ( 
.A(n_545),
.Y(n_566)
);

OAI22xp33_ASAP7_75t_L g567 ( 
.A1(n_526),
.A2(n_391),
.B1(n_322),
.B2(n_276),
.Y(n_567)
);

AND2x6_ASAP7_75t_L g568 ( 
.A(n_501),
.B(n_261),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_533),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_502),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_480),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_499),
.B(n_433),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_517),
.B(n_469),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_516),
.B(n_471),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_535),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_516),
.B(n_473),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_506),
.B(n_466),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_501),
.B(n_466),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_535),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_492),
.B(n_467),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_492),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_535),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_489),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_514),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_487),
.B(n_460),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_543),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_501),
.B(n_467),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_487),
.B(n_468),
.Y(n_588)
);

INVx8_ASAP7_75t_L g589 ( 
.A(n_494),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_475),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_489),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_481),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_519),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_489),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_516),
.A2(n_367),
.B1(n_417),
.B2(n_246),
.Y(n_595)
);

AO21x2_ASAP7_75t_L g596 ( 
.A1(n_503),
.A2(n_314),
.B(n_292),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_493),
.B(n_426),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_543),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_514),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_505),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_487),
.B(n_426),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_543),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_514),
.B(n_430),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_507),
.B(n_261),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_505),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_474),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_505),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_492),
.B(n_430),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_474),
.Y(n_609)
);

NOR2x1p5_ASAP7_75t_L g610 ( 
.A(n_479),
.B(n_197),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_483),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_508),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_509),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_481),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_509),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_509),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_481),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_504),
.B(n_253),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_488),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_488),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_490),
.Y(n_621)
);

CKINVDCx11_ASAP7_75t_R g622 ( 
.A(n_537),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_490),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_508),
.B(n_456),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_478),
.B(n_429),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_500),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_500),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_510),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_510),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_508),
.B(n_449),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_513),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_518),
.B(n_191),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_515),
.B(n_400),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_512),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_513),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_520),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_526),
.B(n_191),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_520),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_493),
.B(n_289),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_481),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_515),
.B(n_400),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_484),
.B(n_323),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_481),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_523),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_523),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_524),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_515),
.B(n_404),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_524),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_495),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_485),
.B(n_278),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_495),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_525),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_525),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_527),
.B(n_192),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_528),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_529),
.B(n_507),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_528),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_530),
.Y(n_658)
);

AO21x2_ASAP7_75t_L g659 ( 
.A1(n_503),
.A2(n_321),
.B(n_316),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_530),
.Y(n_660)
);

AO22x2_ASAP7_75t_L g661 ( 
.A1(n_478),
.A2(n_345),
.B1(n_325),
.B2(n_331),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_532),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_532),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_534),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_491),
.A2(n_427),
.B1(n_326),
.B2(n_261),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_SL g666 ( 
.A(n_519),
.B(n_197),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_476),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_534),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_512),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_497),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_527),
.B(n_192),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_512),
.B(n_200),
.Y(n_672)
);

CKINVDCx16_ASAP7_75t_R g673 ( 
.A(n_539),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_491),
.B(n_280),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_495),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_495),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_497),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_486),
.A2(n_217),
.B1(n_216),
.B2(n_377),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_496),
.B(n_282),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_482),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_497),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_496),
.B(n_287),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_495),
.Y(n_683)
);

OR2x6_ASAP7_75t_L g684 ( 
.A(n_529),
.B(n_344),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_495),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_522),
.B(n_288),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_544),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_529),
.B(n_404),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_497),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_548),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_476),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_511),
.A2(n_319),
.B1(n_317),
.B2(n_307),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_511),
.B(n_200),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_531),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_522),
.B(n_293),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_495),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_498),
.B(n_303),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_SL g698 ( 
.A(n_521),
.B(n_198),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_548),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_531),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_482),
.B(n_348),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_531),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_694),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_584),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_677),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_656),
.B(n_498),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_624),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_589),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_656),
.B(n_498),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_584),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_599),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_693),
.B(n_498),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_568),
.B(n_263),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_558),
.B(n_554),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_SL g715 ( 
.A(n_562),
.B(n_203),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_589),
.Y(n_716)
);

NOR2xp67_ASAP7_75t_L g717 ( 
.A(n_572),
.B(n_507),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_678),
.A2(n_198),
.B1(n_376),
.B2(n_372),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_599),
.B(n_203),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_558),
.B(n_498),
.Y(n_720)
);

A2O1A1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_700),
.A2(n_424),
.B(n_421),
.C(n_422),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_554),
.B(n_498),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_L g723 ( 
.A(n_568),
.B(n_263),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_556),
.B(n_498),
.Y(n_724)
);

NAND2x1_ASAP7_75t_L g725 ( 
.A(n_553),
.B(n_494),
.Y(n_725)
);

BUFx6f_ASAP7_75t_SL g726 ( 
.A(n_667),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_556),
.B(n_541),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_702),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_667),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_702),
.Y(n_730)
);

BUFx6f_ASAP7_75t_SL g731 ( 
.A(n_667),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_601),
.A2(n_379),
.B1(n_306),
.B2(n_310),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_633),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_566),
.B(n_261),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_SL g735 ( 
.A(n_610),
.B(n_573),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_589),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_642),
.B(n_205),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_561),
.B(n_569),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_574),
.B(n_205),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_561),
.B(n_541),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_576),
.B(n_206),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_689),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_633),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_581),
.B(n_542),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_L g745 ( 
.A(n_568),
.B(n_263),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_667),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_569),
.B(n_686),
.Y(n_747)
);

NOR2x1p5_ASAP7_75t_SL g748 ( 
.A(n_583),
.B(n_548),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_581),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_695),
.B(n_541),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_641),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_555),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_650),
.B(n_541),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_612),
.B(n_422),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_669),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_597),
.B(n_206),
.Y(n_756)
);

BUFx5_ASAP7_75t_L g757 ( 
.A(n_575),
.Y(n_757)
);

INVx8_ASAP7_75t_L g758 ( 
.A(n_701),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_589),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_674),
.B(n_679),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_621),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_682),
.B(n_541),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_639),
.B(n_210),
.Y(n_763)
);

AOI22x1_ASAP7_75t_L g764 ( 
.A1(n_606),
.A2(n_355),
.B1(n_550),
.B2(n_547),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_641),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_555),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_566),
.B(n_326),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_566),
.A2(n_661),
.B1(n_568),
.B2(n_647),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_691),
.B(n_424),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_559),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_578),
.B(n_541),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_559),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_587),
.B(n_577),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_612),
.B(n_326),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_669),
.B(n_210),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_560),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_585),
.A2(n_312),
.B1(n_315),
.B2(n_342),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_647),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_634),
.B(n_326),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_570),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_634),
.B(n_541),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_606),
.B(n_545),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_661),
.A2(n_545),
.B1(n_542),
.B2(n_326),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_692),
.A2(n_595),
.B(n_619),
.C(n_609),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_580),
.B(n_347),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_570),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_588),
.A2(n_350),
.B1(n_352),
.B2(n_354),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_621),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_580),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_609),
.B(n_545),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_SL g791 ( 
.A1(n_637),
.A2(n_338),
.B1(n_226),
.B2(n_223),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_619),
.B(n_545),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_688),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_688),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_620),
.A2(n_626),
.B(n_629),
.C(n_627),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_563),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_620),
.B(n_546),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_564),
.B(n_431),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_626),
.B(n_546),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_580),
.B(n_623),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_593),
.B(n_431),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_563),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_623),
.B(n_357),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_654),
.B(n_214),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_671),
.B(n_603),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_628),
.B(n_358),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_666),
.B(n_432),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_SL g808 ( 
.A(n_562),
.B(n_214),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_628),
.B(n_636),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_571),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_627),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_608),
.B(n_432),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_636),
.B(n_359),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_629),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_672),
.B(n_251),
.C(n_242),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_644),
.B(n_363),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_631),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_631),
.B(n_546),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_687),
.B(n_215),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_651),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_651),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_632),
.B(n_215),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_635),
.B(n_546),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_635),
.B(n_546),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_610),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_638),
.B(n_546),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_638),
.B(n_645),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_645),
.B(n_546),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_652),
.B(n_549),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_657),
.B(n_549),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_657),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_644),
.B(n_646),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_651),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_660),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_651),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_662),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_630),
.B(n_680),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_662),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_646),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_648),
.B(n_364),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_661),
.A2(n_542),
.B1(n_494),
.B2(n_547),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_648),
.B(n_549),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_653),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_653),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_567),
.B(n_618),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_655),
.B(n_549),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_655),
.Y(n_847)
);

NOR2x1p5_ASAP7_75t_L g848 ( 
.A(n_565),
.B(n_201),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_658),
.B(n_549),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_568),
.B(n_219),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_684),
.B(n_698),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_684),
.A2(n_339),
.B1(n_221),
.B2(n_222),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_661),
.A2(n_542),
.B1(n_494),
.B2(n_552),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_697),
.A2(n_542),
.B(n_550),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_658),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_680),
.B(n_434),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_663),
.B(n_536),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_663),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_664),
.B(n_536),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_684),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_717),
.B(n_565),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_786),
.B(n_780),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_761),
.Y(n_863)
);

NAND2xp33_ASAP7_75t_L g864 ( 
.A(n_708),
.B(n_568),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_773),
.B(n_664),
.Y(n_865)
);

NAND2x1p5_ASAP7_75t_L g866 ( 
.A(n_708),
.B(n_736),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_786),
.Y(n_867)
);

NOR2x2_ASAP7_75t_L g868 ( 
.A(n_718),
.B(n_701),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_758),
.B(n_701),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_760),
.B(n_668),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_704),
.B(n_625),
.Y(n_871)
);

NOR2xp67_ASAP7_75t_L g872 ( 
.A(n_815),
.B(n_590),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_788),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_707),
.Y(n_874)
);

AO22x1_ASAP7_75t_L g875 ( 
.A1(n_845),
.A2(n_819),
.B1(n_741),
.B2(n_739),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_710),
.B(n_625),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_768),
.A2(n_678),
.B1(n_665),
.B2(n_684),
.Y(n_877)
);

AND2x6_ASAP7_75t_L g878 ( 
.A(n_708),
.B(n_592),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_836),
.B(n_668),
.Y(n_879)
);

NOR2x1_ASAP7_75t_R g880 ( 
.A(n_749),
.B(n_622),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_845),
.A2(n_684),
.B1(n_568),
.B2(n_604),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_844),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_775),
.B(n_590),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_711),
.B(n_763),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_836),
.B(n_670),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_844),
.Y(n_886)
);

INVx5_ASAP7_75t_L g887 ( 
.A(n_708),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_819),
.A2(n_604),
.B1(n_659),
.B2(n_596),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_858),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_737),
.B(n_670),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_749),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_763),
.B(n_611),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_703),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_755),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_747),
.B(n_681),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_805),
.B(n_611),
.Y(n_896)
);

NAND2x1_ASAP7_75t_L g897 ( 
.A(n_736),
.B(n_592),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_798),
.B(n_673),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_739),
.A2(n_604),
.B1(n_659),
.B2(n_596),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_706),
.B(n_681),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_769),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_839),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_709),
.B(n_575),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_741),
.A2(n_604),
.B1(n_659),
.B2(n_596),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_755),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_805),
.B(n_673),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_775),
.B(n_701),
.Y(n_907)
);

OR2x6_ASAP7_75t_L g908 ( 
.A(n_758),
.B(n_701),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_789),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_R g910 ( 
.A(n_735),
.B(n_219),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_715),
.B(n_553),
.Y(n_911)
);

INVx5_ASAP7_75t_L g912 ( 
.A(n_736),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_856),
.B(n_434),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_707),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_728),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_730),
.Y(n_916)
);

BUFx4f_ASAP7_75t_SL g917 ( 
.A(n_825),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_733),
.A2(n_604),
.B1(n_699),
.B2(n_690),
.Y(n_918)
);

AOI22x1_ASAP7_75t_SL g919 ( 
.A1(n_743),
.A2(n_370),
.B1(n_226),
.B2(n_223),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_714),
.B(n_579),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_789),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_827),
.B(n_579),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_811),
.B(n_582),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_851),
.B(n_225),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_814),
.B(n_582),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_751),
.B(n_435),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_817),
.B(n_586),
.Y(n_927)
);

BUFx4f_ASAP7_75t_L g928 ( 
.A(n_758),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_851),
.B(n_225),
.Y(n_929)
);

NAND2x2_ASAP7_75t_L g930 ( 
.A(n_848),
.B(n_378),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_SL g931 ( 
.A1(n_804),
.A2(n_370),
.B1(n_217),
.B2(n_216),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_843),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_831),
.B(n_586),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_765),
.B(n_435),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_847),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_778),
.A2(n_604),
.B1(n_699),
.B2(n_690),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_855),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_756),
.B(n_227),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_752),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_793),
.B(n_436),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_860),
.B(n_436),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_834),
.B(n_598),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_820),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_838),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_794),
.A2(n_604),
.B1(n_602),
.B2(n_598),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_801),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_800),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_800),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_809),
.Y(n_949)
);

NAND3xp33_ASAP7_75t_SL g950 ( 
.A(n_804),
.B(n_212),
.C(n_208),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_837),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_807),
.Y(n_952)
);

NOR2x2_ASAP7_75t_L g953 ( 
.A(n_718),
.B(n_208),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_716),
.A2(n_649),
.B(n_557),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_756),
.B(n_227),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_754),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_860),
.B(n_437),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_719),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_719),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_729),
.B(n_437),
.Y(n_960)
);

NAND2x2_ASAP7_75t_L g961 ( 
.A(n_746),
.B(n_212),
.Y(n_961)
);

INVx5_ASAP7_75t_L g962 ( 
.A(n_736),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_809),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_832),
.Y(n_964)
);

OR2x6_ASAP7_75t_L g965 ( 
.A(n_784),
.B(n_438),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_820),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_754),
.B(n_229),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_768),
.A2(n_602),
.B1(n_591),
.B2(n_594),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_812),
.B(n_229),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_841),
.A2(n_853),
.B1(n_783),
.B2(n_852),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_785),
.B(n_438),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_738),
.B(n_592),
.Y(n_972)
);

INVx5_ASAP7_75t_L g973 ( 
.A(n_716),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_822),
.B(n_230),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_785),
.B(n_439),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_822),
.B(n_439),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_720),
.B(n_442),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_820),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_SL g979 ( 
.A1(n_808),
.A2(n_320),
.B1(n_337),
.B2(n_338),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_766),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_771),
.B(n_614),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_803),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_732),
.B(n_230),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_777),
.B(n_232),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_803),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_787),
.B(n_232),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_726),
.Y(n_987)
);

INVx4_ASAP7_75t_L g988 ( 
.A(n_821),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_832),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_SL g990 ( 
.A1(n_841),
.A2(n_320),
.B1(n_337),
.B2(n_372),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_712),
.B(n_617),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_857),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_853),
.A2(n_281),
.B1(n_258),
.B2(n_267),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_770),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_782),
.B(n_617),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_795),
.A2(n_696),
.B(n_685),
.C(n_683),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_790),
.B(n_617),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_806),
.B(n_442),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_806),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_726),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_859),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_791),
.B(n_557),
.Y(n_1002)
);

AND2x6_ASAP7_75t_SL g1003 ( 
.A(n_731),
.B(n_443),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_734),
.A2(n_767),
.B1(n_764),
.B2(n_744),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_772),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_759),
.B(n_324),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_821),
.B(n_329),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_813),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_705),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_813),
.B(n_649),
.Y(n_1010)
);

INVx5_ASAP7_75t_L g1011 ( 
.A(n_821),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_742),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_816),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_821),
.B(n_329),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_835),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_835),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_792),
.B(n_640),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_835),
.B(n_332),
.Y(n_1018)
);

BUFx4f_ASAP7_75t_L g1019 ( 
.A(n_744),
.Y(n_1019)
);

BUFx4f_ASAP7_75t_L g1020 ( 
.A(n_835),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_776),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_757),
.B(n_734),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_796),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_833),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_802),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_757),
.B(n_640),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_725),
.Y(n_1027)
);

BUFx8_ASAP7_75t_L g1028 ( 
.A(n_731),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_810),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_816),
.B(n_443),
.Y(n_1030)
);

OAI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_750),
.A2(n_753),
.B1(n_762),
.B2(n_824),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_833),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_757),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_944),
.Y(n_1034)
);

AND3x4_ASAP7_75t_L g1035 ( 
.A(n_951),
.B(n_721),
.C(n_268),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_907),
.A2(n_748),
.B(n_767),
.C(n_854),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_875),
.B(n_976),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_867),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_956),
.B(n_840),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_870),
.A2(n_783),
.B1(n_781),
.B2(n_724),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_958),
.A2(n_840),
.B(n_797),
.C(n_799),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_870),
.B(n_757),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_959),
.A2(n_823),
.B(n_818),
.C(n_826),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_893),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_954),
.A2(n_722),
.B(n_727),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_973),
.A2(n_740),
.B(n_651),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_973),
.A2(n_850),
.B(n_829),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_938),
.B(n_830),
.C(n_828),
.Y(n_1048)
);

INVx5_ASAP7_75t_L g1049 ( 
.A(n_943),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_1024),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_865),
.B(n_774),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_973),
.A2(n_713),
.B(n_723),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1004),
.A2(n_779),
.B1(n_774),
.B2(n_842),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_995),
.A2(n_849),
.B(n_846),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_862),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_974),
.A2(n_779),
.B(n_745),
.C(n_448),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_901),
.B(n_332),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_992),
.B(n_1001),
.Y(n_1058)
);

BUFx4_ASAP7_75t_SL g1059 ( 
.A(n_1003),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_891),
.B(n_445),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_952),
.A2(n_685),
.B1(n_683),
.B2(n_676),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_SL g1062 ( 
.A(n_950),
.B(n_304),
.C(n_302),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_946),
.B(n_339),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_952),
.B(n_340),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1022),
.A2(n_696),
.B1(n_676),
.B2(n_675),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_995),
.A2(n_613),
.B(n_594),
.Y(n_1066)
);

AO31x2_ASAP7_75t_L g1067 ( 
.A1(n_970),
.A2(n_605),
.A3(n_600),
.B(n_616),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_894),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_898),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_997),
.A2(n_675),
.B(n_643),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_883),
.B(n_643),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_905),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_941),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_909),
.B(n_340),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1002),
.A2(n_538),
.B(n_540),
.C(n_552),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_887),
.A2(n_616),
.B(n_615),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_906),
.A2(n_374),
.B1(n_373),
.B2(n_371),
.Y(n_1077)
);

AOI21x1_ASAP7_75t_L g1078 ( 
.A1(n_997),
.A2(n_615),
.B(n_607),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_955),
.A2(n_451),
.B(n_448),
.C(n_445),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_915),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_SL g1081 ( 
.A(n_877),
.B(n_371),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_916),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_977),
.B(n_540),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_892),
.B(n_255),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_SL g1085 ( 
.A1(n_877),
.A2(n_416),
.B(n_414),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_982),
.A2(n_374),
.B(n_373),
.C(n_298),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_1024),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_998),
.B(n_279),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_887),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_957),
.B(n_405),
.Y(n_1090)
);

CKINVDCx16_ASAP7_75t_R g1091 ( 
.A(n_910),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1030),
.B(n_295),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_919),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_912),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_970),
.A2(n_300),
.B1(n_301),
.B2(n_313),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_879),
.B(n_318),
.Y(n_1096)
);

OR2x6_ASAP7_75t_L g1097 ( 
.A(n_869),
.B(n_405),
.Y(n_1097)
);

NAND3xp33_ASAP7_75t_L g1098 ( 
.A(n_965),
.B(n_411),
.C(n_410),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_873),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1019),
.A2(n_349),
.B1(n_362),
.B2(n_356),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_874),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_1028),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_985),
.A2(n_494),
.B1(n_411),
.B2(n_410),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1019),
.A2(n_406),
.B1(n_119),
.B2(n_187),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_941),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_896),
.B(n_1),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_913),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_R g1108 ( 
.A(n_914),
.B(n_186),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_957),
.B(n_971),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_863),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_971),
.B(n_494),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_871),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_987),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_SL g1114 ( 
.A1(n_911),
.A2(n_151),
.B(n_149),
.C(n_142),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_975),
.A2(n_2),
.B1(n_5),
.B2(n_8),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_975),
.B(n_5),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_999),
.B(n_8),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1013),
.B(n_11),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_923),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_909),
.B(n_137),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_L g1121 ( 
.A(n_876),
.B(n_11),
.C(n_17),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_902),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_962),
.A2(n_1031),
.B(n_1020),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_1028),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_923),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_925),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1020),
.A2(n_136),
.B(n_120),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_909),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_917),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_965),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_884),
.B(n_26),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1008),
.A2(n_115),
.B1(n_106),
.B2(n_105),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1011),
.A2(n_101),
.B(n_98),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_947),
.A2(n_84),
.B1(n_83),
.B2(n_79),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_969),
.B(n_28),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_895),
.B(n_30),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_924),
.A2(n_929),
.B(n_986),
.C(n_984),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_921),
.B(n_66),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1011),
.A2(n_1016),
.B(n_903),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_895),
.B(n_30),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_983),
.A2(n_31),
.B(n_32),
.C(n_34),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_925),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_993),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_890),
.B(n_36),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_921),
.B(n_74),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_921),
.B(n_64),
.Y(n_1146)
);

BUFx8_ASAP7_75t_SL g1147 ( 
.A(n_1000),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_943),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_869),
.B(n_37),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_926),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_967),
.B(n_40),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_948),
.B(n_40),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_993),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_861),
.B(n_45),
.Y(n_1154)
);

NAND2x1p5_ASAP7_75t_L g1155 ( 
.A(n_1011),
.B(n_46),
.Y(n_1155)
);

BUFx12f_ASAP7_75t_L g1156 ( 
.A(n_869),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_922),
.B(n_47),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_872),
.A2(n_1014),
.B1(n_1007),
.B2(n_1018),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_965),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_935),
.Y(n_1160)
);

BUFx12f_ASAP7_75t_L g1161 ( 
.A(n_908),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_932),
.A2(n_52),
.B(n_54),
.C(n_60),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_SL g1163 ( 
.A(n_928),
.B(n_60),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_927),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_881),
.A2(n_61),
.B1(n_922),
.B2(n_885),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_908),
.B(n_926),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_885),
.A2(n_928),
.B1(n_920),
.B2(n_888),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_927),
.Y(n_1168)
);

OR2x6_ASAP7_75t_L g1169 ( 
.A(n_908),
.B(n_960),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1011),
.B(n_1016),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1016),
.A2(n_903),
.B(n_1017),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_933),
.Y(n_1172)
);

O2A1O1Ixp5_ASAP7_75t_L g1173 ( 
.A1(n_1010),
.A2(n_1006),
.B(n_991),
.C(n_996),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_920),
.B(n_934),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_939),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_990),
.A2(n_904),
.B1(n_899),
.B2(n_968),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1034),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_SL g1178 ( 
.A(n_1091),
.B(n_931),
.C(n_953),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1036),
.A2(n_1016),
.B(n_864),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1055),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1038),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1044),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1174),
.B(n_934),
.Y(n_1183)
);

AO21x2_ASAP7_75t_L g1184 ( 
.A1(n_1123),
.A2(n_991),
.B(n_981),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1042),
.A2(n_1032),
.B(n_866),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1173),
.A2(n_981),
.B(n_1017),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1148),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1167),
.A2(n_1171),
.B(n_1032),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1148),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1058),
.B(n_1112),
.Y(n_1190)
);

O2A1O1Ixp5_ASAP7_75t_L g1191 ( 
.A1(n_1071),
.A2(n_972),
.B(n_900),
.C(n_942),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_1049),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1080),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1049),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1082),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1070),
.A2(n_1047),
.B(n_1046),
.Y(n_1196)
);

NOR2xp67_ASAP7_75t_L g1197 ( 
.A(n_1050),
.B(n_949),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1119),
.B(n_940),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1125),
.B(n_940),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1126),
.B(n_964),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1142),
.B(n_989),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1176),
.A2(n_972),
.A3(n_1026),
.B(n_1033),
.Y(n_1202)
);

AOI21xp33_ASAP7_75t_L g1203 ( 
.A1(n_1081),
.A2(n_979),
.B(n_963),
.Y(n_1203)
);

AND2x2_ASAP7_75t_SL g1204 ( 
.A(n_1163),
.B(n_868),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1176),
.A2(n_1015),
.B(n_978),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1053),
.A2(n_937),
.A3(n_889),
.B(n_882),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1052),
.A2(n_988),
.B(n_897),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1065),
.A2(n_1012),
.B(n_1029),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1164),
.B(n_1009),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1168),
.A2(n_936),
.B1(n_918),
.B2(n_945),
.Y(n_1210)
);

AO21x1_ASAP7_75t_L g1211 ( 
.A1(n_1081),
.A2(n_886),
.B(n_1025),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1084),
.A2(n_1151),
.B(n_1106),
.C(n_1037),
.Y(n_1212)
);

NAND3xp33_ASAP7_75t_L g1213 ( 
.A(n_1121),
.B(n_980),
.C(n_1023),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1041),
.A2(n_1021),
.B(n_1005),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1172),
.B(n_994),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1054),
.A2(n_878),
.B(n_1027),
.Y(n_1216)
);

OA22x2_ASAP7_75t_L g1217 ( 
.A1(n_1035),
.A2(n_961),
.B1(n_930),
.B2(n_880),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1131),
.A2(n_1027),
.B(n_943),
.C(n_966),
.Y(n_1218)
);

NAND3xp33_ASAP7_75t_L g1219 ( 
.A(n_1154),
.B(n_966),
.C(n_978),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_1072),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1040),
.A2(n_878),
.A3(n_966),
.B(n_978),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_1049),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1099),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1051),
.A2(n_1139),
.B(n_1094),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1076),
.A2(n_878),
.B(n_1015),
.Y(n_1225)
);

BUFx12f_ASAP7_75t_L g1226 ( 
.A(n_1124),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_1107),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1144),
.A2(n_1158),
.B(n_1141),
.C(n_1165),
.Y(n_1228)
);

AOI21xp33_ASAP7_75t_L g1229 ( 
.A1(n_1069),
.A2(n_1107),
.B(n_1092),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1089),
.A2(n_1094),
.B(n_1043),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1166),
.B(n_1109),
.Y(n_1231)
);

NAND3xp33_ASAP7_75t_SL g1232 ( 
.A(n_1163),
.B(n_1143),
.C(n_1153),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1150),
.B(n_1166),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1060),
.B(n_1039),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1075),
.A2(n_1061),
.A3(n_1157),
.B(n_1140),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1096),
.B(n_1088),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1056),
.A2(n_1136),
.B(n_1116),
.C(n_1039),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_L g1238 ( 
.A(n_1130),
.B(n_1159),
.C(n_1115),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1089),
.A2(n_1048),
.B(n_1170),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_SL g1240 ( 
.A1(n_1117),
.A2(n_1118),
.B(n_1152),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1048),
.A2(n_1083),
.B(n_1104),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_1085),
.A2(n_1098),
.B(n_1133),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1098),
.A2(n_1086),
.B(n_1062),
.C(n_1162),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1064),
.B(n_1122),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1095),
.A2(n_1090),
.B1(n_1135),
.B2(n_1149),
.Y(n_1245)
);

OR2x6_ASAP7_75t_L g1246 ( 
.A(n_1169),
.B(n_1097),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1050),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1090),
.B(n_1160),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1169),
.A2(n_1087),
.B1(n_1175),
.B2(n_1097),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_SL g1250 ( 
.A(n_1101),
.B(n_1113),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1120),
.A2(n_1074),
.B(n_1127),
.Y(n_1251)
);

O2A1O1Ixp5_ASAP7_75t_SL g1252 ( 
.A1(n_1095),
.A2(n_1057),
.B(n_1134),
.C(n_1100),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1073),
.B(n_1105),
.Y(n_1253)
);

NAND2xp33_ASAP7_75t_R g1254 ( 
.A(n_1108),
.B(n_1145),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1087),
.A2(n_1085),
.B(n_1155),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1128),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1067),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1111),
.A2(n_1114),
.B(n_1079),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1132),
.A2(n_1077),
.B(n_1063),
.C(n_1138),
.Y(n_1259)
);

AO32x2_ASAP7_75t_L g1260 ( 
.A1(n_1067),
.A2(n_1128),
.A3(n_1068),
.B1(n_1155),
.B2(n_1097),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_1138),
.Y(n_1261)
);

AO31x2_ASAP7_75t_L g1262 ( 
.A1(n_1067),
.A2(n_1103),
.A3(n_1149),
.B(n_1156),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1147),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1161),
.A2(n_1146),
.B(n_1129),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1102),
.A2(n_1093),
.B(n_1059),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1072),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1045),
.A2(n_1078),
.B(n_1066),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1174),
.B(n_875),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1036),
.A2(n_1176),
.A3(n_1167),
.B(n_1053),
.Y(n_1269)
);

O2A1O1Ixp5_ASAP7_75t_L g1270 ( 
.A1(n_1123),
.A2(n_875),
.B(n_974),
.C(n_907),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1055),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1036),
.A2(n_973),
.B(n_912),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1045),
.A2(n_1078),
.B(n_1066),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1174),
.B(n_875),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1036),
.A2(n_973),
.B(n_912),
.Y(n_1275)
);

AOI221x1_ASAP7_75t_L g1276 ( 
.A1(n_1176),
.A2(n_1165),
.B1(n_1167),
.B2(n_1036),
.C(n_1037),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1045),
.A2(n_1078),
.B(n_1066),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1110),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1036),
.A2(n_973),
.B(n_912),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1173),
.A2(n_1036),
.B(n_1171),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1137),
.A2(n_845),
.B(n_907),
.C(n_739),
.Y(n_1281)
);

AOI21xp33_ASAP7_75t_L g1282 ( 
.A1(n_1081),
.A2(n_845),
.B(n_883),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1036),
.A2(n_973),
.B(n_912),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1173),
.A2(n_1036),
.B(n_1176),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1174),
.B(n_875),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1036),
.A2(n_973),
.B(n_912),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1174),
.B(n_875),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1137),
.A2(n_845),
.B(n_907),
.C(n_739),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1034),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1176),
.A2(n_1119),
.B1(n_1126),
.B2(n_1125),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1173),
.A2(n_1036),
.B(n_1176),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1107),
.B(n_898),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1166),
.B(n_1109),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1036),
.A2(n_973),
.B(n_912),
.Y(n_1294)
);

O2A1O1Ixp5_ASAP7_75t_L g1295 ( 
.A1(n_1123),
.A2(n_875),
.B(n_974),
.C(n_907),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_SL g1296 ( 
.A1(n_1167),
.A2(n_1176),
.B(n_866),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1036),
.A2(n_973),
.B(n_912),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1058),
.B(n_381),
.Y(n_1298)
);

OAI21xp33_ASAP7_75t_L g1299 ( 
.A1(n_1106),
.A2(n_845),
.B(n_883),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1176),
.A2(n_1119),
.B1(n_1126),
.B2(n_1125),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1081),
.A2(n_526),
.B1(n_898),
.B2(n_1163),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1036),
.A2(n_1176),
.A3(n_1167),
.B(n_1053),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1174),
.B(n_875),
.Y(n_1303)
);

AOI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1123),
.A2(n_1078),
.B(n_1066),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1137),
.A2(n_845),
.B(n_907),
.C(n_739),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1137),
.A2(n_845),
.B(n_907),
.C(n_739),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1137),
.A2(n_845),
.B(n_907),
.C(n_739),
.Y(n_1307)
);

CKINVDCx14_ASAP7_75t_R g1308 ( 
.A(n_1102),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1148),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1107),
.B(n_883),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1174),
.B(n_875),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1174),
.B(n_875),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1174),
.B(n_875),
.Y(n_1313)
);

INVx5_ASAP7_75t_L g1314 ( 
.A(n_1089),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1174),
.B(n_875),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1231),
.B(n_1293),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1290),
.B(n_1300),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1193),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1177),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1182),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1227),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1299),
.A2(n_1238),
.B1(n_1282),
.B2(n_1301),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1292),
.B(n_1227),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1299),
.A2(n_1298),
.B1(n_1212),
.B2(n_1204),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1262),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1284),
.A2(n_1291),
.B(n_1288),
.C(n_1307),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1290),
.B(n_1300),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1238),
.A2(n_1284),
.B1(n_1291),
.B2(n_1261),
.Y(n_1328)
);

BUFx4f_ASAP7_75t_L g1329 ( 
.A(n_1194),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1281),
.A2(n_1306),
.B(n_1305),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1276),
.A2(n_1188),
.B(n_1196),
.Y(n_1331)
);

OA21x2_ASAP7_75t_L g1332 ( 
.A1(n_1186),
.A2(n_1304),
.B(n_1211),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1272),
.A2(n_1279),
.B(n_1275),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1200),
.B(n_1201),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1231),
.B(n_1293),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1278),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1283),
.A2(n_1286),
.B(n_1297),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1263),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1245),
.A2(n_1199),
.B1(n_1198),
.B2(n_1228),
.Y(n_1339)
);

NAND2x1p5_ASAP7_75t_L g1340 ( 
.A(n_1314),
.B(n_1192),
.Y(n_1340)
);

AO32x2_ASAP7_75t_L g1341 ( 
.A1(n_1249),
.A2(n_1269),
.A3(n_1302),
.B1(n_1202),
.B2(n_1210),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1232),
.A2(n_1203),
.B1(n_1236),
.B2(n_1315),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1257),
.A2(n_1241),
.A3(n_1179),
.B(n_1294),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1194),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1195),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1186),
.A2(n_1296),
.B(n_1224),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_1308),
.Y(n_1347)
);

BUFx2_ASAP7_75t_R g1348 ( 
.A(n_1234),
.Y(n_1348)
);

BUFx12f_ASAP7_75t_L g1349 ( 
.A(n_1226),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1289),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1252),
.A2(n_1295),
.B(n_1270),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1264),
.B(n_1246),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1271),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1181),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_R g1355 ( 
.A(n_1254),
.B(n_1250),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1223),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1208),
.A2(n_1216),
.B(n_1207),
.Y(n_1357)
);

NAND2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1314),
.B(n_1192),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1184),
.A2(n_1230),
.B(n_1258),
.Y(n_1359)
);

BUFx2_ASAP7_75t_SL g1360 ( 
.A(n_1220),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1280),
.A2(n_1184),
.B(n_1191),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1214),
.A2(n_1185),
.B(n_1225),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1243),
.B(n_1259),
.C(n_1310),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1214),
.A2(n_1255),
.B(n_1239),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1251),
.A2(n_1240),
.B(n_1280),
.Y(n_1365)
);

INVx6_ASAP7_75t_L g1366 ( 
.A(n_1222),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1268),
.B(n_1274),
.Y(n_1367)
);

AO21x2_ASAP7_75t_L g1368 ( 
.A1(n_1258),
.A2(n_1237),
.B(n_1219),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1210),
.A2(n_1218),
.A3(n_1285),
.B(n_1313),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1266),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1247),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1190),
.B(n_1245),
.Y(n_1372)
);

BUFx8_ASAP7_75t_L g1373 ( 
.A(n_1187),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1246),
.B(n_1205),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1183),
.A2(n_1312),
.B1(n_1311),
.B2(n_1303),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1242),
.A2(n_1197),
.B(n_1287),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1197),
.A2(n_1219),
.B(n_1215),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1256),
.A2(n_1209),
.B(n_1248),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1244),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1213),
.A2(n_1217),
.B(n_1233),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1246),
.B(n_1222),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1260),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1253),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1250),
.A2(n_1229),
.B1(n_1178),
.B2(n_1265),
.Y(n_1384)
);

INVx4_ASAP7_75t_SL g1385 ( 
.A(n_1262),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1221),
.A2(n_1206),
.B(n_1202),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1189),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1189),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1269),
.A2(n_1302),
.A3(n_1206),
.B(n_1202),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1260),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1221),
.A2(n_1269),
.B(n_1302),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1235),
.A2(n_1273),
.B(n_1267),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_SL g1393 ( 
.A1(n_1235),
.A2(n_1288),
.B(n_1305),
.C(n_1281),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1309),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1309),
.B(n_1314),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1284),
.A2(n_1291),
.B(n_1273),
.Y(n_1396)
);

O2A1O1Ixp5_ASAP7_75t_L g1397 ( 
.A1(n_1284),
.A2(n_875),
.B(n_1291),
.C(n_1282),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1263),
.Y(n_1398)
);

NAND2x1p5_ASAP7_75t_L g1399 ( 
.A(n_1314),
.B(n_1192),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1220),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1290),
.B(n_1300),
.Y(n_1401)
);

NOR4xp25_ASAP7_75t_L g1402 ( 
.A(n_1299),
.B(n_1282),
.C(n_1212),
.D(n_1281),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1290),
.B(n_1300),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1290),
.B(n_1300),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1267),
.A2(n_1277),
.B(n_1273),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1276),
.A2(n_1211),
.A3(n_1257),
.B(n_1188),
.Y(n_1406)
);

OAI21xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1282),
.A2(n_1176),
.B(n_1252),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1299),
.A2(n_1282),
.B1(n_1238),
.B2(n_1301),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1194),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1193),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1263),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1290),
.B(n_1300),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1231),
.B(n_1293),
.Y(n_1413)
);

NOR2x1_ASAP7_75t_R g1414 ( 
.A(n_1226),
.B(n_622),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1180),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1290),
.B(n_1300),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1282),
.A2(n_1299),
.B(n_1288),
.C(n_1281),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1299),
.A2(n_1282),
.B(n_1176),
.C(n_1284),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1299),
.B(n_1282),
.Y(n_1419)
);

NAND2x1p5_ASAP7_75t_L g1420 ( 
.A(n_1314),
.B(n_1192),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1267),
.A2(n_1277),
.B(n_1273),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1290),
.B(n_1300),
.Y(n_1422)
);

AO21x2_ASAP7_75t_L g1423 ( 
.A1(n_1284),
.A2(n_1291),
.B(n_1188),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1263),
.Y(n_1424)
);

NAND2x1p5_ASAP7_75t_L g1425 ( 
.A(n_1314),
.B(n_1192),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1267),
.A2(n_1277),
.B(n_1273),
.Y(n_1426)
);

BUFx2_ASAP7_75t_R g1427 ( 
.A(n_1234),
.Y(n_1427)
);

OAI211xp5_ASAP7_75t_L g1428 ( 
.A1(n_1299),
.A2(n_1282),
.B(n_845),
.C(n_678),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1292),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1284),
.A2(n_1291),
.B(n_1275),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1284),
.A2(n_1291),
.B(n_1275),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1204),
.A2(n_1081),
.B1(n_1176),
.B2(n_1238),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1263),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1284),
.A2(n_1291),
.B(n_1188),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1383),
.Y(n_1435)
);

AOI21x1_ASAP7_75t_SL g1436 ( 
.A1(n_1317),
.A2(n_1401),
.B(n_1327),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1430),
.A2(n_1431),
.B(n_1418),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1418),
.A2(n_1374),
.B(n_1322),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1432),
.A2(n_1324),
.B1(n_1408),
.B2(n_1363),
.Y(n_1439)
);

O2A1O1Ixp5_ASAP7_75t_L g1440 ( 
.A1(n_1330),
.A2(n_1351),
.B(n_1430),
.C(n_1431),
.Y(n_1440)
);

NOR2xp67_ASAP7_75t_L g1441 ( 
.A(n_1429),
.B(n_1379),
.Y(n_1441)
);

NAND2x1p5_ASAP7_75t_L g1442 ( 
.A(n_1352),
.B(n_1377),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1329),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1329),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1321),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1319),
.Y(n_1446)
);

O2A1O1Ixp5_ASAP7_75t_L g1447 ( 
.A1(n_1330),
.A2(n_1351),
.B(n_1326),
.C(n_1397),
.Y(n_1447)
);

AOI211xp5_ASAP7_75t_L g1448 ( 
.A1(n_1428),
.A2(n_1322),
.B(n_1402),
.C(n_1419),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1320),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1424),
.Y(n_1450)
);

O2A1O1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1428),
.A2(n_1419),
.B(n_1417),
.C(n_1397),
.Y(n_1451)
);

CKINVDCx14_ASAP7_75t_R g1452 ( 
.A(n_1424),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1323),
.B(n_1367),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1432),
.A2(n_1408),
.B(n_1328),
.C(n_1407),
.Y(n_1454)
);

OA21x2_ASAP7_75t_L g1455 ( 
.A1(n_1361),
.A2(n_1337),
.B(n_1386),
.Y(n_1455)
);

NOR2xp67_ASAP7_75t_L g1456 ( 
.A(n_1429),
.B(n_1400),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1328),
.A2(n_1404),
.B(n_1412),
.C(n_1422),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_SL g1458 ( 
.A(n_1373),
.Y(n_1458)
);

O2A1O1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1393),
.A2(n_1339),
.B(n_1375),
.C(n_1367),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1325),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1372),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1342),
.A2(n_1348),
.B1(n_1427),
.B2(n_1384),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1415),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1374),
.A2(n_1339),
.B(n_1375),
.Y(n_1464)
);

AND2x2_ASAP7_75t_SL g1465 ( 
.A(n_1403),
.B(n_1416),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1348),
.A2(n_1427),
.B1(n_1374),
.B2(n_1334),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1346),
.A2(n_1434),
.B(n_1423),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1340),
.A2(n_1399),
.B(n_1425),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1345),
.Y(n_1469)
);

CKINVDCx16_ASAP7_75t_R g1470 ( 
.A(n_1355),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1340),
.A2(n_1399),
.B(n_1425),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1391),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1316),
.B(n_1335),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1354),
.B(n_1336),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1353),
.A2(n_1370),
.B1(n_1360),
.B2(n_1350),
.Y(n_1475)
);

NOR2xp67_ASAP7_75t_L g1476 ( 
.A(n_1356),
.B(n_1318),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1358),
.A2(n_1420),
.B(n_1395),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1353),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1410),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1413),
.B(n_1387),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1388),
.B(n_1380),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1369),
.B(n_1355),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1338),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1361),
.A2(n_1392),
.B(n_1365),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1389),
.Y(n_1485)
);

BUFx8_ASAP7_75t_L g1486 ( 
.A(n_1349),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1371),
.B(n_1423),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1346),
.A2(n_1434),
.B(n_1359),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1378),
.B(n_1394),
.Y(n_1489)
);

A2O1A1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1364),
.A2(n_1376),
.B(n_1333),
.C(n_1382),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1341),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1389),
.B(n_1368),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1398),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1344),
.B(n_1409),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1389),
.B(n_1406),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1390),
.A2(n_1362),
.B(n_1341),
.C(n_1357),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1373),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1359),
.A2(n_1331),
.B(n_1396),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1389),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1411),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1341),
.B(n_1366),
.Y(n_1501)
);

O2A1O1Ixp5_ASAP7_75t_L g1502 ( 
.A1(n_1343),
.A2(n_1406),
.B(n_1331),
.C(n_1341),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1396),
.B(n_1366),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1347),
.A2(n_1358),
.B1(n_1433),
.B2(n_1332),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1406),
.B(n_1332),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1347),
.A2(n_1433),
.B(n_1414),
.C(n_1343),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1405),
.A2(n_1421),
.B(n_1426),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1343),
.A2(n_1291),
.B(n_1284),
.Y(n_1508)
);

O2A1O1Ixp5_ASAP7_75t_L g1509 ( 
.A1(n_1343),
.A2(n_875),
.B(n_1330),
.C(n_1291),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1385),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1428),
.B(n_1299),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1367),
.B(n_1429),
.Y(n_1512)
);

BUFx12f_ASAP7_75t_L g1513 ( 
.A(n_1349),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1323),
.B(n_1367),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1367),
.B(n_1429),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1323),
.B(n_1367),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1432),
.A2(n_1324),
.B1(n_883),
.B2(n_1204),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1353),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1418),
.A2(n_1288),
.B(n_1281),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1367),
.B(n_1429),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1319),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1319),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1432),
.A2(n_1324),
.B1(n_883),
.B2(n_1204),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1381),
.B(n_1352),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1367),
.B(n_1429),
.Y(n_1525)
);

CKINVDCx20_ASAP7_75t_R g1526 ( 
.A(n_1424),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1430),
.A2(n_1291),
.B(n_1284),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1418),
.A2(n_1288),
.B(n_1281),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1367),
.B(n_1429),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1507),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_SL g1531 ( 
.A1(n_1459),
.A2(n_1457),
.B(n_1517),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1485),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1505),
.B(n_1492),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1501),
.B(n_1491),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1488),
.A2(n_1498),
.B(n_1467),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1495),
.B(n_1496),
.Y(n_1536)
);

BUFx12f_ASAP7_75t_L g1537 ( 
.A(n_1486),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1442),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1460),
.Y(n_1539)
);

INVx4_ASAP7_75t_SL g1540 ( 
.A(n_1482),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1499),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1472),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1465),
.B(n_1457),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1446),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1490),
.B(n_1524),
.Y(n_1545)
);

AOI21xp33_ASAP7_75t_L g1546 ( 
.A1(n_1439),
.A2(n_1451),
.B(n_1448),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1437),
.B(n_1464),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1449),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1465),
.B(n_1527),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1440),
.B(n_1502),
.Y(n_1550)
);

OAI211xp5_ASAP7_75t_L g1551 ( 
.A1(n_1519),
.A2(n_1528),
.B(n_1511),
.C(n_1454),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1502),
.A2(n_1440),
.B(n_1447),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1469),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1487),
.B(n_1508),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1442),
.Y(n_1555)
);

CKINVDCx16_ASAP7_75t_R g1556 ( 
.A(n_1458),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1455),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1489),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1503),
.Y(n_1559)
);

INVx4_ASAP7_75t_L g1560 ( 
.A(n_1510),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1521),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1490),
.A2(n_1454),
.B(n_1438),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1509),
.B(n_1484),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1522),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1512),
.B(n_1515),
.Y(n_1565)
);

AO21x2_ASAP7_75t_L g1566 ( 
.A1(n_1511),
.A2(n_1504),
.B(n_1481),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1524),
.B(n_1479),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1523),
.B(n_1461),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1478),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1441),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1520),
.B(n_1525),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1450),
.Y(n_1572)
);

INVxp67_ASAP7_75t_SL g1573 ( 
.A(n_1529),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1476),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1518),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1474),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1453),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1514),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1516),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1538),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1564),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1545),
.B(n_1538),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1559),
.B(n_1445),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1539),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1544),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1573),
.B(n_1506),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1559),
.B(n_1475),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1554),
.B(n_1534),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1544),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1538),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1573),
.B(n_1456),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1533),
.B(n_1435),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1548),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1545),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1533),
.B(n_1463),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1550),
.B(n_1480),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1545),
.B(n_1494),
.Y(n_1597)
);

NOR2x1_ASAP7_75t_SL g1598 ( 
.A(n_1547),
.B(n_1466),
.Y(n_1598)
);

AO21x2_ASAP7_75t_L g1599 ( 
.A1(n_1535),
.A2(n_1462),
.B(n_1468),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1546),
.A2(n_1470),
.B1(n_1452),
.B2(n_1513),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1542),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1558),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1550),
.B(n_1473),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1546),
.A2(n_1486),
.B1(n_1497),
.B2(n_1526),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1550),
.B(n_1436),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1579),
.B(n_1471),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1542),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1531),
.A2(n_1458),
.B1(n_1443),
.B2(n_1444),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1530),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1604),
.A2(n_1551),
.B1(n_1600),
.B2(n_1543),
.C(n_1586),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1601),
.Y(n_1611)
);

OAI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1586),
.A2(n_1551),
.B1(n_1543),
.B2(n_1547),
.C(n_1549),
.Y(n_1612)
);

OAI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1608),
.A2(n_1547),
.B1(n_1549),
.B2(n_1568),
.C(n_1570),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1592),
.B(n_1556),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1601),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_L g1616 ( 
.A(n_1599),
.B(n_1562),
.Y(n_1616)
);

NAND4xp25_ASAP7_75t_L g1617 ( 
.A(n_1605),
.B(n_1568),
.C(n_1571),
.D(n_1565),
.Y(n_1617)
);

AOI222xp33_ASAP7_75t_L g1618 ( 
.A1(n_1598),
.A2(n_1537),
.B1(n_1565),
.B2(n_1571),
.C1(n_1578),
.C2(n_1572),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1590),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1607),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1588),
.B(n_1540),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1607),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1602),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1608),
.A2(n_1547),
.B1(n_1570),
.B2(n_1560),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1591),
.B(n_1578),
.Y(n_1625)
);

INVx8_ASAP7_75t_L g1626 ( 
.A(n_1582),
.Y(n_1626)
);

OA21x2_ASAP7_75t_L g1627 ( 
.A1(n_1609),
.A2(n_1535),
.B(n_1557),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1588),
.B(n_1540),
.Y(n_1628)
);

OAI31xp33_ASAP7_75t_L g1629 ( 
.A1(n_1605),
.A2(n_1574),
.A3(n_1575),
.B(n_1569),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1585),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1585),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1589),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1589),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1590),
.Y(n_1634)
);

NAND3xp33_ASAP7_75t_L g1635 ( 
.A(n_1583),
.B(n_1574),
.C(n_1552),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1597),
.A2(n_1562),
.B1(n_1566),
.B2(n_1599),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1594),
.B(n_1545),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1597),
.A2(n_1562),
.B1(n_1566),
.B2(n_1567),
.Y(n_1638)
);

OAI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1606),
.A2(n_1577),
.B1(n_1576),
.B2(n_1536),
.C(n_1555),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1593),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1592),
.B(n_1577),
.Y(n_1641)
);

OAI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1606),
.A2(n_1576),
.B1(n_1536),
.B2(n_1555),
.C(n_1558),
.Y(n_1642)
);

OAI33xp33_ASAP7_75t_L g1643 ( 
.A1(n_1581),
.A2(n_1536),
.A3(n_1532),
.B1(n_1541),
.B2(n_1553),
.B3(n_1561),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1580),
.Y(n_1644)
);

OAI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1595),
.A2(n_1576),
.B1(n_1555),
.B2(n_1558),
.C(n_1569),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1588),
.B(n_1540),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1630),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1621),
.B(n_1594),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1618),
.B(n_1582),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1635),
.B(n_1584),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1632),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1596),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1627),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1621),
.B(n_1603),
.Y(n_1654)
);

INVx4_ASAP7_75t_SL g1655 ( 
.A(n_1619),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1623),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1626),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1631),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1637),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1634),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1635),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1633),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_1637),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1640),
.Y(n_1664)
);

INVx4_ASAP7_75t_SL g1665 ( 
.A(n_1619),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_L g1666 ( 
.A(n_1636),
.B(n_1587),
.C(n_1595),
.D(n_1563),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1615),
.B(n_1596),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1620),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1658),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1658),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1660),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1652),
.B(n_1617),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1662),
.Y(n_1673)
);

NAND4xp25_ASAP7_75t_L g1674 ( 
.A(n_1666),
.B(n_1610),
.C(n_1612),
.D(n_1618),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1654),
.B(n_1628),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1661),
.A2(n_1616),
.B(n_1598),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1654),
.B(n_1646),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1656),
.Y(n_1678)
);

NOR3xp33_ASAP7_75t_SL g1679 ( 
.A(n_1666),
.B(n_1613),
.C(n_1617),
.Y(n_1679)
);

NOR2x1_ASAP7_75t_L g1680 ( 
.A(n_1660),
.B(n_1616),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1662),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1654),
.B(n_1646),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1662),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1647),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1647),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1653),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1655),
.B(n_1634),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1651),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1661),
.B(n_1622),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1653),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1664),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1655),
.B(n_1619),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_L g1693 ( 
.A(n_1649),
.B(n_1643),
.C(n_1624),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1655),
.B(n_1619),
.Y(n_1694)
);

NOR2x1_ASAP7_75t_R g1695 ( 
.A(n_1649),
.B(n_1537),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1655),
.B(n_1665),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1655),
.B(n_1619),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1665),
.B(n_1644),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1665),
.B(n_1638),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1665),
.B(n_1659),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1660),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1696),
.B(n_1665),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1696),
.B(n_1665),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1678),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1675),
.B(n_1665),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1679),
.B(n_1648),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1672),
.B(n_1667),
.Y(n_1707)
);

OAI21xp33_ASAP7_75t_L g1708 ( 
.A1(n_1674),
.A2(n_1650),
.B(n_1625),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1672),
.B(n_1641),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1673),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1673),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1681),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1693),
.B(n_1648),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1675),
.B(n_1659),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1677),
.B(n_1659),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1700),
.B(n_1663),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1686),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1674),
.B(n_1689),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1677),
.B(n_1663),
.Y(n_1719)
);

OAI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1676),
.A2(n_1657),
.B1(n_1650),
.B2(n_1663),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1681),
.Y(n_1721)
);

A2O1A1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1693),
.A2(n_1629),
.B(n_1614),
.C(n_1650),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1683),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1695),
.B(n_1537),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1683),
.Y(n_1725)
);

OR2x6_ASAP7_75t_L g1726 ( 
.A(n_1676),
.B(n_1477),
.Y(n_1726)
);

NOR5xp2_ASAP7_75t_L g1727 ( 
.A(n_1684),
.B(n_1645),
.C(n_1639),
.D(n_1642),
.E(n_1651),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1691),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1691),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1682),
.B(n_1657),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1682),
.B(n_1657),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1700),
.B(n_1648),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1689),
.B(n_1668),
.Y(n_1733)
);

AO21x1_ASAP7_75t_L g1734 ( 
.A1(n_1669),
.A2(n_1668),
.B(n_1629),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1685),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1706),
.B(n_1704),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1724),
.B(n_1695),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1702),
.B(n_1687),
.Y(n_1738)
);

INVx4_ASAP7_75t_L g1739 ( 
.A(n_1702),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1703),
.B(n_1687),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1703),
.B(n_1692),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1718),
.B(n_1669),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1735),
.Y(n_1743)
);

CKINVDCx16_ASAP7_75t_R g1744 ( 
.A(n_1724),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1708),
.A2(n_1562),
.B1(n_1699),
.B2(n_1566),
.Y(n_1745)
);

AND3x1_ASAP7_75t_L g1746 ( 
.A(n_1722),
.B(n_1680),
.C(n_1699),
.Y(n_1746)
);

AOI22x1_ASAP7_75t_L g1747 ( 
.A1(n_1727),
.A2(n_1701),
.B1(n_1671),
.B2(n_1500),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1732),
.B(n_1692),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1705),
.B(n_1680),
.Y(n_1749)
);

AO21x2_ASAP7_75t_L g1750 ( 
.A1(n_1734),
.A2(n_1670),
.B(n_1686),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1710),
.Y(n_1751)
);

NAND3x1_ASAP7_75t_L g1752 ( 
.A(n_1713),
.B(n_1697),
.C(n_1694),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1722),
.B(n_1701),
.Y(n_1753)
);

INVx3_ASAP7_75t_SL g1754 ( 
.A(n_1726),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1714),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1716),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1716),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1711),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1716),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1709),
.B(n_1483),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1732),
.B(n_1705),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1738),
.B(n_1730),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1746),
.B(n_1734),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1736),
.B(n_1707),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1747),
.A2(n_1720),
.B1(n_1726),
.B2(n_1566),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1755),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1743),
.B(n_1714),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_SL g1768 ( 
.A(n_1744),
.B(n_1694),
.Y(n_1768)
);

AOI33xp33_ASAP7_75t_L g1769 ( 
.A1(n_1745),
.A2(n_1712),
.A3(n_1721),
.B1(n_1723),
.B2(n_1725),
.B3(n_1729),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1755),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1755),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1743),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1738),
.B(n_1730),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1751),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1756),
.B(n_1715),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1751),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1758),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1758),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1756),
.B(n_1715),
.Y(n_1779)
);

O2A1O1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1753),
.A2(n_1726),
.B(n_1733),
.C(n_1688),
.Y(n_1780)
);

INVx2_ASAP7_75t_SL g1781 ( 
.A(n_1739),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1762),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1762),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1781),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1773),
.B(n_1739),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1768),
.B(n_1740),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1781),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1775),
.B(n_1739),
.Y(n_1788)
);

XNOR2x1_ASAP7_75t_L g1789 ( 
.A(n_1764),
.B(n_1747),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1766),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1763),
.B(n_1742),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1763),
.B(n_1742),
.Y(n_1792)
);

AOI222xp33_ASAP7_75t_L g1793 ( 
.A1(n_1791),
.A2(n_1765),
.B1(n_1772),
.B2(n_1767),
.C1(n_1746),
.C2(n_1779),
.Y(n_1793)
);

OAI211xp5_ASAP7_75t_L g1794 ( 
.A1(n_1791),
.A2(n_1765),
.B(n_1780),
.C(n_1739),
.Y(n_1794)
);

AOI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1792),
.A2(n_1750),
.B1(n_1759),
.B2(n_1757),
.C(n_1774),
.Y(n_1795)
);

OAI211xp5_ASAP7_75t_SL g1796 ( 
.A1(n_1792),
.A2(n_1769),
.B(n_1737),
.C(n_1776),
.Y(n_1796)
);

AOI211xp5_ASAP7_75t_L g1797 ( 
.A1(n_1786),
.A2(n_1788),
.B(n_1785),
.C(n_1754),
.Y(n_1797)
);

NOR3xp33_ASAP7_75t_L g1798 ( 
.A(n_1782),
.B(n_1744),
.C(n_1777),
.Y(n_1798)
);

AOI222xp33_ASAP7_75t_L g1799 ( 
.A1(n_1783),
.A2(n_1778),
.B1(n_1771),
.B2(n_1770),
.C1(n_1757),
.C2(n_1759),
.Y(n_1799)
);

AOI211x1_ASAP7_75t_L g1800 ( 
.A1(n_1790),
.A2(n_1740),
.B(n_1741),
.C(n_1761),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1787),
.B(n_1741),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1784),
.B(n_1761),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1802),
.B(n_1789),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1800),
.Y(n_1804)
);

BUFx2_ASAP7_75t_L g1805 ( 
.A(n_1801),
.Y(n_1805)
);

XOR2x2_ASAP7_75t_L g1806 ( 
.A(n_1798),
.B(n_1797),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1799),
.Y(n_1807)
);

OAI321xp33_ASAP7_75t_L g1808 ( 
.A1(n_1796),
.A2(n_1752),
.A3(n_1748),
.B1(n_1750),
.B2(n_1726),
.C(n_1754),
.Y(n_1808)
);

XNOR2x1_ASAP7_75t_L g1809 ( 
.A(n_1806),
.B(n_1493),
.Y(n_1809)
);

NOR3xp33_ASAP7_75t_L g1810 ( 
.A(n_1803),
.B(n_1795),
.C(n_1794),
.Y(n_1810)
);

XNOR2x1_ASAP7_75t_L g1811 ( 
.A(n_1807),
.B(n_1793),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1805),
.Y(n_1812)
);

NAND2xp33_ASAP7_75t_L g1813 ( 
.A(n_1804),
.B(n_1752),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1804),
.B(n_1748),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1812),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1814),
.Y(n_1816)
);

NOR4xp25_ASAP7_75t_L g1817 ( 
.A(n_1813),
.B(n_1808),
.C(n_1769),
.D(n_1750),
.Y(n_1817)
);

O2A1O1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1810),
.A2(n_1750),
.B(n_1754),
.C(n_1749),
.Y(n_1818)
);

AOI211xp5_ASAP7_75t_SL g1819 ( 
.A1(n_1811),
.A2(n_1749),
.B(n_1760),
.C(n_1728),
.Y(n_1819)
);

NOR2x1p5_ASAP7_75t_L g1820 ( 
.A(n_1815),
.B(n_1809),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1817),
.A2(n_1749),
.B1(n_1698),
.B2(n_1670),
.Y(n_1821)
);

XNOR2xp5_ASAP7_75t_L g1822 ( 
.A(n_1816),
.B(n_1749),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1822),
.B(n_1819),
.Y(n_1823)
);

OAI322xp33_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1818),
.A3(n_1821),
.B1(n_1820),
.B2(n_1733),
.C1(n_1717),
.C2(n_1690),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1824),
.A2(n_1717),
.B(n_1731),
.Y(n_1825)
);

CKINVDCx16_ASAP7_75t_R g1826 ( 
.A(n_1824),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1825),
.A2(n_1719),
.B(n_1731),
.Y(n_1827)
);

XNOR2xp5_ASAP7_75t_L g1828 ( 
.A(n_1826),
.B(n_1719),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1828),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1829),
.Y(n_1830)
);

INVxp67_ASAP7_75t_SL g1831 ( 
.A(n_1830),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1831),
.B(n_1827),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1832),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1833),
.A2(n_1686),
.B1(n_1690),
.B2(n_1697),
.C(n_1698),
.Y(n_1834)
);

AOI211xp5_ASAP7_75t_L g1835 ( 
.A1(n_1834),
.A2(n_1690),
.B(n_1443),
.C(n_1444),
.Y(n_1835)
);


endmodule