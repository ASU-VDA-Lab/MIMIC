module fake_jpeg_14514_n_181 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_181);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

INVx8_ASAP7_75t_SL g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

OR2x2_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_1),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_80),
.Y(n_89)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_1),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_54),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_76),
.B1(n_68),
.B2(n_62),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_68),
.B1(n_72),
.B2(n_71),
.Y(n_120)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_59),
.C(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_49),
.B(n_56),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_119),
.B(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_115),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_66),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_122),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_76),
.B1(n_55),
.B2(n_67),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_123),
.B1(n_4),
.B2(n_7),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_52),
.B1(n_55),
.B2(n_51),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_55),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_141),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_119),
.A2(n_67),
.B1(n_51),
.B2(n_61),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_130),
.B(n_139),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_21),
.B(n_23),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_120),
.B(n_118),
.Y(n_130)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_75),
.B(n_3),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_144),
.B1(n_9),
.B2(n_13),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_145),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_102),
.B(n_8),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_36),
.C(n_12),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_154),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_139),
.B1(n_142),
.B2(n_135),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_161),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_152),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_14),
.C(n_18),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_159),
.B(n_41),
.Y(n_168)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_25),
.C(n_29),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_30),
.B(n_34),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_151),
.C(n_146),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_167),
.B(n_158),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_159),
.B(n_155),
.C(n_43),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_170),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_164),
.A2(n_157),
.B1(n_126),
.B2(n_132),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_171),
.B1(n_163),
.B2(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_162),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_176),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_173),
.C(n_174),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_165),
.Y(n_181)
);


endmodule