module fake_jpeg_7297_n_59 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;

BUFx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_32),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_13),
.Y(n_45)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_1),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_26),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_4),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_28),
.B(n_22),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_28),
.B1(n_34),
.B2(n_36),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_42),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_11),
.C(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_45),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_14),
.C(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_16),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_17),
.C(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_49),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_44),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_53),
.B(n_51),
.C(n_44),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_52),
.B(n_50),
.C(n_37),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_52),
.Y(n_59)
);


endmodule