module real_aes_7355_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_1), .A2(n_149), .B(n_152), .C(n_232), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_2), .A2(n_178), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g509 ( .A(n_3), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_4), .B(n_208), .Y(n_207) );
AOI21xp33_ASAP7_75t_L g492 ( .A1(n_5), .A2(n_178), .B(n_493), .Y(n_492) );
AND2x6_ASAP7_75t_L g149 ( .A(n_6), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g245 ( .A(n_7), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_8), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_8), .B(n_44), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_9), .A2(n_177), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_10), .B(n_161), .Y(n_234) );
INVx1_ASAP7_75t_L g497 ( .A(n_11), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_12), .B(n_202), .Y(n_532) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_13), .A2(n_452), .B1(n_453), .B2(n_459), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_13), .Y(n_459) );
INVx1_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
INVx1_ASAP7_75t_L g544 ( .A(n_15), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_16), .A2(n_81), .B1(n_457), .B2(n_458), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_16), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_17), .A2(n_186), .B(n_267), .C(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_18), .B(n_208), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_19), .B(n_475), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_20), .B(n_178), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_21), .B(n_192), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_22), .A2(n_202), .B(n_253), .C(n_255), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_23), .A2(n_105), .B1(n_115), .B2(n_753), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_24), .B(n_208), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_25), .B(n_161), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_26), .A2(n_188), .B(n_269), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_27), .B(n_161), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g143 ( .A(n_28), .Y(n_143) );
INVx1_ASAP7_75t_L g215 ( .A(n_29), .Y(n_215) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_30), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_31), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_32), .B(n_161), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_33), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g184 ( .A(n_34), .Y(n_184) );
INVx1_ASAP7_75t_L g487 ( .A(n_35), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_36), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_36), .Y(n_454) );
INVx2_ASAP7_75t_L g147 ( .A(n_37), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_38), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_39), .A2(n_202), .B(n_203), .C(n_205), .Y(n_201) );
INVxp67_ASAP7_75t_L g187 ( .A(n_40), .Y(n_187) );
CKINVDCx14_ASAP7_75t_R g200 ( .A(n_41), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_42), .A2(n_152), .B(n_214), .C(n_218), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_43), .A2(n_149), .B(n_152), .C(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g114 ( .A(n_44), .Y(n_114) );
INVx1_ASAP7_75t_L g486 ( .A(n_45), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_46), .A2(n_163), .B(n_243), .C(n_244), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_47), .B(n_161), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_48), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_49), .Y(n_180) );
INVx1_ASAP7_75t_L g251 ( .A(n_50), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_51), .Y(n_488) );
AOI222xp33_ASAP7_75t_SL g449 ( .A1(n_52), .A2(n_450), .B1(n_451), .B2(n_460), .C1(n_746), .C2(n_749), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g432 ( .A1(n_53), .A2(n_62), .B1(n_433), .B2(n_434), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_53), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_54), .B(n_178), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_55), .A2(n_152), .B1(n_255), .B2(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_56), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_57), .Y(n_506) );
CKINVDCx14_ASAP7_75t_R g241 ( .A(n_58), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_59), .A2(n_205), .B(n_243), .C(n_496), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_60), .A2(n_123), .B1(n_124), .B2(n_437), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_60), .Y(n_437) );
INVx1_ASAP7_75t_L g494 ( .A(n_61), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_62), .Y(n_434) );
INVx1_ASAP7_75t_L g150 ( .A(n_63), .Y(n_150) );
INVx1_ASAP7_75t_L g140 ( .A(n_64), .Y(n_140) );
INVx1_ASAP7_75t_SL g204 ( .A(n_65), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_66), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g431 ( .A1(n_67), .A2(n_432), .B1(n_435), .B2(n_436), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_67), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_68), .B(n_208), .Y(n_257) );
INVx1_ASAP7_75t_L g156 ( .A(n_69), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_SL g474 ( .A1(n_70), .A2(n_205), .B(n_475), .C(n_476), .Y(n_474) );
INVxp67_ASAP7_75t_L g477 ( .A(n_71), .Y(n_477) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_73), .A2(n_178), .B(n_240), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_74), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_75), .A2(n_178), .B(n_264), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_76), .Y(n_490) );
INVx1_ASAP7_75t_L g550 ( .A(n_77), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_78), .A2(n_177), .B(n_179), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g212 ( .A(n_79), .Y(n_212) );
INVx1_ASAP7_75t_L g265 ( .A(n_80), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_81), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_82), .A2(n_149), .B(n_152), .C(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_83), .A2(n_178), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g268 ( .A(n_84), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_85), .B(n_185), .Y(n_521) );
INVx2_ASAP7_75t_L g138 ( .A(n_86), .Y(n_138) );
INVx1_ASAP7_75t_L g233 ( .A(n_87), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_88), .B(n_475), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_89), .A2(n_149), .B(n_152), .C(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g109 ( .A(n_90), .Y(n_109) );
OR2x2_ASAP7_75t_L g441 ( .A(n_90), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g461 ( .A(n_90), .B(n_443), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_91), .A2(n_152), .B(n_155), .C(n_165), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_92), .B(n_170), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_93), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_94), .A2(n_149), .B(n_152), .C(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_95), .Y(n_536) );
INVx1_ASAP7_75t_L g473 ( .A(n_96), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_97), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_98), .B(n_185), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_99), .B(n_136), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_100), .B(n_136), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_101), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g254 ( .A(n_102), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_103), .A2(n_178), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g754 ( .A(n_106), .Y(n_754) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g443 ( .A(n_108), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g745 ( .A(n_109), .B(n_443), .Y(n_745) );
NOR2x2_ASAP7_75t_L g748 ( .A(n_109), .B(n_442), .Y(n_748) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_448), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g752 ( .A(n_119), .Y(n_752) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_438), .B(n_445), .Y(n_121) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
XOR2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_431), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g460 ( .A1(n_125), .A2(n_461), .B1(n_462), .B2(n_743), .Y(n_460) );
INVx2_ASAP7_75t_L g750 ( .A(n_125), .Y(n_750) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_365), .Y(n_125) );
NAND5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_294), .C(n_324), .D(n_345), .E(n_351), .Y(n_126) );
AOI221xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_224), .B1(n_258), .B2(n_260), .C(n_271), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_221), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_193), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_SL g345 ( .A1(n_132), .A2(n_209), .B(n_346), .C(n_349), .Y(n_345) );
AND2x2_ASAP7_75t_L g415 ( .A(n_132), .B(n_210), .Y(n_415) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_171), .Y(n_132) );
AND2x2_ASAP7_75t_L g273 ( .A(n_133), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g277 ( .A(n_133), .B(n_274), .Y(n_277) );
OR2x2_ASAP7_75t_L g303 ( .A(n_133), .B(n_210), .Y(n_303) );
AND2x2_ASAP7_75t_L g305 ( .A(n_133), .B(n_196), .Y(n_305) );
AND2x2_ASAP7_75t_L g323 ( .A(n_133), .B(n_195), .Y(n_323) );
INVx1_ASAP7_75t_L g356 ( .A(n_133), .Y(n_356) );
INVx2_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
BUFx2_ASAP7_75t_L g223 ( .A(n_134), .Y(n_223) );
AND2x2_ASAP7_75t_L g259 ( .A(n_134), .B(n_196), .Y(n_259) );
AND2x2_ASAP7_75t_L g412 ( .A(n_134), .B(n_210), .Y(n_412) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_142), .B(n_167), .Y(n_134) );
INVx3_ASAP7_75t_L g208 ( .A(n_135), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_135), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_135), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_SL g523 ( .A(n_135), .B(n_524), .Y(n_523) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_136), .A2(n_471), .B(n_478), .Y(n_470) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_138), .B(n_139), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_151), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_144), .A2(n_170), .B(n_212), .C(n_213), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_144), .A2(n_230), .B(n_231), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_144), .A2(n_166), .B1(n_484), .B2(n_488), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_144), .A2(n_506), .B(n_507), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_144), .A2(n_550), .B(n_551), .Y(n_549) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
AND2x4_ASAP7_75t_L g178 ( .A(n_145), .B(n_149), .Y(n_178) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g256 ( .A(n_147), .Y(n_256) );
INVx1_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
INVx3_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
INVx1_ASAP7_75t_L g475 ( .A(n_148), .Y(n_475) );
INVx4_ASAP7_75t_SL g166 ( .A(n_149), .Y(n_166) );
BUFx3_ASAP7_75t_L g218 ( .A(n_149), .Y(n_218) );
INVx5_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx3_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_153), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_160), .C(n_162), .Y(n_155) );
O2A1O1Ixp5_ASAP7_75t_L g232 ( .A1(n_157), .A2(n_162), .B(n_233), .C(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g485 ( .A1(n_158), .A2(n_159), .B1(n_486), .B2(n_487), .Y(n_485) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g188 ( .A(n_159), .Y(n_188) );
INVx4_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
INVx2_ASAP7_75t_L g243 ( .A(n_161), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_162), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_162), .A2(n_553), .B(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g269 ( .A(n_164), .Y(n_269) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g179 ( .A1(n_166), .A2(n_180), .B(n_181), .C(n_182), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_166), .A2(n_181), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_SL g240 ( .A1(n_166), .A2(n_181), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g250 ( .A1(n_166), .A2(n_181), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_166), .A2(n_181), .B(n_265), .C(n_266), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_166), .A2(n_181), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_166), .A2(n_181), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_166), .A2(n_181), .B(n_541), .C(n_542), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVx1_ASAP7_75t_L g192 ( .A(n_169), .Y(n_192) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_169), .A2(n_528), .B(n_535), .Y(n_527) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_170), .A2(n_239), .B(n_246), .Y(n_238) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_170), .A2(n_539), .B(n_545), .Y(n_538) );
AND2x2_ASAP7_75t_L g293 ( .A(n_171), .B(n_194), .Y(n_293) );
OR2x2_ASAP7_75t_L g297 ( .A(n_171), .B(n_210), .Y(n_297) );
AND2x2_ASAP7_75t_L g322 ( .A(n_171), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g369 ( .A(n_171), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_171), .B(n_331), .Y(n_417) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_190), .Y(n_171) );
INVx1_ASAP7_75t_L g275 ( .A(n_172), .Y(n_275) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_172), .A2(n_549), .B(n_555), .Y(n_548) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_SL g517 ( .A1(n_173), .A2(n_518), .B(n_519), .Y(n_517) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_174), .A2(n_483), .B(n_489), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_174), .B(n_490), .Y(n_489) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_174), .A2(n_505), .B(n_512), .Y(n_504) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_176), .A2(n_191), .B(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_183), .B(n_189), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B1(n_187), .B2(n_188), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_185), .A2(n_215), .B(n_216), .C(n_217), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_185), .A2(n_509), .B(n_510), .C(n_511), .Y(n_508) );
INVx5_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_186), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_186), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_186), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_188), .B(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_188), .B(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_188), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g217 ( .A(n_189), .Y(n_217) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OAI322xp33_ASAP7_75t_L g418 ( .A1(n_193), .A2(n_354), .A3(n_377), .B1(n_398), .B2(n_419), .C1(n_421), .C2(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_194), .B(n_274), .Y(n_421) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_209), .Y(n_194) );
AND2x2_ASAP7_75t_L g222 ( .A(n_195), .B(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g290 ( .A(n_195), .B(n_210), .Y(n_290) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g331 ( .A(n_196), .B(n_210), .Y(n_331) );
AND2x2_ASAP7_75t_L g375 ( .A(n_196), .B(n_209), .Y(n_375) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_207), .Y(n_196) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_197), .A2(n_249), .B(n_257), .Y(n_248) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_197), .A2(n_263), .B(n_270), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_202), .B(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_206), .Y(n_533) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_208), .A2(n_492), .B(n_498), .Y(n_491) );
AND2x2_ASAP7_75t_L g258 ( .A(n_209), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g276 ( .A(n_209), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_209), .B(n_305), .Y(n_429) );
INVx3_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g221 ( .A(n_210), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_210), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g343 ( .A(n_210), .B(n_274), .Y(n_343) );
AND2x2_ASAP7_75t_L g370 ( .A(n_210), .B(n_305), .Y(n_370) );
OR2x2_ASAP7_75t_L g426 ( .A(n_210), .B(n_277), .Y(n_426) );
OR2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_219), .Y(n_210) );
INVx1_ASAP7_75t_SL g312 ( .A(n_221), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_222), .B(n_343), .Y(n_344) );
AND2x2_ASAP7_75t_L g378 ( .A(n_222), .B(n_368), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_222), .B(n_301), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_222), .B(n_423), .Y(n_422) );
OAI31xp33_ASAP7_75t_L g396 ( .A1(n_224), .A2(n_258), .A3(n_397), .B(n_399), .Y(n_396) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_237), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_225), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g379 ( .A(n_225), .B(n_314), .Y(n_379) );
OR2x2_ASAP7_75t_L g386 ( .A(n_225), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g398 ( .A(n_225), .B(n_287), .Y(n_398) );
CKINVDCx16_ASAP7_75t_R g225 ( .A(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g332 ( .A(n_226), .B(n_333), .Y(n_332) );
BUFx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g260 ( .A(n_227), .B(n_261), .Y(n_260) );
INVx4_ASAP7_75t_L g281 ( .A(n_227), .Y(n_281) );
AND2x2_ASAP7_75t_L g318 ( .A(n_227), .B(n_262), .Y(n_318) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_235), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_228), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_228), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_228), .B(n_437), .Y(n_555) );
AND2x2_ASAP7_75t_L g317 ( .A(n_237), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g387 ( .A(n_237), .Y(n_387) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_247), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_238), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g287 ( .A(n_238), .B(n_248), .Y(n_287) );
INVx2_ASAP7_75t_L g307 ( .A(n_238), .Y(n_307) );
AND2x2_ASAP7_75t_L g321 ( .A(n_238), .B(n_248), .Y(n_321) );
AND2x2_ASAP7_75t_L g328 ( .A(n_238), .B(n_284), .Y(n_328) );
BUFx3_ASAP7_75t_L g338 ( .A(n_238), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_238), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g283 ( .A(n_247), .Y(n_283) );
AND2x2_ASAP7_75t_L g291 ( .A(n_247), .B(n_281), .Y(n_291) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g261 ( .A(n_248), .B(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
INVx2_ASAP7_75t_L g511 ( .A(n_255), .Y(n_511) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_SL g298 ( .A(n_259), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_259), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_259), .B(n_368), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_260), .B(n_338), .Y(n_391) );
INVx1_ASAP7_75t_SL g425 ( .A(n_260), .Y(n_425) );
INVx1_ASAP7_75t_SL g333 ( .A(n_261), .Y(n_333) );
INVx1_ASAP7_75t_SL g284 ( .A(n_262), .Y(n_284) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_262), .Y(n_295) );
OR2x2_ASAP7_75t_L g306 ( .A(n_262), .B(n_281), .Y(n_306) );
AND2x2_ASAP7_75t_L g320 ( .A(n_262), .B(n_281), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_262), .B(n_310), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_276), .B(n_278), .C(n_289), .Y(n_271) );
AOI31xp33_ASAP7_75t_L g388 ( .A1(n_272), .A2(n_389), .A3(n_390), .B(n_391), .Y(n_388) );
AND2x2_ASAP7_75t_L g361 ( .A(n_273), .B(n_290), .Y(n_361) );
BUFx3_ASAP7_75t_L g301 ( .A(n_274), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_274), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g337 ( .A(n_274), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_274), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g292 ( .A(n_277), .Y(n_292) );
OAI222xp33_ASAP7_75t_L g401 ( .A1(n_277), .A2(n_402), .B1(n_405), .B2(n_406), .C1(n_407), .C2(n_408), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_285), .Y(n_278) );
INVx1_ASAP7_75t_L g407 ( .A(n_279), .Y(n_407) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_281), .B(n_284), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_281), .B(n_307), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_281), .B(n_282), .Y(n_377) );
INVx1_ASAP7_75t_L g428 ( .A(n_281), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_282), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g430 ( .A(n_282), .Y(n_430) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx2_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_284), .Y(n_353) );
AOI32xp33_ASAP7_75t_L g289 ( .A1(n_285), .A2(n_290), .A3(n_291), .B1(n_292), .B2(n_293), .Y(n_289) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_287), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g364 ( .A(n_287), .Y(n_364) );
OR2x2_ASAP7_75t_L g405 ( .A(n_287), .B(n_306), .Y(n_405) );
INVx1_ASAP7_75t_L g341 ( .A(n_288), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_290), .B(n_301), .Y(n_326) );
INVx3_ASAP7_75t_L g335 ( .A(n_290), .Y(n_335) );
AOI322xp5_ASAP7_75t_L g351 ( .A1(n_290), .A2(n_335), .A3(n_352), .B1(n_354), .B2(n_357), .C1(n_361), .C2(n_362), .Y(n_351) );
AND2x2_ASAP7_75t_L g327 ( .A(n_291), .B(n_328), .Y(n_327) );
INVxp67_ASAP7_75t_L g404 ( .A(n_291), .Y(n_404) );
A2O1A1O1Ixp25_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_299), .C(n_307), .D(n_308), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_295), .B(n_338), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g308 ( .A1(n_297), .A2(n_309), .B1(n_312), .B2(n_313), .C(n_316), .Y(n_308) );
INVx1_ASAP7_75t_SL g423 ( .A(n_297), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_304), .B(n_306), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_301), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI221xp5_ASAP7_75t_SL g393 ( .A1(n_303), .A2(n_387), .B1(n_394), .B2(n_395), .C(n_396), .Y(n_393) );
OAI222xp33_ASAP7_75t_L g424 ( .A1(n_304), .A2(n_425), .B1(n_426), .B2(n_427), .C1(n_429), .C2(n_430), .Y(n_424) );
AND2x2_ASAP7_75t_L g382 ( .A(n_305), .B(n_368), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_305), .A2(n_320), .B(n_367), .Y(n_394) );
INVx1_ASAP7_75t_L g408 ( .A(n_305), .Y(n_408) );
INVx2_ASAP7_75t_SL g311 ( .A(n_306), .Y(n_311) );
AND2x2_ASAP7_75t_L g314 ( .A(n_307), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_SL g348 ( .A(n_310), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_310), .B(n_320), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_311), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_311), .B(n_321), .Y(n_350) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI21xp5_ASAP7_75t_SL g316 ( .A1(n_317), .A2(n_319), .B(n_322), .Y(n_316) );
INVx1_ASAP7_75t_SL g334 ( .A(n_318), .Y(n_334) );
AND2x2_ASAP7_75t_L g381 ( .A(n_318), .B(n_364), .Y(n_381) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g420 ( .A(n_320), .B(n_338), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_321), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g406 ( .A(n_322), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B1(n_329), .B2(n_336), .C(n_339), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B1(n_334), .B2(n_335), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_333), .A2(n_340), .B1(n_342), .B2(n_344), .Y(n_339) );
OR2x2_ASAP7_75t_L g410 ( .A(n_334), .B(n_338), .Y(n_410) );
OR2x2_ASAP7_75t_L g413 ( .A(n_334), .B(n_348), .Y(n_413) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_355), .A2(n_410), .B1(n_411), .B2(n_413), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND3xp33_ASAP7_75t_SL g365 ( .A(n_366), .B(n_380), .C(n_392), .Y(n_365) );
AOI222xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B1(n_373), .B2(n_376), .C1(n_378), .C2(n_379), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_368), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g390 ( .A(n_370), .Y(n_390) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B1(n_383), .B2(n_385), .C(n_388), .Y(n_380) );
INVx1_ASAP7_75t_L g395 ( .A(n_381), .Y(n_395) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI21xp33_ASAP7_75t_L g414 ( .A1(n_385), .A2(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
NOR5xp2_ASAP7_75t_L g392 ( .A(n_393), .B(n_401), .C(n_409), .D(n_418), .E(n_424), .Y(n_392) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_432), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g447 ( .A(n_441), .Y(n_447) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_445), .B(n_449), .C(n_751), .Y(n_448) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_461), .A2(n_463), .B1(n_743), .B2(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_SL g463 ( .A(n_464), .B(n_680), .Y(n_463) );
NOR4xp25_ASAP7_75t_L g464 ( .A(n_465), .B(n_610), .C(n_641), .D(n_660), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g465 ( .A(n_466), .B(n_568), .C(n_583), .D(n_601), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_514), .B1(n_546), .B2(n_556), .C1(n_561), .C2(n_563), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_499), .Y(n_467) );
INVx1_ASAP7_75t_L g624 ( .A(n_468), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_479), .Y(n_468) );
AND2x2_ASAP7_75t_L g500 ( .A(n_469), .B(n_491), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_469), .B(n_503), .Y(n_653) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g560 ( .A(n_470), .B(n_481), .Y(n_560) );
AND2x2_ASAP7_75t_L g569 ( .A(n_470), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g595 ( .A(n_470), .Y(n_595) );
AND2x2_ASAP7_75t_L g616 ( .A(n_470), .B(n_481), .Y(n_616) );
BUFx2_ASAP7_75t_L g639 ( .A(n_470), .Y(n_639) );
AND2x2_ASAP7_75t_L g663 ( .A(n_470), .B(n_482), .Y(n_663) );
AND2x2_ASAP7_75t_L g727 ( .A(n_470), .B(n_491), .Y(n_727) );
AND2x2_ASAP7_75t_L g628 ( .A(n_479), .B(n_559), .Y(n_628) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_480), .B(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_491), .Y(n_480) );
OR2x2_ASAP7_75t_L g588 ( .A(n_481), .B(n_504), .Y(n_588) );
AND2x2_ASAP7_75t_L g600 ( .A(n_481), .B(n_559), .Y(n_600) );
BUFx2_ASAP7_75t_L g732 ( .A(n_481), .Y(n_732) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g502 ( .A(n_482), .B(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g582 ( .A(n_482), .B(n_504), .Y(n_582) );
AND2x2_ASAP7_75t_L g635 ( .A(n_482), .B(n_491), .Y(n_635) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_482), .Y(n_671) );
AND2x2_ASAP7_75t_L g558 ( .A(n_491), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_SL g570 ( .A(n_491), .Y(n_570) );
INVx2_ASAP7_75t_L g581 ( .A(n_491), .Y(n_581) );
BUFx2_ASAP7_75t_L g605 ( .A(n_491), .Y(n_605) );
AND2x2_ASAP7_75t_SL g662 ( .A(n_491), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
AOI332xp33_ASAP7_75t_L g583 ( .A1(n_500), .A2(n_584), .A3(n_588), .B1(n_589), .B2(n_593), .B3(n_596), .C1(n_597), .C2(n_599), .Y(n_583) );
NAND2x1_ASAP7_75t_L g668 ( .A(n_500), .B(n_559), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_500), .B(n_573), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_SL g601 ( .A1(n_501), .A2(n_602), .B(n_605), .C(n_606), .Y(n_601) );
AND2x2_ASAP7_75t_L g740 ( .A(n_501), .B(n_581), .Y(n_740) );
INVx3_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g637 ( .A(n_502), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g642 ( .A(n_502), .B(n_639), .Y(n_642) );
INVx1_ASAP7_75t_L g573 ( .A(n_503), .Y(n_573) );
AND2x2_ASAP7_75t_L g676 ( .A(n_503), .B(n_635), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_503), .B(n_616), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_503), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_503), .B(n_594), .Y(n_702) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g559 ( .A(n_504), .Y(n_559) );
OAI31xp33_ASAP7_75t_L g741 ( .A1(n_514), .A2(n_662), .A3(n_669), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_525), .Y(n_514) );
AND2x2_ASAP7_75t_L g546 ( .A(n_515), .B(n_547), .Y(n_546) );
NAND2x1_ASAP7_75t_SL g564 ( .A(n_515), .B(n_565), .Y(n_564) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_515), .Y(n_651) );
AND2x2_ASAP7_75t_L g656 ( .A(n_515), .B(n_567), .Y(n_656) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_516), .A2(n_569), .B(n_571), .C(n_574), .Y(n_568) );
OR2x2_ASAP7_75t_L g585 ( .A(n_516), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g598 ( .A(n_516), .Y(n_598) );
AND2x2_ASAP7_75t_L g604 ( .A(n_516), .B(n_548), .Y(n_604) );
INVx2_ASAP7_75t_L g622 ( .A(n_516), .Y(n_622) );
AND2x2_ASAP7_75t_L g633 ( .A(n_516), .B(n_587), .Y(n_633) );
AND2x2_ASAP7_75t_L g665 ( .A(n_516), .B(n_623), .Y(n_665) );
AND2x2_ASAP7_75t_L g669 ( .A(n_516), .B(n_592), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_516), .B(n_525), .Y(n_674) );
AND2x2_ASAP7_75t_L g708 ( .A(n_516), .B(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_516), .B(n_611), .Y(n_742) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_523), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_525), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g650 ( .A(n_525), .Y(n_650) );
AND2x2_ASAP7_75t_L g712 ( .A(n_525), .B(n_633), .Y(n_712) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_537), .Y(n_525) );
OR2x2_ASAP7_75t_L g566 ( .A(n_526), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g576 ( .A(n_526), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_526), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g684 ( .A(n_526), .Y(n_684) );
AND2x2_ASAP7_75t_L g701 ( .A(n_526), .B(n_548), .Y(n_701) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g592 ( .A(n_527), .B(n_537), .Y(n_592) );
AND2x2_ASAP7_75t_L g621 ( .A(n_527), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g632 ( .A(n_527), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_527), .B(n_587), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_534), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_533), .Y(n_530) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g547 ( .A(n_538), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g567 ( .A(n_538), .Y(n_567) );
AND2x2_ASAP7_75t_L g623 ( .A(n_538), .B(n_587), .Y(n_623) );
INVx1_ASAP7_75t_L g725 ( .A(n_546), .Y(n_725) );
INVx1_ASAP7_75t_L g729 ( .A(n_547), .Y(n_729) );
INVx2_ASAP7_75t_L g587 ( .A(n_548), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_558), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_558), .B(n_663), .Y(n_721) );
OR2x2_ASAP7_75t_L g562 ( .A(n_559), .B(n_560), .Y(n_562) );
INVx1_ASAP7_75t_SL g614 ( .A(n_559), .Y(n_614) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_565), .A2(n_618), .B1(n_620), .B2(n_624), .C(n_625), .Y(n_617) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g645 ( .A(n_566), .B(n_609), .Y(n_645) );
INVx2_ASAP7_75t_L g577 ( .A(n_567), .Y(n_577) );
INVx1_ASAP7_75t_L g603 ( .A(n_567), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_567), .B(n_587), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_567), .B(n_590), .Y(n_697) );
INVx1_ASAP7_75t_L g705 ( .A(n_567), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_569), .B(n_573), .Y(n_619) );
AND2x4_ASAP7_75t_L g594 ( .A(n_570), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g707 ( .A(n_573), .B(n_663), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_578), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_576), .B(n_608), .Y(n_607) );
INVxp67_ASAP7_75t_L g715 ( .A(n_577), .Y(n_715) );
INVxp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g615 ( .A(n_581), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g687 ( .A(n_581), .B(n_663), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_581), .B(n_600), .Y(n_693) );
AOI322xp5_ASAP7_75t_L g647 ( .A1(n_582), .A2(n_616), .A3(n_623), .B1(n_648), .B2(n_651), .C1(n_652), .C2(n_654), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_582), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g713 ( .A(n_585), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g659 ( .A(n_586), .Y(n_659) );
INVx2_ASAP7_75t_L g590 ( .A(n_587), .Y(n_590) );
INVx1_ASAP7_75t_L g649 ( .A(n_587), .Y(n_649) );
CKINVDCx16_ASAP7_75t_R g596 ( .A(n_588), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g685 ( .A(n_590), .B(n_598), .Y(n_685) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g597 ( .A(n_592), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g640 ( .A(n_592), .B(n_633), .Y(n_640) );
AND2x2_ASAP7_75t_L g644 ( .A(n_592), .B(n_604), .Y(n_644) );
OAI21xp33_ASAP7_75t_SL g654 ( .A1(n_593), .A2(n_655), .B(n_657), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g724 ( .A1(n_593), .A2(n_725), .B1(n_726), .B2(n_728), .Y(n_724) );
INVx3_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g599 ( .A(n_594), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_594), .B(n_614), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_596), .B(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g736 ( .A(n_603), .Y(n_736) );
INVx4_ASAP7_75t_L g609 ( .A(n_604), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_604), .B(n_631), .Y(n_679) );
INVx1_ASAP7_75t_SL g691 ( .A(n_605), .Y(n_691) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NOR2xp67_ASAP7_75t_L g704 ( .A(n_609), .B(n_705), .Y(n_704) );
OAI211xp5_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_612), .B(n_617), .C(n_634), .Y(n_610) );
OAI221xp5_ASAP7_75t_SL g730 ( .A1(n_612), .A2(n_650), .B1(n_729), .B2(n_731), .C(n_733), .Y(n_730) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_614), .B(n_727), .Y(n_726) );
OAI31xp33_ASAP7_75t_L g706 ( .A1(n_615), .A2(n_692), .A3(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g646 ( .A(n_616), .Y(n_646) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g696 ( .A(n_621), .Y(n_696) );
AND2x2_ASAP7_75t_L g709 ( .A(n_623), .B(n_632), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B(n_629), .Y(n_625) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVxp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_633), .B(n_736), .Y(n_735) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B(n_640), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI221xp5_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_643), .B1(n_645), .B2(n_646), .C(n_647), .Y(n_641) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_642), .A2(n_711), .B(n_713), .C(n_716), .Y(n_710) );
CKINVDCx16_ASAP7_75t_R g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_645), .B(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g672 ( .A(n_653), .Y(n_672) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g658 ( .A(n_656), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g700 ( .A(n_656), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B(n_666), .C(n_675), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_664), .A2(n_674), .B1(n_738), .B2(n_739), .C(n_741), .Y(n_737) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B1(n_670), .B2(n_673), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI21xp5_ASAP7_75t_SL g675 ( .A1(n_676), .A2(n_677), .B(n_678), .Y(n_675) );
INVx1_ASAP7_75t_SL g738 ( .A(n_677), .Y(n_738) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR4xp25_ASAP7_75t_L g680 ( .A(n_681), .B(n_710), .C(n_730), .D(n_737), .Y(n_680) );
OAI211xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_686), .B(n_688), .C(n_706), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
INVxp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
O2A1O1Ixp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_692), .B(n_694), .C(n_698), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g717 ( .A(n_695), .Y(n_717) );
OR2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
OR2x2_ASAP7_75t_L g728 ( .A(n_696), .B(n_729), .Y(n_728) );
OAI21xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_702), .B(n_703), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_720), .B2(n_722), .C(n_724), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_727), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
endmodule