module fake_jpeg_22303_n_121 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_20),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_26),
.B(n_13),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_48),
.B(n_24),
.C(n_21),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_30),
.A2(n_13),
.B1(n_24),
.B2(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_37),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_60),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_50),
.B1(n_31),
.B2(n_36),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_51),
.B1(n_14),
.B2(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_68),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_65),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_38),
.C(n_16),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_1),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_14),
.B1(n_51),
.B2(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_20),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_45),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_78),
.Y(n_92)
);

OAI32xp33_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_43),
.A3(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_94),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_65),
.B1(n_60),
.B2(n_56),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_11),
.C(n_8),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_76),
.C(n_77),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_96),
.B(n_97),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_71),
.B(n_73),
.C(n_77),
.D(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_74),
.C(n_83),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_83),
.B1(n_74),
.B2(n_28),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_84),
.B1(n_90),
.B2(n_85),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_93),
.B(n_91),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_44),
.B(n_22),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_72),
.B1(n_44),
.B2(n_63),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_109),
.B(n_44),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_72),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_100),
.B1(n_99),
.B2(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_104),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_106),
.B(n_105),
.Y(n_114)
);

XOR2x2_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_5),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_116),
.Y(n_118)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_116),
.C1(n_113),
.C2(n_112),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_2),
.C(n_3),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_118),
.Y(n_121)
);


endmodule