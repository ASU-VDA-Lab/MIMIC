module real_jpeg_14403_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_288;
wire n_215;
wire n_221;
wire n_249;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_3),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_3),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_3),
.B(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_3),
.B(n_32),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_3),
.B(n_77),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_4),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_4),
.B(n_44),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_4),
.B(n_30),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_4),
.B(n_50),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_4),
.B(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_4),
.B(n_53),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_4),
.B(n_32),
.Y(n_155)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_7),
.B(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_7),
.B(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_7),
.B(n_30),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_7),
.B(n_50),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_8),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_8),
.B(n_53),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_8),
.B(n_44),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_8),
.B(n_50),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_8),
.B(n_63),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_11),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_11),
.B(n_44),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_11),
.B(n_50),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_11),
.B(n_63),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_11),
.B(n_32),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_11),
.B(n_77),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_11),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_12),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_12),
.B(n_63),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_25),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_14),
.B(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_14),
.B(n_50),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_14),
.B(n_77),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_14),
.B(n_30),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_15),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_15),
.B(n_50),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_15),
.B(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_15),
.B(n_44),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_159),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_158),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_20),
.B(n_123),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.C(n_101),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_21),
.B(n_86),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_22),
.B(n_55),
.C(n_72),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.C(n_47),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_23),
.B(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_24),
.B(n_29),
.C(n_36),
.Y(n_100)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_29),
.B(n_155),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_29),
.A2(n_35),
.B1(n_154),
.B2(n_155),
.Y(n_236)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_33),
.B(n_46),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_33),
.B(n_67),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_37),
.A2(n_38),
.B1(n_47),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_38),
.A2(n_39),
.B(n_42),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_40),
.B(n_113),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_40),
.B(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_46),
.B(n_112),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_47),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.C(n_52),
.Y(n_47)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_48),
.B(n_49),
.CI(n_52),
.CON(n_104),
.SN(n_104)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_72),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_68),
.C(n_70),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.C(n_65),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_57),
.A2(n_58),
.B1(n_84),
.B2(n_85),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_57),
.A2(n_58),
.B1(n_62),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_69),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_SL g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_60),
.B(n_67),
.Y(n_253)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_62),
.Y(n_173)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_65),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_66),
.B(n_113),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_79),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_75),
.B(n_76),
.C(n_79),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_80),
.B(n_83),
.C(n_84),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_82),
.A2(n_83),
.B1(n_106),
.B2(n_107),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_84),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_84),
.A2(n_85),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_84),
.B(n_223),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_94),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_95),
.C(n_100),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_88),
.B(n_91),
.C(n_92),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.C(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_99),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_101),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_115),
.C(n_118),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_102),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.C(n_108),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_103),
.A2(n_104),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_104),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_105),
.B(n_108),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.C(n_114),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_111),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_157),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_147),
.B2(n_148),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_137),
.B2(n_138),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_145),
.B2(n_146),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_153),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_208),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_184),
.B(n_207),
.Y(n_161)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_162),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_182),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_182),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_170),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_167),
.B1(n_170),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_181),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_171),
.B(n_174),
.CI(n_181),
.CON(n_190),
.SN(n_190)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_179),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_175),
.A2(n_176),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_185),
.B(n_188),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_195),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_189),
.A2(n_190),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_190),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_191),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_287)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.C(n_201),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_197),
.B(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_200),
.B(n_201),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.C(n_205),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_289),
.C(n_290),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_283),
.B(n_288),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_268),
.B(n_282),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_238),
.B(n_267),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_225),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_213),
.B(n_225),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.C(n_222),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_228),
.B1(n_229),
.B2(n_231),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_214),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_264),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.CI(n_217),
.CON(n_214),
.SN(n_214)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_265),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_220),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_232),
.B2(n_237),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_231),
.C(n_237),
.Y(n_269)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_235),
.C(n_236),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_261),
.B(n_266),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_251),
.B(n_260),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_246),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_249),
.C(n_250),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_255),
.B(n_259),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_254),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_270),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_276),
.C(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_280),
.B2(n_281),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);


endmodule