module fake_jpeg_20077_n_274 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_33),
.Y(n_45)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_21),
.B1(n_29),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_50),
.B1(n_54),
.B2(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_21),
.B1(n_29),
.B2(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_15),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_31),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_60),
.B(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_21),
.B1(n_29),
.B2(n_24),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVxp67_ASAP7_75t_SL g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_57),
.Y(n_66)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_24),
.B1(n_31),
.B2(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_32),
.B1(n_36),
.B2(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_73),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_48),
.B1(n_50),
.B2(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_36),
.B1(n_32),
.B2(n_21),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_70),
.B1(n_52),
.B2(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_51),
.C(n_45),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_79),
.C(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_59),
.C(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_77),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_56),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_37),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_92),
.B1(n_64),
.B2(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_74),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_68),
.B1(n_55),
.B2(n_60),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_96),
.B1(n_66),
.B2(n_78),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_91),
.Y(n_111)
);

AO21x1_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_58),
.B(n_54),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_90),
.B1(n_93),
.B2(n_66),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_88),
.B(n_43),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_57),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_53),
.B1(n_57),
.B2(n_49),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_53),
.B1(n_46),
.B2(n_58),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_81),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_55),
.B1(n_60),
.B2(n_37),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_114),
.B1(n_96),
.B2(n_85),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_95),
.C(n_31),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_103),
.B1(n_108),
.B2(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_115),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_67),
.B(n_65),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_106),
.B(n_18),
.Y(n_147)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_76),
.B(n_75),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_63),
.B1(n_69),
.B2(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_38),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_74),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_74),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_119),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_66),
.B1(n_71),
.B2(n_77),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_17),
.B1(n_20),
.B2(n_18),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_89),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_118),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_97),
.B(n_88),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_23),
.B(n_16),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_132),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_90),
.B1(n_93),
.B2(n_97),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_86),
.B(n_61),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_23),
.B(n_16),
.Y(n_163)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_136),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_113),
.C(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_147),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_95),
.B1(n_61),
.B2(n_17),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVxp33_ASAP7_75t_SL g141 ( 
.A(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_142),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_20),
.B1(n_18),
.B2(n_14),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_61),
.C(n_14),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_31),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_31),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_31),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_164),
.B1(n_170),
.B2(n_127),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_156),
.Y(n_182)
);

NOR4xp25_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_19),
.C(n_16),
.D(n_20),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_153),
.B(n_166),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_14),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_161),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_169),
.B1(n_171),
.B2(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_23),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_163),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_30),
.B1(n_43),
.B2(n_2),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_126),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_167),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_19),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_128),
.A2(n_131),
.B1(n_122),
.B2(n_136),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_123),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_122),
.B1(n_146),
.B2(n_123),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_165),
.Y(n_203)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_135),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_179),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_135),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_134),
.C(n_129),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_185),
.C(n_187),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_134),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_181),
.B(n_30),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_127),
.C(n_25),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_148),
.B1(n_164),
.B2(n_3),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_38),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_158),
.C(n_149),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_19),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_154),
.A2(n_13),
.B1(n_30),
.B2(n_3),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_19),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_194),
.A2(n_157),
.B(n_160),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_197),
.A2(n_196),
.B(n_203),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_152),
.B(n_155),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_191),
.B(n_183),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_204),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_203),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_184),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_176),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_205),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_155),
.C(n_173),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_210),
.C(n_193),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_173),
.C(n_152),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_181),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_187),
.Y(n_216)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_215),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_219),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_189),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_197),
.C(n_198),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_223),
.C(n_202),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_185),
.C(n_178),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_228),
.B(n_235),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_234),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_200),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_200),
.C(n_199),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_0),
.B(n_1),
.Y(n_249)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_208),
.A3(n_202),
.B1(n_212),
.B2(n_211),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_237),
.A2(n_219),
.B1(n_225),
.B2(n_224),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_199),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_238),
.A2(n_220),
.B1(n_215),
.B2(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_245),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_231),
.A2(n_218),
.B(n_226),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_242),
.A2(n_0),
.B(n_3),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_217),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_249),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_213),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_248),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_216),
.B1(n_214),
.B2(n_13),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_19),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_232),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_254),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_255),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_236),
.B1(n_1),
.B2(n_3),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_13),
.Y(n_255)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_258),
.A2(n_257),
.A3(n_253),
.B1(n_252),
.B2(n_7),
.C1(n_9),
.C2(n_10),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_248),
.A3(n_25),
.B1(n_12),
.B2(n_22),
.C1(n_9),
.C2(n_4),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_256),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_262),
.Y(n_265)
);

NOR3xp33_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_4),
.C(n_5),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_5),
.B(n_6),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_265),
.A3(n_7),
.B1(n_10),
.B2(n_6),
.C1(n_12),
.C2(n_22),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_267),
.A2(n_264),
.B1(n_261),
.B2(n_259),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.C(n_25),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_12),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_271),
.B(n_12),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_12),
.B(n_6),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_7),
.B1(n_12),
.B2(n_257),
.Y(n_274)
);


endmodule