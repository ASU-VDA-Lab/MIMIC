module fake_jpeg_5910_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_1),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_6),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_18),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_2),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_10),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_15),
.C(n_4),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_14),
.B1(n_10),
.B2(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_21),
.B1(n_14),
.B2(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_34),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_33),
.Y(n_38)
);

NOR2xp67_ASAP7_75t_R g32 ( 
.A(n_29),
.B(n_3),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_29),
.B(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_25),
.B(n_11),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_40),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_35),
.C(n_11),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_42),
.B(n_45),
.C(n_46),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_41),
.Y(n_49)
);


endmodule