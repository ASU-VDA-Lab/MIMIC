module fake_jpeg_25555_n_341 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_9),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_39),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR3xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_0),
.C(n_1),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_45),
.Y(n_65)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_35),
.B1(n_34),
.B2(n_14),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_66),
.B1(n_41),
.B2(n_45),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_42),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_35),
.B1(n_34),
.B2(n_14),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_58),
.A2(n_42),
.B1(n_36),
.B2(n_49),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_64),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_34),
.B1(n_14),
.B2(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_37),
.B1(n_46),
.B2(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_99),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_41),
.B1(n_45),
.B2(n_43),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_81),
.Y(n_130)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_75),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_76),
.B(n_78),
.Y(n_128)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_79),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_60),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_36),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_87),
.C(n_93),
.Y(n_138)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_88),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_86),
.B(n_89),
.Y(n_150)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_51),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_67),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_45),
.B1(n_43),
.B2(n_40),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_110),
.B1(n_40),
.B2(n_20),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_93),
.Y(n_143)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_51),
.B(n_24),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_96),
.Y(n_133)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_69),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_104),
.B1(n_109),
.B2(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_23),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_62),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_23),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_27),
.Y(n_119)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_63),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_113),
.B1(n_101),
.B2(n_82),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_56),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_148),
.B1(n_86),
.B2(n_92),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_119),
.B(n_149),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_89),
.B(n_39),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_15),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_15),
.C(n_21),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_144),
.C(n_138),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_34),
.B1(n_20),
.B2(n_32),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_108),
.B1(n_101),
.B2(n_32),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_90),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_70),
.A2(n_32),
.B1(n_16),
.B2(n_28),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_142),
.B1(n_19),
.B2(n_16),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_77),
.A2(n_32),
.B1(n_16),
.B2(n_28),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_84),
.B(n_74),
.C(n_81),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_84),
.A2(n_83),
.B1(n_94),
.B2(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_85),
.B(n_26),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_72),
.Y(n_152)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_153),
.A2(n_173),
.B1(n_180),
.B2(n_181),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_154),
.B(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_112),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_157),
.B(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_163),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_133),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_164),
.A2(n_169),
.B1(n_185),
.B2(n_145),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_124),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_170),
.B(n_177),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_91),
.Y(n_166)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_149),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_167),
.Y(n_190)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

NAND2x1_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_90),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_21),
.Y(n_171)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_116),
.B1(n_117),
.B2(n_126),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_141),
.Y(n_200)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_117),
.B(n_73),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_90),
.B1(n_73),
.B2(n_76),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_176),
.B1(n_177),
.B2(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_19),
.B(n_29),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_130),
.A2(n_73),
.B1(n_30),
.B2(n_31),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_181)
);

OAI22x1_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_15),
.B1(n_21),
.B2(n_26),
.Y(n_182)
);

AOI22x1_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_135),
.B1(n_147),
.B2(n_15),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_29),
.B(n_28),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_184),
.B(n_136),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_R g184 ( 
.A(n_120),
.B(n_119),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_123),
.B(n_21),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_201),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_179),
.B(n_170),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_188),
.B(n_211),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_151),
.B(n_141),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_202),
.B1(n_204),
.B2(n_153),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_151),
.C(n_139),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_200),
.C(n_208),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_140),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_178),
.A2(n_121),
.B1(n_118),
.B2(n_137),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_121),
.B1(n_118),
.B2(n_137),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_206),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_142),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_33),
.B1(n_22),
.B2(n_18),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_147),
.C(n_135),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_154),
.A2(n_30),
.B(n_19),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_31),
.B(n_27),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_217),
.B(n_0),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_27),
.B(n_26),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_160),
.B(n_47),
.C(n_44),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_26),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_219),
.A2(n_225),
.B1(n_229),
.B2(n_188),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_216),
.A2(n_160),
.B1(n_169),
.B2(n_157),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_220),
.A2(n_245),
.B1(n_192),
.B2(n_210),
.Y(n_259)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_221),
.B(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_166),
.Y(n_224)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_164),
.B1(n_180),
.B2(n_155),
.Y(n_225)
);

AOI32xp33_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_181),
.A3(n_165),
.B1(n_156),
.B2(n_168),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_213),
.B(n_205),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_232),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_158),
.B1(n_175),
.B2(n_145),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_231),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_212),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_233),
.A2(n_246),
.B1(n_190),
.B2(n_192),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_234),
.B(n_235),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_33),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_207),
.A2(n_33),
.B1(n_22),
.B2(n_18),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_33),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_22),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_195),
.A2(n_47),
.A3(n_44),
.B1(n_22),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_237),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_47),
.B1(n_44),
.B2(n_3),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_247),
.A2(n_248),
.B1(n_255),
.B2(n_259),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_190),
.B1(n_187),
.B2(n_208),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_256),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_193),
.CI(n_195),
.CON(n_256),
.SN(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_193),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_267),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_265),
.B1(n_268),
.B2(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_200),
.C(n_198),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_269),
.C(n_242),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_219),
.A2(n_206),
.B1(n_201),
.B2(n_217),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_215),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_221),
.A2(n_215),
.B1(n_1),
.B2(n_3),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_246),
.C(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_273),
.A2(n_233),
.B1(n_256),
.B2(n_267),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_227),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_278),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_249),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_281),
.C(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_279),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_227),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_229),
.C(n_224),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_223),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_283),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_220),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_240),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_287),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_259),
.A2(n_225),
.B1(n_228),
.B2(n_233),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_265),
.B(n_233),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_0),
.C(n_3),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_296),
.B(n_284),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_261),
.B(n_260),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_280),
.B(n_5),
.Y(n_311)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_266),
.B1(n_248),
.B2(n_263),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_302),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_266),
.B1(n_250),
.B2(n_254),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_303),
.B(n_280),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_276),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_308),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_313),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_274),
.B1(n_278),
.B2(n_282),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_310),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_295),
.B(n_299),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_4),
.C(n_6),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_314),
.C(n_294),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_6),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_301),
.B1(n_292),
.B2(n_289),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_316),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_303),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_291),
.C(n_294),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_299),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_328),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_317),
.B1(n_320),
.B2(n_318),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_295),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_321),
.Y(n_333)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_324),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_333),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_314),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

AOI21x1_ASAP7_75t_SL g336 ( 
.A1(n_334),
.A2(n_330),
.B(n_325),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_335),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_325),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_321),
.B(n_309),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_10),
.Y(n_341)
);


endmodule