module fake_jpeg_2636_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_55),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_57),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_69),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_38),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_73),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_75),
.Y(n_94)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_40),
.B1(n_47),
.B2(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_40),
.Y(n_98)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_39),
.C(n_46),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_44),
.C(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_85),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_1),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_60),
.B(n_41),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_60),
.B1(n_40),
.B2(n_52),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_99),
.B(n_100),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_37),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_77),
.B(n_75),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_97),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_8),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_48),
.B(n_49),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_78),
.B1(n_84),
.B2(n_4),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_113),
.B1(n_114),
.B2(n_10),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_99),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_110),
.Y(n_128)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_1),
.CI(n_3),
.CON(n_110),
.SN(n_110)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_115),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_9),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_115),
.B(n_96),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_21),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_123),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_102),
.B1(n_109),
.B2(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_127),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_11),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_25),
.C(n_33),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_22),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_136),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_124),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_124),
.B1(n_131),
.B2(n_121),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_139),
.A2(n_120),
.B1(n_130),
.B2(n_12),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_125),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_141),
.A2(n_135),
.B(n_17),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_137),
.B1(n_128),
.B2(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_144),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_145),
.B(n_140),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_14),
.C(n_19),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_20),
.C(n_26),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_32),
.Y(n_152)
);


endmodule