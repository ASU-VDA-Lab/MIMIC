module fake_jpeg_27286_n_34 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_34);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_2),
.B(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_15),
.B(n_0),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_19),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_0),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_14),
.B(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_1),
.C(n_8),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_9),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_21),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_20),
.B1(n_24),
.B2(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_34)
);


endmodule