module fake_jpeg_4387_n_267 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_37),
.B(n_39),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_40),
.B(n_43),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_5),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_47),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_49),
.Y(n_100)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_52),
.B(n_53),
.Y(n_123)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_54),
.B(n_55),
.Y(n_125)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_32),
.B1(n_20),
.B2(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_56),
.A2(n_63),
.B1(n_99),
.B2(n_23),
.Y(n_103)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_18),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g107 ( 
.A(n_59),
.B(n_74),
.Y(n_107)
);

AND2x6_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

OA22x2_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_32),
.B1(n_17),
.B2(n_23),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_66),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_29),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_67),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_69),
.B(n_71),
.Y(n_101)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_30),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_41),
.B(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_27),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_76),
.B(n_78),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_40),
.A2(n_17),
.B1(n_34),
.B2(n_28),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_34),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_12),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_81),
.B(n_86),
.Y(n_119)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_39),
.B(n_12),
.Y(n_87)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_90),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_36),
.B(n_13),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_36),
.B(n_11),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_36),
.B(n_4),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_39),
.A2(n_23),
.B1(n_16),
.B2(n_19),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_116),
.B1(n_93),
.B2(n_88),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_61),
.A2(n_19),
.B1(n_14),
.B2(n_33),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_120),
.B1(n_93),
.B2(n_82),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_14),
.B1(n_24),
.B2(n_21),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_77),
.A2(n_33),
.B1(n_24),
.B2(n_21),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_74),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_139),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_82),
.B1(n_65),
.B2(n_51),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_135),
.B1(n_146),
.B2(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_57),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_132),
.B(n_142),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_126),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_84),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_137),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_88),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_0),
.Y(n_176)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_95),
.Y(n_140)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_145),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_62),
.B1(n_57),
.B2(n_94),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_101),
.B(n_124),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_21),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_157),
.B(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_86),
.B1(n_68),
.B2(n_67),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_154),
.A2(n_155),
.B1(n_7),
.B2(n_129),
.Y(n_184)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_4),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_24),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_117),
.B(n_110),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_160),
.A2(n_157),
.B(n_150),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_171),
.B(n_178),
.Y(n_190)
);

AO21x2_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_121),
.B(n_105),
.Y(n_163)
);

OAI22x1_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_164),
.B1(n_157),
.B2(n_150),
.Y(n_188)
);

OAI22x1_ASAP7_75t_SL g164 ( 
.A1(n_128),
.A2(n_121),
.B1(n_105),
.B2(n_102),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_110),
.B1(n_102),
.B2(n_111),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_141),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_111),
.B(n_1),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_131),
.B1(n_142),
.B2(n_152),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_0),
.C(n_1),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_179),
.C(n_168),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_181),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_136),
.A2(n_0),
.B(n_2),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_0),
.B(n_2),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_184),
.B(n_181),
.Y(n_205)
);

CKINVDCx12_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_3),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_193),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_206),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_196),
.B1(n_205),
.B2(n_166),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_164),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_149),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_198),
.B(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_134),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_154),
.B(n_141),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_163),
.B1(n_172),
.B2(n_166),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_153),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

AO22x2_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_163),
.B1(n_165),
.B2(n_160),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_207),
.A2(n_190),
.B1(n_203),
.B2(n_158),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_162),
.C(n_175),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_219),
.C(n_197),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_210),
.A2(n_194),
.B1(n_198),
.B2(n_199),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_196),
.B1(n_206),
.B2(n_158),
.Y(n_231)
);

OAI22x1_ASAP7_75t_SL g217 ( 
.A1(n_191),
.A2(n_175),
.B1(n_170),
.B2(n_167),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_192),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_183),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_189),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.C(n_228),
.Y(n_237)
);

XNOR2x2_ASAP7_75t_SL g226 ( 
.A(n_207),
.B(n_190),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_226),
.A2(n_227),
.B(n_207),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_204),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_195),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_218),
.C(n_215),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_207),
.B1(n_209),
.B2(n_229),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_233),
.Y(n_239)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_236),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_242),
.B(n_222),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_224),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_230),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_211),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_247),
.B(n_248),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_225),
.C(n_228),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_223),
.C(n_235),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_249),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_215),
.B(n_217),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_195),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_251),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_236),
.Y(n_253)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_SL g254 ( 
.A(n_246),
.B(n_237),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_255),
.B(n_239),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_250),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_255),
.C(n_256),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_261),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_174),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_265),
.A2(n_260),
.B(n_264),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_266),
.Y(n_267)
);


endmodule