module fake_jpeg_13780_n_175 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_152;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_14),
.B(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_33),
.B(n_45),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

CKINVDCx9p33_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_14),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_1),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_12),
.B(n_25),
.C(n_5),
.Y(n_85)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_26),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_54),
.Y(n_71)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_1),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_12),
.Y(n_55)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_15),
.B(n_2),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_3),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_60),
.A2(n_4),
.B1(n_7),
.B2(n_82),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_17),
.B1(n_28),
.B2(n_30),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_48),
.B1(n_41),
.B2(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_13),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_81),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_23),
.B1(n_16),
.B2(n_29),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_50),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_13),
.B1(n_23),
.B2(n_16),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_84),
.B1(n_76),
.B2(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_3),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_31),
.B(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_44),
.B(n_25),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_36),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_34),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_35),
.B1(n_42),
.B2(n_40),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_57),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_108),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_37),
.B1(n_38),
.B2(n_43),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_69),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_71),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_117),
.B(n_118),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_68),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_66),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_58),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_130),
.Y(n_142)
);

OAI22x1_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_109),
.B1(n_89),
.B2(n_103),
.Y(n_131)
);

OAI22x1_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_134),
.B1(n_126),
.B2(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_108),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_139),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_101),
.B1(n_105),
.B2(n_95),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_140),
.B1(n_124),
.B2(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_91),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_67),
.B1(n_78),
.B2(n_61),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_119),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_135),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_149),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_126),
.B(n_128),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_123),
.B(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_123),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_152),
.A2(n_146),
.B(n_144),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_145),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_137),
.B1(n_130),
.B2(n_113),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_154),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_133),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_155),
.C(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_122),
.B1(n_119),
.B2(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_162),
.C(n_111),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_119),
.C(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_151),
.B1(n_156),
.B2(n_121),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_124),
.B1(n_111),
.B2(n_125),
.Y(n_168)
);

AOI31xp33_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_159),
.A3(n_124),
.B(n_125),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_99),
.B1(n_80),
.B2(n_78),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_169),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_166),
.B1(n_165),
.B2(n_163),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_168),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_170),
.C(n_171),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_57),
.B(n_73),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_87),
.Y(n_175)
);


endmodule