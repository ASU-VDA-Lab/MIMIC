module fake_jpeg_25857_n_39 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_39);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_0),
.B(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_0),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_2),
.C(n_3),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_27),
.B(n_16),
.Y(n_31)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_2),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_18),
.B1(n_5),
.B2(n_8),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_30),
.B1(n_4),
.B2(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_18),
.B1(n_12),
.B2(n_14),
.Y(n_30)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_35),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

AO21x1_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_28),
.B(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_28),
.Y(n_39)
);


endmodule