module fake_ibex_262_n_1520 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_285, n_139, n_247, n_274, n_288, n_55, n_130, n_275, n_291, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_267, n_268, n_8, n_118, n_224, n_273, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_287, n_110, n_193, n_293, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_27, n_165, n_242, n_278, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_296, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_282, n_14, n_0, n_239, n_289, n_94, n_134, n_12, n_266, n_42, n_77, n_112, n_257, n_294, n_150, n_286, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_284, n_80, n_172, n_215, n_250, n_279, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_281, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_280, n_269, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_283, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_297, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_270, n_295, n_230, n_96, n_185, n_271, n_241, n_68, n_117, n_292, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_298, n_158, n_211, n_290, n_218, n_259, n_132, n_174, n_276, n_277, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_272, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1520);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_285;
input n_139;
input n_247;
input n_274;
input n_288;
input n_55;
input n_130;
input n_275;
input n_291;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_267;
input n_268;
input n_8;
input n_118;
input n_224;
input n_273;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_287;
input n_110;
input n_193;
input n_293;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_27;
input n_165;
input n_242;
input n_278;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_296;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_282;
input n_14;
input n_0;
input n_239;
input n_289;
input n_94;
input n_134;
input n_12;
input n_266;
input n_42;
input n_77;
input n_112;
input n_257;
input n_294;
input n_150;
input n_286;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_284;
input n_80;
input n_172;
input n_215;
input n_250;
input n_279;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_281;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_280;
input n_269;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_283;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_297;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_270;
input n_295;
input n_230;
input n_96;
input n_185;
input n_271;
input n_241;
input n_68;
input n_117;
input n_292;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_158;
input n_211;
input n_290;
input n_218;
input n_259;
input n_132;
input n_174;
input n_276;
input n_277;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_272;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1520;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_1509;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_1042;
wire n_822;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1477;
wire n_1184;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1495;
wire n_303;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_1340;
wire n_339;
wire n_348;
wire n_674;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_923;
wire n_642;
wire n_933;
wire n_1037;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_839;
wire n_768;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1415;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_1455;
wire n_484;
wire n_480;
wire n_354;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_581;
wire n_416;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g299 ( 
.A(n_213),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_289),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_86),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_150),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_144),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_46),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_175),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_1),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_86),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_33),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_163),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_138),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_115),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_151),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_37),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_132),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_198),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_141),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_221),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_201),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_109),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_134),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_23),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_41),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_215),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_160),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_252),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_27),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_143),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_166),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_154),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_148),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_176),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_52),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_155),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_292),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_199),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_41),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_298),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_69),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_233),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_261),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_71),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_1),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_38),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_229),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_205),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_217),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_245),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_243),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_142),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_18),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_67),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_12),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_207),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_260),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_259),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_120),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_188),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_129),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_227),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_76),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_22),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_250),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_220),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_280),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_109),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_177),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_178),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_234),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_279),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_152),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_285),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_277),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_262),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_79),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_44),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_90),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_212),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_208),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_94),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_275),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_173),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_288),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_77),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_20),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_237),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_62),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_195),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_190),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_125),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_225),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_102),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_7),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_78),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_46),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_77),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_284),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_258),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_294),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_104),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_264),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_265),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_135),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_297),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_219),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_270),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_222),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_196),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_290),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_111),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_267),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_113),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_80),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_183),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_191),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_197),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_56),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_286),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_249),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_247),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_51),
.Y(n_422)
);

BUFx8_ASAP7_75t_SL g423 ( 
.A(n_18),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_10),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_283),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_76),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_127),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_105),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_204),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_99),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_296),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_22),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_8),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_124),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_228),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_232),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_218),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_216),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_291),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_193),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_230),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_210),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_203),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_45),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_157),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_253),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_107),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_47),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_60),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_194),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_74),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_254),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_118),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_164),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_192),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_251),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_37),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_209),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_73),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_73),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_246),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_244),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_238),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_170),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_149),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_242),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_206),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_293),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_272),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_295),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_248),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_202),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_74),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_161),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_52),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_78),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_145),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_269),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_256),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_189),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_273),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_39),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_235),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_159),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_276),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_282),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_28),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_255),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_90),
.Y(n_489)
);

BUFx8_ASAP7_75t_SL g490 ( 
.A(n_153),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_271),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_47),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_168),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_278),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_241),
.Y(n_495)
);

BUFx2_ASAP7_75t_SL g496 ( 
.A(n_110),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_136),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_35),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_181),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_111),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_107),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_231),
.Y(n_502)
);

BUFx10_ASAP7_75t_L g503 ( 
.A(n_34),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_69),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_274),
.Y(n_505)
);

BUFx8_ASAP7_75t_SL g506 ( 
.A(n_126),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_200),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_6),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_223),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_13),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_236),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_65),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_158),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_239),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_6),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_287),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_266),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_116),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_240),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_156),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_36),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_263),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_131),
.Y(n_523)
);

CKINVDCx14_ASAP7_75t_R g524 ( 
.A(n_133),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_121),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_257),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_179),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_214),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_95),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_211),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_224),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_93),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_226),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_103),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_477),
.Y(n_535)
);

INVxp67_ASAP7_75t_SL g536 ( 
.A(n_422),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g537 ( 
.A(n_362),
.B(n_385),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_372),
.B(n_0),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_490),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_490),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_317),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_374),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_506),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_422),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_423),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_305),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_506),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_305),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_429),
.B(n_0),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_300),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_423),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_324),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_384),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_391),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_402),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_501),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_394),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_353),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_406),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_414),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_308),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_408),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_330),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_341),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_309),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_353),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_419),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_328),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_451),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_340),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_408),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_507),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g574 ( 
.A(n_408),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_345),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_451),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_503),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_352),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_378),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_439),
.B(n_2),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_482),
.Y(n_581)
);

INVxp33_ASAP7_75t_SL g582 ( 
.A(n_301),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_393),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_411),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_311),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_520),
.Y(n_586)
);

INVxp67_ASAP7_75t_SL g587 ( 
.A(n_520),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_503),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_520),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_424),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_311),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_426),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_366),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_447),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_482),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_366),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_448),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_318),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_463),
.B(n_2),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_521),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_459),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_476),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_307),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_489),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_299),
.B(n_3),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_503),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_504),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_R g608 ( 
.A(n_524),
.B(n_114),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_515),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_375),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_375),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_532),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_380),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_392),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_524),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_586),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_547),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_559),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_547),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_598),
.Y(n_620)
);

NOR2x1_ASAP7_75t_L g621 ( 
.A(n_614),
.B(n_303),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_586),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_561),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_563),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_572),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_603),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_R g627 ( 
.A(n_539),
.B(n_380),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_574),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_540),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_587),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_535),
.B(n_318),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_589),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_598),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_543),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_546),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_548),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_536),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_551),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_554),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_544),
.B(n_315),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_541),
.B(n_316),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_606),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_537),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_550),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_562),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_559),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_567),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_557),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_566),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_542),
.B(n_615),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_569),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_571),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_567),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_575),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_578),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_577),
.B(n_337),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_579),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_582),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_582),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_555),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_588),
.B(n_337),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_558),
.B(n_612),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_615),
.B(n_392),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_564),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_583),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_584),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_590),
.B(n_592),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_594),
.B(n_315),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_597),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_601),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_602),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_604),
.B(n_342),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_556),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_607),
.B(n_355),
.Y(n_674)
);

AND2x6_ASAP7_75t_L g675 ( 
.A(n_538),
.B(n_342),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_609),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_570),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_549),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_580),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_599),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_570),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_605),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_608),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_565),
.B(n_355),
.Y(n_684)
);

CKINVDCx8_ASAP7_75t_R g685 ( 
.A(n_560),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_568),
.B(n_364),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_573),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_585),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_591),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_593),
.Y(n_690)
);

CKINVDCx8_ASAP7_75t_R g691 ( 
.A(n_596),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_610),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_553),
.Y(n_693)
);

BUFx8_ASAP7_75t_L g694 ( 
.A(n_545),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_611),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_553),
.Y(n_696)
);

AND2x6_ASAP7_75t_L g697 ( 
.A(n_613),
.B(n_349),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_545),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_552),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_552),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_576),
.B(n_304),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_576),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_581),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_SL g704 ( 
.A1(n_581),
.A2(n_321),
.B1(n_323),
.B2(n_314),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_595),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_595),
.B(n_364),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_600),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_600),
.B(n_407),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_606),
.B(n_392),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_603),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_586),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_559),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_603),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_547),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_586),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_547),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_586),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_586),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_547),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_586),
.B(n_407),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_603),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_586),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_547),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_586),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_606),
.B(n_466),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_563),
.B(n_334),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_R g727 ( 
.A(n_547),
.B(n_410),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_606),
.B(n_466),
.Y(n_728)
);

XOR2xp5_ASAP7_75t_L g729 ( 
.A(n_553),
.B(n_410),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_586),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_586),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_547),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_603),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_586),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_586),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_614),
.B(n_319),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_547),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_586),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_547),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_586),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_606),
.B(n_466),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_614),
.B(n_349),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_586),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_R g744 ( 
.A(n_547),
.B(n_453),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_547),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_586),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_547),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_586),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_598),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_547),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_586),
.B(n_454),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_547),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_547),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_623),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_658),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_678),
.B(n_443),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_679),
.B(n_502),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_662),
.B(n_302),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_680),
.B(n_306),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_633),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_618),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_722),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_656),
.B(n_465),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_633),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_738),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_633),
.Y(n_766)
);

BUFx10_ASAP7_75t_L g767 ( 
.A(n_662),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_738),
.Y(n_768)
);

BUFx10_ASAP7_75t_L g769 ( 
.A(n_642),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_626),
.B(n_338),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_738),
.Y(n_771)
);

AND2x6_ASAP7_75t_L g772 ( 
.A(n_709),
.B(n_398),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_740),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_659),
.B(n_496),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_669),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_725),
.B(n_398),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_683),
.B(n_310),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_644),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_644),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_682),
.B(n_312),
.Y(n_780)
);

AND2x6_ASAP7_75t_L g781 ( 
.A(n_728),
.B(n_741),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_710),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_635),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_636),
.Y(n_784)
);

AND3x4_ASAP7_75t_L g785 ( 
.A(n_699),
.B(n_521),
.C(n_397),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_740),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_648),
.Y(n_787)
);

AND2x6_ASAP7_75t_L g788 ( 
.A(n_621),
.B(n_403),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_733),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_648),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_682),
.B(n_313),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_625),
.A2(n_488),
.B1(n_519),
.B2(n_465),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_648),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_656),
.B(n_488),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_628),
.B(n_322),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_652),
.Y(n_796)
);

OAI22xp33_ASAP7_75t_L g797 ( 
.A1(n_706),
.A2(n_519),
.B1(n_401),
.B2(n_395),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_654),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_713),
.B(n_343),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_657),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_630),
.B(n_325),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_748),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_676),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_641),
.A2(n_354),
.B1(n_363),
.B2(n_344),
.Y(n_804)
);

INVx6_ASAP7_75t_L g805 ( 
.A(n_694),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_632),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_637),
.B(n_326),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_726),
.B(n_327),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_720),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_672),
.B(n_329),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_672),
.B(n_331),
.Y(n_811)
);

AND2x6_ASAP7_75t_SL g812 ( 
.A(n_698),
.B(n_320),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_646),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_720),
.Y(n_814)
);

AND2x6_ASAP7_75t_L g815 ( 
.A(n_663),
.B(n_403),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_661),
.B(n_333),
.Y(n_816)
);

NOR2x1p5_ASAP7_75t_L g817 ( 
.A(n_617),
.B(n_619),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_647),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_689),
.B(n_332),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_721),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_629),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_620),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_742),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_634),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_664),
.B(n_367),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_684),
.B(n_336),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_706),
.A2(n_534),
.B1(n_377),
.B2(n_381),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_749),
.Y(n_828)
);

NOR2x1p5_ASAP7_75t_L g829 ( 
.A(n_714),
.B(n_376),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_727),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_708),
.B(n_386),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_661),
.B(n_388),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_684),
.B(n_686),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_708),
.B(n_396),
.Y(n_834)
);

INVx5_ASAP7_75t_L g835 ( 
.A(n_697),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_631),
.B(n_500),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_631),
.A2(n_667),
.B1(n_736),
.B2(n_645),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_751),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_742),
.B(n_339),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_616),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_649),
.B(n_413),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_687),
.B(n_347),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_651),
.Y(n_843)
);

AND2x4_ASAP7_75t_SL g844 ( 
.A(n_689),
.B(n_346),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_744),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_622),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_655),
.B(n_348),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_643),
.B(n_418),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_665),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_666),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_711),
.Y(n_851)
);

BUFx10_ASAP7_75t_L g852 ( 
.A(n_716),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_670),
.B(n_428),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_671),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_640),
.B(n_430),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_715),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_717),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_640),
.B(n_432),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_718),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_693),
.B(n_433),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_697),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_690),
.B(n_350),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_627),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_701),
.B(n_444),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_696),
.B(n_702),
.Y(n_865)
);

AND2x6_ASAP7_75t_L g866 ( 
.A(n_724),
.B(n_351),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_638),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_675),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_668),
.B(n_449),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_730),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_731),
.B(n_356),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_734),
.B(n_357),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_735),
.B(n_359),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_743),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_746),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_668),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_675),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_692),
.B(n_360),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_674),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_674),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_639),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_688),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_697),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_697),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_695),
.B(n_457),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_753),
.Y(n_886)
);

HAxp5_ASAP7_75t_SL g887 ( 
.A(n_729),
.B(n_361),
.CON(n_887),
.SN(n_887)
);

INVx5_ASAP7_75t_L g888 ( 
.A(n_689),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_685),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_704),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_719),
.B(n_368),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_723),
.B(n_369),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_660),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_705),
.B(n_370),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_703),
.B(n_371),
.Y(n_895)
);

AND2x2_ASAP7_75t_SL g896 ( 
.A(n_700),
.B(n_694),
.Y(n_896)
);

AND2x6_ASAP7_75t_L g897 ( 
.A(n_691),
.B(n_365),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_673),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_732),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_737),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_739),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_745),
.Y(n_902)
);

AND3x1_ASAP7_75t_L g903 ( 
.A(n_653),
.B(n_681),
.C(n_677),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_747),
.B(n_750),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_752),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_707),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_712),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_623),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_626),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_656),
.B(n_460),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_722),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_624),
.A2(n_405),
.B1(n_434),
.B2(n_399),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_624),
.A2(n_446),
.B1(n_455),
.B2(n_440),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_626),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_623),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_722),
.Y(n_916)
);

AO21x2_ASAP7_75t_L g917 ( 
.A1(n_720),
.A2(n_464),
.B(n_462),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_624),
.B(n_373),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_623),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_678),
.B(n_379),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_727),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_624),
.B(n_382),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_626),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_623),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_623),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_722),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_678),
.B(n_383),
.Y(n_927)
);

NAND2x1p5_ASAP7_75t_L g928 ( 
.A(n_658),
.B(n_467),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_662),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_662),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_662),
.B(n_473),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_662),
.B(n_475),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_623),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_727),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_662),
.B(n_387),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_722),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_656),
.B(n_487),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_722),
.Y(n_938)
);

BUFx4f_ASAP7_75t_L g939 ( 
.A(n_697),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_662),
.B(n_492),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_624),
.B(n_389),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_722),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_722),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_656),
.B(n_498),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_650),
.B(n_510),
.C(n_508),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_678),
.B(n_390),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_623),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_623),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_722),
.Y(n_949)
);

XOR2xp5_ASAP7_75t_L g950 ( 
.A(n_887),
.B(n_512),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_929),
.B(n_529),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_SL g952 ( 
.A(n_820),
.B(n_400),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_846),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_876),
.Y(n_954)
);

NOR2x1p5_ASAP7_75t_L g955 ( 
.A(n_889),
.B(n_404),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_930),
.A2(n_833),
.B1(n_858),
.B2(n_855),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_909),
.B(n_3),
.Y(n_957)
);

OR2x6_ASAP7_75t_L g958 ( 
.A(n_805),
.B(n_889),
.Y(n_958)
);

AND2x6_ASAP7_75t_SL g959 ( 
.A(n_774),
.B(n_470),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_880),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_767),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_846),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_879),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_767),
.B(n_409),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_806),
.Y(n_965)
);

NAND2xp33_ASAP7_75t_SL g966 ( 
.A(n_861),
.B(n_412),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_856),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_856),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_769),
.Y(n_969)
);

OAI221xp5_ASAP7_75t_L g970 ( 
.A1(n_890),
.A2(n_480),
.B1(n_491),
.B2(n_486),
.C(n_485),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_809),
.B(n_415),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_855),
.A2(n_495),
.B1(n_513),
.B2(n_494),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_840),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_914),
.B(n_4),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_814),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_835),
.B(n_416),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_923),
.B(n_4),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_858),
.A2(n_522),
.B1(n_523),
.B2(n_517),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_835),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_940),
.B(n_782),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_838),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_869),
.B(n_417),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_831),
.B(n_420),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_789),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_769),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_834),
.B(n_837),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_910),
.B(n_421),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_843),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_754),
.B(n_425),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_853),
.A2(n_530),
.B1(n_431),
.B2(n_435),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_L g991 ( 
.A(n_797),
.B(n_436),
.C(n_427),
.Y(n_991)
);

NAND2x1_ASAP7_75t_L g992 ( 
.A(n_849),
.B(n_469),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_910),
.B(n_437),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_908),
.B(n_438),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_850),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_851),
.A2(n_497),
.B(n_533),
.Y(n_996)
);

NAND2xp33_ASAP7_75t_L g997 ( 
.A(n_868),
.B(n_441),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_937),
.B(n_944),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_915),
.B(n_442),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_937),
.B(n_5),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_SL g1001 ( 
.A(n_867),
.B(n_450),
.C(n_445),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_944),
.B(n_452),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_854),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_919),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_835),
.B(n_531),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_924),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_861),
.B(n_456),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_755),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_925),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_933),
.B(n_458),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_761),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_947),
.B(n_461),
.Y(n_1012)
);

OAI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_882),
.A2(n_471),
.B1(n_472),
.B2(n_468),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_875),
.Y(n_1014)
);

NAND2x1_ASAP7_75t_L g1015 ( 
.A(n_765),
.B(n_335),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_948),
.B(n_474),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_781),
.A2(n_479),
.B1(n_481),
.B2(n_478),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_898),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_841),
.B(n_483),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_826),
.B(n_484),
.Y(n_1020)
);

INVxp67_ASAP7_75t_SL g1021 ( 
.A(n_763),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_763),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_851),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_796),
.B(n_493),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_865),
.A2(n_8),
.B(n_5),
.C(n_7),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_931),
.B(n_9),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_868),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_798),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_756),
.A2(n_358),
.B(n_525),
.C(n_335),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_SL g1030 ( 
.A(n_889),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_758),
.B(n_499),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_800),
.B(n_505),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_935),
.B(n_509),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_805),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_765),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_803),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_783),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_932),
.B(n_511),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_757),
.B(n_514),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_781),
.A2(n_518),
.B1(n_526),
.B2(n_516),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_770),
.B(n_9),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_SL g1042 ( 
.A(n_939),
.B(n_527),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_832),
.B(n_528),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_901),
.B(n_853),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_832),
.B(n_10),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_799),
.B(n_11),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_801),
.A2(n_358),
.B(n_335),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_781),
.A2(n_358),
.B1(n_525),
.B2(n_335),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_888),
.B(n_358),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_772),
.B(n_11),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_772),
.B(n_12),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_939),
.B(n_525),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_784),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_762),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_773),
.Y(n_1055)
);

AO22x1_ASAP7_75t_L g1056 ( 
.A1(n_785),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_825),
.B(n_14),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_857),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_928),
.B(n_15),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_772),
.B(n_16),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_794),
.B(n_16),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_794),
.B(n_17),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_868),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_772),
.B(n_776),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_859),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_776),
.B(n_17),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_864),
.B(n_860),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_819),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_781),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_L g1070 ( 
.A(n_912),
.B(n_19),
.C(n_21),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_901),
.B(n_23),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_776),
.B(n_24),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_815),
.B(n_24),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_792),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_836),
.B(n_25),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_848),
.B(n_26),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_815),
.B(n_28),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_815),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_815),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_839),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_877),
.B(n_35),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_819),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_827),
.B(n_36),
.Y(n_1083)
);

NAND3xp33_ASAP7_75t_L g1084 ( 
.A(n_913),
.B(n_38),
.C(n_39),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_759),
.B(n_40),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_911),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_L g1087 ( 
.A(n_866),
.B(n_117),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_808),
.B(n_40),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_866),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_774),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_836),
.A2(n_45),
.B1(n_42),
.B2(n_43),
.Y(n_1091)
);

AND2x6_ASAP7_75t_SL g1092 ( 
.A(n_904),
.B(n_48),
.Y(n_1092)
);

AND3x1_ASAP7_75t_L g1093 ( 
.A(n_906),
.B(n_48),
.C(n_49),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_795),
.B(n_49),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_866),
.A2(n_53),
.B1(n_50),
.B2(n_51),
.Y(n_1095)
);

NAND3xp33_ASAP7_75t_SL g1096 ( 
.A(n_830),
.B(n_50),
.C(n_53),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_848),
.B(n_54),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_888),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_920),
.B(n_54),
.Y(n_1099)
);

AND2x2_ASAP7_75t_SL g1100 ( 
.A(n_903),
.B(n_55),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_927),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_866),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_844),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_917),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_823),
.B(n_61),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_945),
.B(n_61),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_946),
.B(n_62),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_823),
.B(n_63),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_901),
.B(n_63),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_813),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_870),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_SL g1112 ( 
.A(n_883),
.B(n_119),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_778),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_847),
.B(n_64),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_885),
.B(n_66),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_818),
.B(n_67),
.Y(n_1116)
);

NOR2xp67_ASAP7_75t_L g1117 ( 
.A(n_893),
.B(n_68),
.Y(n_1117)
);

INVx8_ASAP7_75t_L g1118 ( 
.A(n_897),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_804),
.A2(n_71),
.B1(n_68),
.B2(n_70),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_911),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_956),
.B(n_881),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_954),
.Y(n_1122)
);

INVx3_ASAP7_75t_SL g1123 ( 
.A(n_958),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_960),
.B(n_807),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_963),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_R g1126 ( 
.A(n_1011),
.B(n_921),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_1110),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_975),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_981),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_965),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_979),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1023),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1030),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_1030),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_984),
.B(n_907),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_988),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_969),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_995),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1003),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1018),
.B(n_821),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_985),
.B(n_1044),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1067),
.B(n_900),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1027),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_958),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_986),
.B(n_918),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_958),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1004),
.B(n_922),
.Y(n_1147)
);

INVxp67_ASAP7_75t_SL g1148 ( 
.A(n_1082),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1027),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1057),
.A2(n_1025),
.B(n_1046),
.C(n_1080),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1006),
.B(n_941),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1009),
.B(n_816),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1058),
.Y(n_1153)
);

NOR3xp33_ASAP7_75t_SL g1154 ( 
.A(n_998),
.B(n_934),
.C(n_892),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1118),
.B(n_824),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1065),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_SL g1157 ( 
.A1(n_1100),
.A2(n_896),
.B1(n_905),
.B2(n_899),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_959),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_973),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1111),
.B(n_874),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_1118),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_SL g1162 ( 
.A(n_1074),
.B(n_891),
.C(n_895),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_SL g1163 ( 
.A(n_1074),
.B(n_777),
.C(n_894),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_SL g1164 ( 
.A(n_980),
.B(n_878),
.C(n_862),
.Y(n_1164)
);

AO22x1_ASAP7_75t_L g1165 ( 
.A1(n_1000),
.A2(n_897),
.B1(n_863),
.B2(n_845),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1021),
.B(n_906),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1028),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1000),
.B(n_957),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1044),
.B(n_900),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1068),
.B(n_886),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1036),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_SL g1172 ( 
.A(n_1061),
.B(n_791),
.C(n_780),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_SL g1173 ( 
.A(n_1034),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1022),
.B(n_902),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1090),
.B(n_961),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1037),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1053),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_1118),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_959),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_979),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1071),
.Y(n_1181)
);

INVxp67_ASAP7_75t_L g1182 ( 
.A(n_974),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_SL g1183 ( 
.A(n_1062),
.B(n_842),
.C(n_811),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1027),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1008),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1116),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1092),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1098),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1014),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1013),
.B(n_902),
.Y(n_1190)
);

NOR3xp33_ASAP7_75t_SL g1191 ( 
.A(n_1059),
.B(n_970),
.C(n_987),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_972),
.B(n_788),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_1071),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1075),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_978),
.B(n_788),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_953),
.Y(n_1196)
);

AND3x1_ASAP7_75t_SL g1197 ( 
.A(n_955),
.B(n_817),
.C(n_829),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1115),
.B(n_902),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_R g1199 ( 
.A(n_952),
.B(n_852),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_R g1200 ( 
.A(n_966),
.B(n_852),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1108),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1109),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1109),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1045),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1043),
.B(n_810),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1092),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1035),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1091),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1103),
.B(n_884),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_962),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_1063),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_977),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_991),
.A2(n_897),
.B1(n_788),
.B2(n_779),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1049),
.Y(n_1214)
);

AO22x1_ASAP7_75t_L g1215 ( 
.A1(n_1066),
.A2(n_897),
.B1(n_788),
.B2(n_812),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1001),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1041),
.B(n_1026),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_SL g1218 ( 
.A(n_1042),
.B(n_786),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_996),
.B(n_822),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1083),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1035),
.B(n_822),
.Y(n_1221)
);

BUFx8_ASAP7_75t_L g1222 ( 
.A(n_1056),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_967),
.Y(n_1223)
);

AOI221xp5_ASAP7_75t_L g1224 ( 
.A1(n_1076),
.A2(n_871),
.B1(n_872),
.B2(n_873),
.C(n_828),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1049),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1055),
.B(n_786),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_996),
.B(n_982),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_968),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_993),
.B(n_760),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1105),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1002),
.B(n_764),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1097),
.B(n_766),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_R g1233 ( 
.A(n_1066),
.B(n_768),
.Y(n_1233)
);

INVx6_ASAP7_75t_L g1234 ( 
.A(n_1117),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_971),
.A2(n_771),
.B1(n_790),
.B2(n_787),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1101),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1055),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1064),
.B(n_768),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1054),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_983),
.B(n_802),
.Y(n_1240)
);

NOR3xp33_ASAP7_75t_SL g1241 ( 
.A(n_1096),
.B(n_793),
.C(n_775),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1119),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1093),
.Y(n_1243)
);

NOR3xp33_ASAP7_75t_SL g1244 ( 
.A(n_1031),
.B(n_1033),
.C(n_951),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_992),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1208),
.B(n_1019),
.Y(n_1246)
);

NOR2xp67_ASAP7_75t_L g1247 ( 
.A(n_1127),
.B(n_1069),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1161),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1150),
.A2(n_1029),
.A3(n_1047),
.B(n_1113),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1162),
.A2(n_1163),
.B(n_1220),
.C(n_1243),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1236),
.B(n_1242),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1145),
.B(n_990),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_SL g1253 ( 
.A1(n_1193),
.A2(n_1051),
.B(n_1050),
.Y(n_1253)
);

AOI21xp33_ASAP7_75t_L g1254 ( 
.A1(n_1230),
.A2(n_1088),
.B(n_1227),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1219),
.A2(n_1085),
.A3(n_1107),
.B(n_1099),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1193),
.B(n_1199),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1201),
.A2(n_1077),
.A3(n_1073),
.B(n_1094),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1128),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1124),
.A2(n_1087),
.B(n_1224),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1147),
.A2(n_1114),
.B(n_1112),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1131),
.A2(n_1120),
.B(n_1086),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1131),
.A2(n_1015),
.B(n_1052),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1133),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1129),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1161),
.Y(n_1265)
);

AOI21xp33_ASAP7_75t_L g1266 ( 
.A1(n_1142),
.A2(n_1072),
.B(n_1060),
.Y(n_1266)
);

NAND3xp33_ASAP7_75t_L g1267 ( 
.A(n_1183),
.B(n_1048),
.C(n_1104),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1134),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1191),
.B(n_1038),
.Y(n_1269)
);

AO22x2_ASAP7_75t_L g1270 ( 
.A1(n_1121),
.A2(n_1190),
.B1(n_1167),
.B2(n_1070),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1130),
.Y(n_1271)
);

BUFx4_ASAP7_75t_SL g1272 ( 
.A(n_1155),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1161),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1122),
.B(n_989),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1204),
.A2(n_1084),
.B(n_1070),
.C(n_1106),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1136),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1135),
.B(n_950),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1132),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1138),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1167),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1214),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1151),
.A2(n_1112),
.B(n_1081),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1241),
.A2(n_1084),
.B(n_1079),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1168),
.B(n_1093),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1235),
.A2(n_999),
.B(n_994),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1139),
.B(n_1010),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1153),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1160),
.A2(n_1016),
.B(n_1012),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1152),
.A2(n_1020),
.B(n_1024),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1217),
.B(n_964),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1126),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1156),
.B(n_1171),
.Y(n_1292)
);

OAI22x1_ASAP7_75t_L g1293 ( 
.A1(n_1187),
.A2(n_1078),
.B1(n_1039),
.B2(n_1089),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1211),
.A2(n_949),
.A3(n_942),
.B(n_1032),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1181),
.A2(n_1102),
.B1(n_1095),
.B2(n_1040),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1137),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1146),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1210),
.A2(n_936),
.A3(n_938),
.B(n_916),
.Y(n_1298)
);

AO22x1_ASAP7_75t_L g1299 ( 
.A1(n_1222),
.A2(n_1042),
.B1(n_75),
.B2(n_70),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1176),
.Y(n_1300)
);

NOR3xp33_ASAP7_75t_L g1301 ( 
.A(n_1157),
.B(n_1007),
.C(n_1005),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1177),
.B(n_1017),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1194),
.B(n_802),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1202),
.A2(n_936),
.B1(n_938),
.B2(n_916),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1125),
.B(n_926),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1205),
.B(n_926),
.Y(n_1306)
);

OA22x2_ASAP7_75t_L g1307 ( 
.A1(n_1206),
.A2(n_976),
.B1(n_79),
.B2(n_72),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1164),
.A2(n_997),
.B(n_938),
.C(n_943),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1159),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1240),
.A2(n_943),
.B(n_936),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1180),
.A2(n_943),
.B(n_123),
.Y(n_1311)
);

AO32x2_ASAP7_75t_L g1312 ( 
.A1(n_1212),
.A2(n_72),
.A3(n_75),
.B1(n_80),
.B2(n_81),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1189),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1178),
.B(n_81),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1166),
.B(n_82),
.Y(n_1315)
);

AOI21xp33_ASAP7_75t_L g1316 ( 
.A1(n_1229),
.A2(n_82),
.B(n_83),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1192),
.A2(n_83),
.B(n_84),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1198),
.B(n_84),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1195),
.A2(n_128),
.B(n_122),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1198),
.B(n_85),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1213),
.A2(n_85),
.B(n_87),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1203),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1280),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1298),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1281),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1298),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1251),
.B(n_1278),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1258),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1296),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1264),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1298),
.Y(n_1331)
);

INVxp33_ASAP7_75t_L g1332 ( 
.A(n_1297),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1268),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1281),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1279),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1272),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1284),
.A2(n_1222),
.B1(n_1200),
.B2(n_1158),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1277),
.B(n_1179),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1259),
.A2(n_1182),
.B1(n_1140),
.B2(n_1234),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1314),
.B(n_1178),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1276),
.B(n_1174),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1313),
.Y(n_1342)
);

CKINVDCx6p67_ASAP7_75t_R g1343 ( 
.A(n_1263),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1311),
.A2(n_1239),
.B(n_1210),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1291),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1314),
.Y(n_1346)
);

AO21x2_ASAP7_75t_L g1347 ( 
.A1(n_1254),
.A2(n_1321),
.B(n_1260),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1287),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1309),
.Y(n_1349)
);

NAND2xp33_ASAP7_75t_L g1350 ( 
.A(n_1270),
.B(n_1143),
.Y(n_1350)
);

AOI21xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1299),
.A2(n_1216),
.B(n_1186),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1261),
.A2(n_1207),
.B(n_1209),
.Y(n_1352)
);

NAND3xp33_ASAP7_75t_L g1353 ( 
.A(n_1250),
.B(n_1172),
.C(n_1244),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1246),
.B(n_1215),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1269),
.A2(n_1252),
.B1(n_1267),
.B2(n_1247),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1310),
.A2(n_1207),
.B(n_1196),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_L g1357 ( 
.A(n_1248),
.B(n_1185),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1294),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1315),
.A2(n_1234),
.B1(n_1155),
.B2(n_1148),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1290),
.A2(n_1231),
.B1(n_1169),
.B2(n_1170),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1275),
.A2(n_1282),
.B(n_1317),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1271),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1253),
.A2(n_1228),
.B(n_1223),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1355),
.A2(n_1270),
.B1(n_1293),
.B2(n_1307),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1328),
.Y(n_1365)
);

NAND2xp33_ASAP7_75t_SL g1366 ( 
.A(n_1333),
.B(n_1233),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1340),
.A2(n_1322),
.B1(n_1295),
.B2(n_1320),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1330),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1327),
.B(n_1300),
.Y(n_1369)
);

OR2x6_ASAP7_75t_SL g1370 ( 
.A(n_1353),
.B(n_1197),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1358),
.A2(n_1340),
.B(n_1326),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1358),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1335),
.Y(n_1373)
);

CKINVDCx6p67_ASAP7_75t_R g1374 ( 
.A(n_1343),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1349),
.Y(n_1375)
);

OR2x6_ASAP7_75t_L g1376 ( 
.A(n_1340),
.B(n_1256),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1348),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1340),
.A2(n_1316),
.B1(n_1288),
.B2(n_1301),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1339),
.A2(n_1302),
.B1(n_1289),
.B2(n_1283),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1325),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1354),
.A2(n_1283),
.B1(n_1266),
.B2(n_1318),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1362),
.Y(n_1382)
);

BUFx12f_ASAP7_75t_L g1383 ( 
.A(n_1345),
.Y(n_1383)
);

AO31x2_ASAP7_75t_L g1384 ( 
.A1(n_1324),
.A2(n_1285),
.A3(n_1308),
.B(n_1304),
.Y(n_1384)
);

NAND2xp33_ASAP7_75t_R g1385 ( 
.A(n_1361),
.B(n_1265),
.Y(n_1385)
);

AO31x2_ASAP7_75t_L g1386 ( 
.A1(n_1324),
.A2(n_1319),
.A3(n_1292),
.B(n_1286),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1337),
.A2(n_1274),
.B1(n_1144),
.B2(n_1306),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1357),
.B(n_1265),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1323),
.B(n_1273),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1341),
.B(n_1312),
.Y(n_1390)
);

AO31x2_ASAP7_75t_L g1391 ( 
.A1(n_1326),
.A2(n_1305),
.A3(n_1255),
.B(n_1257),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1346),
.A2(n_1169),
.B1(n_1237),
.B2(n_1245),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1349),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1374),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1383),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1382),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1375),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1364),
.A2(n_1359),
.B1(n_1360),
.B2(n_1350),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1389),
.B(n_1329),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1376),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1376),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1376),
.A2(n_1350),
.B1(n_1325),
.B2(n_1334),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1364),
.A2(n_1332),
.B1(n_1342),
.B2(n_1327),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1365),
.B(n_1342),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1388),
.A2(n_1334),
.B1(n_1336),
.B2(n_1333),
.Y(n_1405)
);

NOR2x1_ASAP7_75t_SL g1406 ( 
.A(n_1380),
.B(n_1248),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1387),
.A2(n_1332),
.B1(n_1323),
.B2(n_1341),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1387),
.A2(n_1273),
.B1(n_1343),
.B2(n_1123),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1378),
.A2(n_1351),
.B1(n_1225),
.B2(n_1331),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1393),
.Y(n_1410)
);

OR2x6_ASAP7_75t_L g1411 ( 
.A(n_1371),
.B(n_1331),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1378),
.A2(n_1347),
.B(n_1363),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1367),
.A2(n_1347),
.B1(n_1361),
.B2(n_1338),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1366),
.A2(n_1165),
.B1(n_1141),
.B2(n_1232),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1388),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1379),
.A2(n_1381),
.B1(n_1368),
.B2(n_1377),
.Y(n_1416)
);

AND2x4_ASAP7_75t_SL g1417 ( 
.A(n_1380),
.B(n_1141),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1397),
.B(n_1372),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1404),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1411),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1397),
.B(n_1410),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1410),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1417),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1396),
.B(n_1372),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1415),
.B(n_1391),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1411),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1411),
.B(n_1391),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1401),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1399),
.B(n_1391),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1401),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1400),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1401),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1400),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1413),
.B(n_1391),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1413),
.B(n_1390),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1400),
.Y(n_1436)
);

AOI221x1_ASAP7_75t_L g1437 ( 
.A1(n_1426),
.A2(n_1408),
.B1(n_1409),
.B2(n_1412),
.C(n_1407),
.Y(n_1437)
);

AOI33xp33_ASAP7_75t_L g1438 ( 
.A1(n_1435),
.A2(n_1403),
.A3(n_1405),
.B1(n_1398),
.B2(n_1416),
.B3(n_1394),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1423),
.Y(n_1439)
);

OAI33xp33_ASAP7_75t_L g1440 ( 
.A1(n_1419),
.A2(n_1373),
.A3(n_1369),
.B1(n_1395),
.B2(n_1370),
.B3(n_1403),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1423),
.A2(n_1398),
.B1(n_1402),
.B2(n_1417),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1435),
.A2(n_1416),
.B1(n_1379),
.B2(n_1381),
.C(n_1392),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1429),
.B(n_1384),
.Y(n_1443)
);

AOI322xp5_ASAP7_75t_L g1444 ( 
.A1(n_1434),
.A2(n_1392),
.A3(n_1395),
.B1(n_1414),
.B2(n_1345),
.C1(n_1312),
.C2(n_1406),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1423),
.A2(n_1361),
.B1(n_1347),
.B2(n_1363),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1424),
.B(n_1386),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1431),
.A2(n_1356),
.B(n_1344),
.Y(n_1447)
);

AOI211x1_ASAP7_75t_L g1448 ( 
.A1(n_1433),
.A2(n_1426),
.B(n_1427),
.C(n_1434),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1427),
.B(n_1384),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1443),
.B(n_1420),
.Y(n_1450)
);

NAND2x1p5_ASAP7_75t_SL g1451 ( 
.A(n_1439),
.B(n_1436),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1439),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1438),
.B(n_1443),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1446),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1449),
.B(n_1418),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1445),
.B(n_1418),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1438),
.B(n_1425),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1448),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1441),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1444),
.B(n_1421),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1442),
.B(n_1425),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1447),
.Y(n_1462)
);

OR2x2_ASAP7_75t_SL g1463 ( 
.A(n_1440),
.B(n_1436),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1437),
.Y(n_1464)
);

INVxp33_ASAP7_75t_L g1465 ( 
.A(n_1464),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1460),
.B(n_1433),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1452),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1460),
.B(n_1422),
.Y(n_1468)
);

NAND2x1_ASAP7_75t_SL g1469 ( 
.A(n_1458),
.B(n_1431),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1451),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1470),
.B(n_1459),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1467),
.B(n_1431),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1467),
.B(n_1450),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1472),
.A2(n_1470),
.B1(n_1453),
.B2(n_1457),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1471),
.A2(n_1465),
.B1(n_1461),
.B2(n_1466),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1475),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1474),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1475),
.B(n_1465),
.C(n_1471),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1476),
.B(n_1471),
.Y(n_1479)
);

AOI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1476),
.A2(n_1468),
.B1(n_1462),
.B2(n_1473),
.C(n_1472),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1478),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1477),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1481),
.B(n_1454),
.Y(n_1483)
);

NAND4xp25_ASAP7_75t_L g1484 ( 
.A(n_1479),
.B(n_1170),
.C(n_1456),
.D(n_1462),
.Y(n_1484)
);

NOR3xp33_ASAP7_75t_L g1485 ( 
.A(n_1480),
.B(n_1188),
.C(n_1175),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1482),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1482),
.B(n_1463),
.Y(n_1487)
);

AOI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1486),
.A2(n_1462),
.B1(n_1173),
.B2(n_1451),
.C(n_1456),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1487),
.A2(n_1455),
.B1(n_1154),
.B2(n_1385),
.Y(n_1489)
);

OAI221xp5_ASAP7_75t_L g1490 ( 
.A1(n_1485),
.A2(n_1469),
.B1(n_1218),
.B2(n_1385),
.C(n_1428),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1483),
.B(n_1303),
.C(n_1226),
.Y(n_1491)
);

OAI321xp33_ASAP7_75t_L g1492 ( 
.A1(n_1484),
.A2(n_1432),
.A3(n_1430),
.B1(n_1312),
.B2(n_92),
.C(n_93),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1486),
.A2(n_1221),
.B1(n_1422),
.B2(n_1226),
.C(n_1238),
.Y(n_1493)
);

AOI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1492),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.C(n_100),
.Y(n_1494)
);

AOI21xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1489),
.A2(n_101),
.B(n_103),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1488),
.A2(n_1352),
.B1(n_1262),
.B2(n_1184),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1493),
.A2(n_1143),
.B1(n_1149),
.B2(n_1184),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1491),
.B(n_105),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1490),
.B(n_106),
.Y(n_1499)
);

INVxp67_ASAP7_75t_SL g1500 ( 
.A(n_1499),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1498),
.B(n_108),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1496),
.B(n_112),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1497),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_1495),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1494),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1501),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1505),
.B(n_130),
.Y(n_1507)
);

AOI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1504),
.A2(n_1257),
.B1(n_1249),
.B2(n_137),
.C(n_139),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1506),
.A2(n_1500),
.B1(n_1503),
.B2(n_1502),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1507),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1508),
.B(n_140),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1509),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1512),
.A2(n_1510),
.B1(n_1511),
.B2(n_1249),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1513),
.Y(n_1514)
);

AOI21xp33_ASAP7_75t_L g1515 ( 
.A1(n_1514),
.A2(n_146),
.B(n_147),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1515),
.Y(n_1516)
);

AOI322xp5_ASAP7_75t_L g1517 ( 
.A1(n_1516),
.A2(n_1386),
.A3(n_1384),
.B1(n_162),
.B2(n_165),
.C1(n_167),
.C2(n_169),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_SL g1518 ( 
.A1(n_1516),
.A2(n_171),
.B1(n_172),
.B2(n_174),
.Y(n_1518)
);

AOI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1518),
.A2(n_180),
.B1(n_182),
.B2(n_184),
.C(n_185),
.Y(n_1519)
);

AOI211xp5_ASAP7_75t_L g1520 ( 
.A1(n_1519),
.A2(n_1517),
.B(n_186),
.C(n_187),
.Y(n_1520)
);


endmodule