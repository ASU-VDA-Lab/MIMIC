module fake_aes_9280_n_38 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
OAI22xp5_ASAP7_75t_SL g15 ( .A1(n_11), .A2(n_1), .B1(n_10), .B2(n_4), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_5), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_14), .B(n_2), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_1), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_16), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_0), .Y(n_23) );
NAND2xp5_ASAP7_75t_SL g24 ( .A(n_16), .B(n_0), .Y(n_24) );
INVx1_ASAP7_75t_SL g25 ( .A(n_23), .Y(n_25) );
OR2x6_ASAP7_75t_L g26 ( .A(n_24), .B(n_15), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_27), .B(n_25), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_28), .B(n_26), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NAND2xp33_ASAP7_75t_R g31 ( .A(n_29), .B(n_2), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_22), .Y(n_32) );
OAI211xp5_ASAP7_75t_SL g33 ( .A1(n_32), .A2(n_17), .B(n_18), .C(n_16), .Y(n_33) );
NOR2xp67_ASAP7_75t_L g34 ( .A(n_31), .B(n_29), .Y(n_34) );
OAI22xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_19), .B1(n_20), .B2(n_3), .Y(n_35) );
OAI22x1_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_3), .B1(n_19), .B2(n_7), .Y(n_36) );
OAI22xp5_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_20), .B1(n_6), .B2(n_13), .Y(n_37) );
AOI22x1_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_20), .B1(n_36), .B2(n_16), .Y(n_38) );
endmodule