module real_aes_909_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g242 ( .A(n_0), .B(n_163), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_1), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_2), .B(n_147), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_3), .B(n_165), .Y(n_493) );
INVx1_ASAP7_75t_L g154 ( .A(n_4), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_5), .B(n_147), .Y(n_146) );
NAND2xp33_ASAP7_75t_SL g233 ( .A(n_6), .B(n_153), .Y(n_233) );
INVx1_ASAP7_75t_L g214 ( .A(n_7), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_8), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_9), .Y(n_109) );
AND2x2_ASAP7_75t_L g141 ( .A(n_10), .B(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g495 ( .A(n_11), .B(n_204), .Y(n_495) );
AND2x2_ASAP7_75t_L g503 ( .A(n_12), .B(n_230), .Y(n_503) );
INVx2_ASAP7_75t_L g143 ( .A(n_13), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_14), .B(n_165), .Y(n_512) );
XNOR2xp5_ASAP7_75t_L g773 ( .A(n_15), .B(n_774), .Y(n_773) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_16), .B(n_108), .C(n_110), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_16), .Y(n_126) );
AOI221x1_ASAP7_75t_L g227 ( .A1(n_17), .A2(n_156), .B1(n_228), .B2(n_230), .C(n_232), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_18), .B(n_147), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_19), .B(n_147), .Y(n_526) );
INVx1_ASAP7_75t_L g113 ( .A(n_20), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_21), .A2(n_89), .B1(n_147), .B2(n_215), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_22), .A2(n_156), .B(n_161), .Y(n_155) );
AOI221xp5_ASAP7_75t_SL g191 ( .A1(n_23), .A2(n_37), .B1(n_147), .B2(n_156), .C(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_24), .B(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g144 ( .A(n_25), .B(n_88), .Y(n_144) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_25), .A2(n_88), .B(n_143), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_26), .B(n_165), .Y(n_203) );
INVxp67_ASAP7_75t_L g226 ( .A(n_27), .Y(n_226) );
AND2x2_ASAP7_75t_L g187 ( .A(n_28), .B(n_177), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_29), .A2(n_156), .B(n_241), .Y(n_240) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_30), .A2(n_230), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_31), .B(n_165), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_32), .A2(n_156), .B(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_33), .B(n_165), .Y(n_521) );
AND2x2_ASAP7_75t_L g153 ( .A(n_34), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g157 ( .A(n_34), .B(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g222 ( .A(n_34), .Y(n_222) );
INVxp67_ASAP7_75t_L g110 ( .A(n_35), .Y(n_110) );
OR2x6_ASAP7_75t_L g128 ( .A(n_35), .B(n_129), .Y(n_128) );
INVxp33_ASAP7_75t_L g799 ( .A(n_36), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_38), .B(n_147), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_39), .A2(n_81), .B1(n_156), .B2(n_220), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_40), .B(n_165), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_41), .B(n_147), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_42), .A2(n_73), .B1(n_795), .B2(n_796), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_42), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_43), .B(n_163), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_44), .A2(n_156), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g245 ( .A(n_45), .B(n_177), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_46), .B(n_163), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_47), .B(n_177), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_48), .B(n_147), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g792 ( .A1(n_49), .A2(n_793), .B1(n_794), .B2(n_797), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_49), .Y(n_797) );
INVx1_ASAP7_75t_L g150 ( .A(n_50), .Y(n_150) );
INVx1_ASAP7_75t_L g160 ( .A(n_50), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_51), .B(n_165), .Y(n_501) );
AND2x2_ASAP7_75t_L g537 ( .A(n_52), .B(n_177), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_53), .B(n_147), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_54), .B(n_163), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_55), .B(n_163), .Y(n_520) );
AND2x2_ASAP7_75t_L g178 ( .A(n_56), .B(n_177), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_57), .B(n_147), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_58), .B(n_165), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_59), .B(n_147), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_60), .A2(n_156), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_61), .B(n_163), .Y(n_174) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_62), .B(n_142), .Y(n_206) );
AND2x2_ASAP7_75t_L g532 ( .A(n_63), .B(n_142), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_64), .A2(n_156), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_65), .B(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_SL g258 ( .A(n_66), .B(n_204), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_67), .B(n_163), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_68), .B(n_163), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_69), .A2(n_92), .B1(n_156), .B2(n_220), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_70), .B(n_165), .Y(n_529) );
INVx1_ASAP7_75t_L g152 ( .A(n_71), .Y(n_152) );
INVx1_ASAP7_75t_L g158 ( .A(n_71), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_72), .B(n_163), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_73), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_74), .A2(n_156), .B(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_75), .A2(n_156), .B(n_483), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_76), .A2(n_156), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g523 ( .A(n_77), .B(n_142), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_78), .B(n_177), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_79), .B(n_147), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_80), .A2(n_83), .B1(n_147), .B2(n_215), .Y(n_256) );
INVx1_ASAP7_75t_L g112 ( .A(n_82), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_84), .B(n_163), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_85), .B(n_163), .Y(n_194) );
AND2x2_ASAP7_75t_L g486 ( .A(n_86), .B(n_204), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_87), .A2(n_156), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_90), .B(n_165), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_91), .A2(n_156), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_93), .B(n_165), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_94), .A2(n_102), .B1(n_775), .B2(n_776), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_94), .Y(n_775) );
INVxp67_ASAP7_75t_L g229 ( .A(n_95), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_96), .B(n_147), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_97), .B(n_165), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_98), .A2(n_156), .B(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g531 ( .A(n_99), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_100), .A2(n_773), .B1(n_778), .B2(n_781), .Y(n_777) );
BUFx2_ASAP7_75t_L g118 ( .A(n_101), .Y(n_118) );
BUFx2_ASAP7_75t_SL g787 ( .A(n_101), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_102), .Y(n_776) );
AOI21xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_114), .B(n_798), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx3_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g802 ( .A(n_106), .Y(n_802) );
NAND2xp5_ASAP7_75t_SL g106 ( .A(n_107), .B(n_111), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_112), .B(n_113), .Y(n_129) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_131), .B(n_785), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_119), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI21xp33_ASAP7_75t_SL g788 ( .A1(n_120), .A2(n_789), .B(n_790), .Y(n_788) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_130), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g789 ( .A(n_125), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x6_ASAP7_75t_SL g471 ( .A(n_126), .B(n_128), .Y(n_471) );
OR2x6_ASAP7_75t_SL g772 ( .A(n_126), .B(n_127), .Y(n_772) );
OR2x2_ASAP7_75t_L g784 ( .A(n_126), .B(n_128), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
OAI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_773), .B(n_777), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_468), .B1(n_472), .B2(n_772), .Y(n_133) );
OAI22x1_ASAP7_75t_L g790 ( .A1(n_134), .A2(n_135), .B1(n_791), .B2(n_792), .Y(n_790) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_135), .A2(n_468), .B1(n_473), .B2(n_779), .Y(n_778) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_379), .Y(n_135) );
NOR3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_301), .C(n_351), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_268), .Y(n_137) );
AOI221xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_188), .B1(n_207), .B2(n_250), .C(n_260), .Y(n_138) );
INVx1_ASAP7_75t_SL g350 ( .A(n_139), .Y(n_350) );
AND2x4_ASAP7_75t_SL g139 ( .A(n_140), .B(n_168), .Y(n_139) );
INVx2_ASAP7_75t_L g272 ( .A(n_140), .Y(n_272) );
OR2x2_ASAP7_75t_L g294 ( .A(n_140), .B(n_285), .Y(n_294) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_140), .Y(n_309) );
INVx5_ASAP7_75t_L g316 ( .A(n_140), .Y(n_316) );
AND2x4_ASAP7_75t_L g322 ( .A(n_140), .B(n_180), .Y(n_322) );
AND2x2_ASAP7_75t_SL g325 ( .A(n_140), .B(n_252), .Y(n_325) );
OR2x2_ASAP7_75t_L g334 ( .A(n_140), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g341 ( .A(n_140), .B(n_169), .Y(n_341) );
AND2x2_ASAP7_75t_L g442 ( .A(n_140), .B(n_179), .Y(n_442) );
OR2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x4_ASAP7_75t_L g167 ( .A(n_143), .B(n_144), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_155), .B(n_167), .Y(n_145) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_153), .Y(n_147) );
INVx1_ASAP7_75t_L g234 ( .A(n_148), .Y(n_234) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
AND2x6_ASAP7_75t_L g163 ( .A(n_149), .B(n_158), .Y(n_163) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g165 ( .A(n_151), .B(n_160), .Y(n_165) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx5_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
AND2x2_ASAP7_75t_L g159 ( .A(n_154), .B(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_154), .Y(n_218) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
BUFx3_ASAP7_75t_L g219 ( .A(n_157), .Y(n_219) );
INVx2_ASAP7_75t_L g224 ( .A(n_158), .Y(n_224) );
AND2x4_ASAP7_75t_L g220 ( .A(n_159), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g217 ( .A(n_160), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B(n_166), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_163), .B(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_166), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_166), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_166), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_166), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_166), .A2(n_242), .B(n_243), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_166), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_166), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_166), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_166), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_166), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_166), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_166), .A2(n_542), .B(n_543), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_167), .B(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_167), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_167), .B(n_229), .Y(n_228) );
NOR3xp33_ASAP7_75t_L g232 ( .A(n_167), .B(n_233), .C(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_167), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_167), .A2(n_539), .B(n_540), .Y(n_538) );
INVx3_ASAP7_75t_SL g293 ( .A(n_168), .Y(n_293) );
AND2x2_ASAP7_75t_L g337 ( .A(n_168), .B(n_252), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_168), .A2(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g378 ( .A(n_168), .B(n_316), .Y(n_378) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_179), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_169), .B(n_180), .Y(n_259) );
OR2x2_ASAP7_75t_L g263 ( .A(n_169), .B(n_180), .Y(n_263) );
INVx1_ASAP7_75t_L g271 ( .A(n_169), .Y(n_271) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_169), .Y(n_283) );
INVx2_ASAP7_75t_L g291 ( .A(n_169), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_169), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g400 ( .A(n_169), .B(n_285), .Y(n_400) );
AND2x2_ASAP7_75t_L g415 ( .A(n_169), .B(n_252), .Y(n_415) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_176), .B(n_178), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_175), .Y(n_170) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_176), .A2(n_181), .B(n_187), .Y(n_180) );
AO21x2_ASAP7_75t_L g335 ( .A1(n_176), .A2(n_181), .B(n_187), .Y(n_335) );
AOI21x1_ASAP7_75t_L g488 ( .A1(n_176), .A2(n_489), .B(n_495), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_177), .A2(n_191), .B(n_195), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_177), .A2(n_481), .B(n_482), .Y(n_480) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_177), .A2(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g284 ( .A(n_180), .B(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_180), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_186), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_188), .B(n_408), .Y(n_407) );
NOR2x1p5_ASAP7_75t_L g188 ( .A(n_189), .B(n_196), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g236 ( .A(n_190), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_190), .B(n_197), .Y(n_266) );
INVx1_ASAP7_75t_L g276 ( .A(n_190), .Y(n_276) );
INVx2_ASAP7_75t_L g299 ( .A(n_190), .Y(n_299) );
INVx2_ASAP7_75t_L g305 ( .A(n_190), .Y(n_305) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_190), .Y(n_375) );
OR2x2_ASAP7_75t_L g406 ( .A(n_190), .B(n_197), .Y(n_406) );
OR2x2_ASAP7_75t_L g422 ( .A(n_196), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x4_ASAP7_75t_SL g210 ( .A(n_197), .B(n_211), .Y(n_210) );
AND2x4_ASAP7_75t_L g248 ( .A(n_197), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g286 ( .A(n_197), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g298 ( .A(n_197), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g311 ( .A(n_197), .B(n_277), .Y(n_311) );
OR2x2_ASAP7_75t_L g319 ( .A(n_197), .B(n_211), .Y(n_319) );
INVx2_ASAP7_75t_L g346 ( .A(n_197), .Y(n_346) );
INVx1_ASAP7_75t_L g364 ( .A(n_197), .Y(n_364) );
NOR2xp33_ASAP7_75t_R g397 ( .A(n_197), .B(n_237), .Y(n_397) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_206), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_204), .Y(n_198) );
INVx2_ASAP7_75t_SL g254 ( .A(n_204), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_204), .A2(n_526), .B(n_527), .Y(n_525) );
BUFx4f_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g231 ( .A(n_205), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_208), .B(n_246), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_208), .A2(n_289), .B1(n_292), .B2(n_295), .Y(n_288) );
OR2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_235), .Y(n_208) );
INVx1_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g303 ( .A(n_210), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g338 ( .A(n_210), .B(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g417 ( .A(n_210), .B(n_395), .Y(n_417) );
INVx3_ASAP7_75t_L g249 ( .A(n_211), .Y(n_249) );
AND2x4_ASAP7_75t_L g277 ( .A(n_211), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_211), .B(n_237), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_211), .B(n_299), .Y(n_344) );
AND2x2_ASAP7_75t_L g349 ( .A(n_211), .B(n_346), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_211), .B(n_236), .Y(n_386) );
INVx1_ASAP7_75t_L g456 ( .A(n_211), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_211), .B(n_374), .Y(n_467) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_227), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_215), .B1(n_220), .B2(n_225), .Y(n_212) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_219), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
NOR2x1p5_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx3_ASAP7_75t_L g516 ( .A(n_230), .Y(n_516) );
INVx4_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AOI21x1_ASAP7_75t_L g238 ( .A1(n_231), .A2(n_239), .B(n_245), .Y(n_238) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_231), .A2(n_497), .B(n_503), .Y(n_496) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g247 ( .A(n_237), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_237), .B(n_249), .Y(n_267) );
INVx2_ASAP7_75t_L g278 ( .A(n_237), .Y(n_278) );
AND2x2_ASAP7_75t_L g304 ( .A(n_237), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g320 ( .A(n_237), .B(n_299), .Y(n_320) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_237), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_237), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g409 ( .A(n_237), .Y(n_409) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_244), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_247), .B(n_276), .Y(n_287) );
AOI221x1_ASAP7_75t_SL g381 ( .A1(n_248), .A2(n_382), .B1(n_385), .B2(n_387), .C(n_391), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_248), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g439 ( .A(n_248), .B(n_304), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_248), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g370 ( .A(n_249), .B(n_298), .Y(n_370) );
AND2x2_ASAP7_75t_L g408 ( .A(n_249), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_259), .Y(n_251) );
AND2x2_ASAP7_75t_L g261 ( .A(n_252), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g356 ( .A(n_252), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_252), .B(n_272), .Y(n_361) );
AND2x4_ASAP7_75t_L g390 ( .A(n_252), .B(n_291), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_252), .B(n_322), .Y(n_426) );
OR2x2_ASAP7_75t_L g444 ( .A(n_252), .B(n_375), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_252), .B(n_335), .Y(n_454) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g285 ( .A(n_253), .Y(n_285) );
AOI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_258), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g310 ( .A(n_259), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_259), .A2(n_318), .B1(n_321), .B2(n_323), .Y(n_317) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx2_ASAP7_75t_L g273 ( .A(n_261), .Y(n_273) );
AND2x2_ASAP7_75t_L g412 ( .A(n_262), .B(n_272), .Y(n_412) );
AND2x2_ASAP7_75t_L g458 ( .A(n_262), .B(n_325), .Y(n_458) );
AND2x2_ASAP7_75t_L g463 ( .A(n_262), .B(n_314), .Y(n_463) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AOI32xp33_ASAP7_75t_L g432 ( .A1(n_264), .A2(n_334), .A3(n_414), .B1(n_433), .B2(n_435), .Y(n_432) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g300 ( .A(n_267), .Y(n_300) );
AOI211xp5_ASAP7_75t_SL g268 ( .A1(n_269), .A2(n_274), .B(n_279), .C(n_288), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_272), .B(n_273), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_271), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_272), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g452 ( .A(n_272), .Y(n_452) );
AND2x2_ASAP7_75t_L g362 ( .A(n_274), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_SL g274 ( .A(n_275), .B(n_277), .Y(n_274) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_275), .Y(n_462) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_276), .Y(n_331) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_276), .Y(n_431) );
INVx1_ASAP7_75t_L g328 ( .A(n_277), .Y(n_328) );
AND2x2_ASAP7_75t_L g394 ( .A(n_277), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_277), .B(n_405), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_286), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI21xp33_ASAP7_75t_L g360 ( .A1(n_281), .A2(n_361), .B(n_362), .Y(n_360) );
AND2x2_ASAP7_75t_SL g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g290 ( .A(n_285), .B(n_291), .Y(n_290) );
BUFx2_ASAP7_75t_L g314 ( .A(n_285), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_290), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g421 ( .A(n_290), .Y(n_421) );
AND2x2_ASAP7_75t_L g451 ( .A(n_290), .B(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_291), .Y(n_428) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_293), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g368 ( .A(n_294), .Y(n_368) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g327 ( .A(n_298), .B(n_328), .Y(n_327) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_299), .Y(n_395) );
AND2x2_ASAP7_75t_L g404 ( .A(n_300), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_324), .Y(n_301) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_306), .B1(n_311), .B2(n_312), .C(n_317), .Y(n_302) );
INVx1_ASAP7_75t_L g423 ( .A(n_304), .Y(n_423) );
INVxp33_ASAP7_75t_SL g455 ( .A(n_304), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_306), .A2(n_402), .B(n_410), .Y(n_401) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_310), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g323 ( .A(n_311), .Y(n_323) );
AND2x2_ASAP7_75t_L g358 ( .A(n_311), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g377 ( .A(n_311), .B(n_378), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_311), .A2(n_439), .B1(n_440), .B2(n_443), .Y(n_438) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
OR2x2_ASAP7_75t_L g333 ( .A(n_314), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_314), .B(n_322), .Y(n_372) );
AND2x4_ASAP7_75t_L g389 ( .A(n_316), .B(n_335), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_316), .B(n_390), .Y(n_436) );
AND2x2_ASAP7_75t_L g448 ( .A(n_316), .B(n_400), .Y(n_448) );
NAND2xp33_ASAP7_75t_L g433 ( .A(n_318), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_SL g376 ( .A(n_319), .Y(n_376) );
INVx1_ASAP7_75t_L g447 ( .A(n_320), .Y(n_447) );
INVx2_ASAP7_75t_SL g399 ( .A(n_322), .Y(n_399) );
AOI211xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_326), .B(n_329), .C(n_347), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI211xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B(n_336), .C(n_340), .Y(n_329) );
OR2x6_ASAP7_75t_SL g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g359 ( .A(n_331), .Y(n_359) );
INVx1_ASAP7_75t_SL g384 ( .A(n_334), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_334), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_339), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g425 ( .A1(n_343), .A2(n_426), .B1(n_427), .B2(n_429), .Y(n_425) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
OAI211xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_357), .B(n_360), .C(n_365), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_369), .B1(n_371), .B2(n_373), .C(n_377), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_376), .A2(n_458), .B1(n_459), .B2(n_463), .C1(n_464), .C2(n_466), .Y(n_457) );
INVx2_ASAP7_75t_L g392 ( .A(n_378), .Y(n_392) );
NOR3xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_418), .C(n_437), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_401), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_389), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_390), .B(n_452), .Y(n_465) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_396), .B2(n_398), .Y(n_391) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVxp33_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_399), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_407), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_407), .A2(n_411), .B1(n_413), .B2(n_416), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
CKINVDCx16_ASAP7_75t_R g416 ( .A(n_417), .Y(n_416) );
OAI211xp5_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_422), .B(n_424), .C(n_432), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_445), .C(n_457), .Y(n_437) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_449), .B(n_456), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_453), .B(n_455), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
CKINVDCx11_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
INVx5_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_676), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_601), .C(n_637), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_575), .Y(n_475) );
AOI211xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_504), .B(n_533), .C(n_558), .Y(n_476) );
AND2x2_ASAP7_75t_L g666 ( .A(n_477), .B(n_535), .Y(n_666) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_487), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_478), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g699 ( .A(n_478), .B(n_581), .Y(n_699) );
AND2x2_ASAP7_75t_L g715 ( .A(n_478), .B(n_550), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_478), .B(n_725), .Y(n_724) );
NAND2x1p5_ASAP7_75t_L g748 ( .A(n_478), .B(n_749), .Y(n_748) );
INVx4_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_SL g545 ( .A(n_479), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g570 ( .A(n_479), .Y(n_570) );
AND2x2_ASAP7_75t_L g617 ( .A(n_479), .B(n_560), .Y(n_617) );
AND2x2_ASAP7_75t_L g636 ( .A(n_479), .B(n_487), .Y(n_636) );
BUFx2_ASAP7_75t_L g641 ( .A(n_479), .Y(n_641) );
AND2x2_ASAP7_75t_L g685 ( .A(n_479), .B(n_496), .Y(n_685) );
AND2x4_ASAP7_75t_L g757 ( .A(n_479), .B(n_758), .Y(n_757) );
NOR2x1_ASAP7_75t_L g769 ( .A(n_479), .B(n_549), .Y(n_769) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_486), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_487), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g688 ( .A(n_487), .Y(n_688) );
BUFx2_ASAP7_75t_L g737 ( .A(n_487), .Y(n_737) );
INVx1_ASAP7_75t_L g759 ( .A(n_487), .Y(n_759) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_496), .Y(n_487) );
INVx3_ASAP7_75t_L g546 ( .A(n_488), .Y(n_546) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_488), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_494), .Y(n_489) );
INVx2_ASAP7_75t_L g549 ( .A(n_496), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_496), .B(n_546), .Y(n_550) );
INVx2_ASAP7_75t_L g625 ( .A(n_496), .Y(n_625) );
OR2x2_ASAP7_75t_L g632 ( .A(n_496), .B(n_581), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_502), .Y(n_497) );
AND2x2_ASAP7_75t_L g587 ( .A(n_504), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g621 ( .A(n_504), .B(n_584), .Y(n_621) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
AND2x2_ASAP7_75t_L g657 ( .A(n_505), .B(n_556), .Y(n_657) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g614 ( .A(n_506), .B(n_515), .Y(n_614) );
AND2x2_ASAP7_75t_L g733 ( .A(n_506), .B(n_524), .Y(n_733) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g555 ( .A(n_507), .Y(n_555) );
INVx1_ASAP7_75t_L g573 ( .A(n_507), .Y(n_573) );
AND2x2_ASAP7_75t_L g629 ( .A(n_507), .B(n_515), .Y(n_629) );
AND2x2_ASAP7_75t_L g634 ( .A(n_507), .B(n_536), .Y(n_634) );
OR2x2_ASAP7_75t_L g697 ( .A(n_507), .B(n_524), .Y(n_697) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_507), .Y(n_706) );
AND2x2_ASAP7_75t_L g535 ( .A(n_514), .B(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g574 ( .A(n_514), .Y(n_574) );
NOR2x1_ASAP7_75t_SL g514 ( .A(n_515), .B(n_524), .Y(n_514) );
AO21x1_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_517), .B(n_523), .Y(n_515) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_516), .A2(n_517), .B(n_523), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
AND2x2_ASAP7_75t_L g552 ( .A(n_524), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g600 ( .A(n_524), .Y(n_600) );
NAND2x1_ASAP7_75t_L g610 ( .A(n_524), .B(n_536), .Y(n_610) );
OR2x2_ASAP7_75t_L g615 ( .A(n_524), .B(n_553), .Y(n_615) );
BUFx2_ASAP7_75t_L g671 ( .A(n_524), .Y(n_671) );
AND2x2_ASAP7_75t_L g707 ( .A(n_524), .B(n_586), .Y(n_707) );
AND2x2_ASAP7_75t_L g718 ( .A(n_524), .B(n_556), .Y(n_718) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_532), .Y(n_524) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_544), .B1(n_550), .B2(n_551), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_535), .A2(n_715), .B1(n_765), .B2(n_770), .Y(n_764) );
INVx4_ASAP7_75t_L g553 ( .A(n_536), .Y(n_553) );
INVx2_ASAP7_75t_L g584 ( .A(n_536), .Y(n_584) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_536), .Y(n_655) );
OR2x2_ASAP7_75t_L g670 ( .A(n_536), .B(n_556), .Y(n_670) );
OR2x2_ASAP7_75t_SL g696 ( .A(n_536), .B(n_697), .Y(n_696) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_SL g544 ( .A(n_545), .B(n_547), .Y(n_544) );
INVx2_ASAP7_75t_SL g577 ( .A(n_545), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_545), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g645 ( .A(n_545), .B(n_593), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_545), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g567 ( .A(n_546), .Y(n_567) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_546), .Y(n_592) );
AND2x2_ASAP7_75t_L g648 ( .A(n_546), .B(n_625), .Y(n_648) );
INVx1_ASAP7_75t_L g758 ( .A(n_546), .Y(n_758) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_548), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_548), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g566 ( .A(n_549), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_550), .B(n_699), .Y(n_698) );
AOI321xp33_ASAP7_75t_L g720 ( .A1(n_551), .A2(n_622), .A3(n_690), .B1(n_721), .B2(n_722), .C(n_726), .Y(n_720) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_552), .Y(n_619) );
AND2x2_ASAP7_75t_L g644 ( .A(n_552), .B(n_573), .Y(n_644) );
AND2x2_ASAP7_75t_L g719 ( .A(n_552), .B(n_629), .Y(n_719) );
INVx1_ASAP7_75t_L g588 ( .A(n_553), .Y(n_588) );
BUFx2_ASAP7_75t_L g598 ( .A(n_553), .Y(n_598) );
NOR2xp67_ASAP7_75t_L g705 ( .A(n_553), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g643 ( .A(n_554), .Y(n_643) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
BUFx2_ASAP7_75t_L g650 ( .A(n_555), .Y(n_650) );
INVx2_ASAP7_75t_L g586 ( .A(n_556), .Y(n_586) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_556), .Y(n_609) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AOI21xp33_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_568), .B(n_571), .Y(n_558) );
NOR2xp67_ASAP7_75t_L g702 ( .A(n_559), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_566), .Y(n_560) );
INVx3_ASAP7_75t_L g593 ( .A(n_561), .Y(n_593) );
AND2x2_ASAP7_75t_L g624 ( .A(n_561), .B(n_625), .Y(n_624) );
AND2x4_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x4_ASAP7_75t_L g581 ( .A(n_562), .B(n_563), .Y(n_581) );
INVx1_ASAP7_75t_L g664 ( .A(n_566), .Y(n_664) );
INVx1_ASAP7_75t_SL g749 ( .A(n_567), .Y(n_749) );
INVxp33_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_570), .B(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g675 ( .A(n_570), .B(n_632), .Y(n_675) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND2x2_ASAP7_75t_L g679 ( .A(n_572), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_572), .B(n_694), .Y(n_693) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_573), .B(n_610), .Y(n_665) );
NOR4xp25_ASAP7_75t_L g760 ( .A(n_573), .B(n_604), .C(n_761), .D(n_762), .Y(n_760) );
OR2x2_ASAP7_75t_L g728 ( .A(n_574), .B(n_729), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_582), .B1(n_587), .B2(n_589), .C(n_594), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AND2x2_ASAP7_75t_L g603 ( .A(n_578), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g640 ( .A(n_579), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g660 ( .A(n_580), .Y(n_660) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx3_ASAP7_75t_L g683 ( .A(n_581), .Y(n_683) );
AND2x2_ASAP7_75t_L g690 ( .A(n_581), .B(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
OR2x2_ASAP7_75t_L g627 ( .A(n_584), .B(n_628), .Y(n_627) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_586), .B(n_600), .Y(n_599) );
INVxp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx2_ASAP7_75t_L g604 ( .A(n_591), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_591), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g596 ( .A(n_593), .Y(n_596) );
OAI321xp33_ASAP7_75t_L g708 ( .A1(n_593), .A2(n_701), .A3(n_709), .B1(n_714), .B2(n_716), .C(n_720), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
OR2x2_ASAP7_75t_L g663 ( .A(n_596), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g763 ( .A(n_599), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_600), .B(n_643), .Y(n_642) );
NAND2xp33_ASAP7_75t_SL g743 ( .A(n_600), .B(n_614), .Y(n_743) );
OAI211xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B(n_616), .C(n_620), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_611), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g712 ( .A(n_609), .Y(n_712) );
INVx3_ASAP7_75t_L g651 ( .A(n_610), .Y(n_651) );
OR2x2_ASAP7_75t_L g754 ( .A(n_610), .B(n_628), .Y(n_754) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_612), .A2(n_696), .B1(n_698), .B2(n_700), .Y(n_695) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_SL g694 ( .A(n_615), .Y(n_694) );
OR2x2_ASAP7_75t_L g771 ( .A(n_615), .B(n_628), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AOI21xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_622), .B(n_626), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_624), .B(n_641), .Y(n_740) );
AND2x2_ASAP7_75t_L g746 ( .A(n_624), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g691 ( .A(n_625), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_630), .B1(n_633), .B2(n_635), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_628), .A2(n_671), .B(n_673), .C(n_675), .Y(n_672) );
INVx2_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_631), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_631), .B(n_723), .Y(n_745) );
INVx2_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g717 ( .A(n_634), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_636), .A2(n_668), .B(n_671), .C(n_672), .Y(n_667) );
NAND3xp33_ASAP7_75t_SL g637 ( .A(n_638), .B(n_652), .C(n_667), .Y(n_637) );
AOI222xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .B1(n_644), .B2(n_645), .C1(n_646), .C2(n_649), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g701 ( .A(n_641), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_641), .B(n_674), .Y(n_727) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g661 ( .A(n_648), .Y(n_661) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
OR2x2_ASAP7_75t_L g766 ( .A(n_650), .B(n_683), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_651), .A2(n_742), .B1(n_744), .B2(n_746), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_658), .B1(n_662), .B2(n_665), .C(n_666), .Y(n_652) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI21xp5_ASAP7_75t_SL g726 ( .A1(n_659), .A2(n_727), .B(n_728), .Y(n_726) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx2_ASAP7_75t_L g674 ( .A(n_660), .Y(n_674) );
AND2x2_ASAP7_75t_L g768 ( .A(n_660), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g752 ( .A(n_664), .Y(n_752) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g681 ( .A(n_670), .B(n_671), .Y(n_681) );
INVx1_ASAP7_75t_L g734 ( .A(n_670), .Y(n_734) );
NOR3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_708), .C(n_730), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_682), .B(n_684), .C(n_689), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_679), .A2(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .B(n_695), .C(n_702), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g713 ( .A(n_696), .Y(n_713) );
INVxp67_ASAP7_75t_SL g738 ( .A(n_697), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_699), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g761 ( .A(n_699), .Y(n_761) );
AND2x2_ASAP7_75t_L g751 ( .A(n_701), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g721 ( .A(n_703), .Y(n_721) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g729 ( .A(n_705), .Y(n_729) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_711), .B(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g750 ( .A1(n_717), .A2(n_751), .B1(n_753), .B2(n_755), .C(n_760), .Y(n_750) );
OAI21xp33_ASAP7_75t_SL g765 ( .A1(n_722), .A2(n_766), .B(n_767), .Y(n_765) );
INVx2_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND4xp25_ASAP7_75t_L g730 ( .A(n_731), .B(n_741), .C(n_750), .D(n_764), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_735), .B1(n_738), .B2(n_739), .Y(n_731) );
AND2x4_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
CKINVDCx11_ASAP7_75t_R g780 ( .A(n_772), .Y(n_780) );
INVx1_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
INVx3_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
INVxp33_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_802), .Y(n_801) );
endmodule