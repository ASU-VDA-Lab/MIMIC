module fake_ariane_468_n_8149 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_33, n_19, n_40, n_106, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_108, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_8149);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_33;
input n_19;
input n_40;
input n_106;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_108;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_8149;

wire n_2752;
wire n_4474;
wire n_3527;
wire n_7329;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_8139;
wire n_416;
wire n_4962;
wire n_1430;
wire n_7832;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_7922;
wire n_7805;
wire n_2790;
wire n_7542;
wire n_2207;
wire n_7053;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_462;
wire n_1131;
wire n_8037;
wire n_5479;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_232;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_6358;
wire n_6293;
wire n_2482;
wire n_1682;
wire n_7001;
wire n_958;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_146;
wire n_4853;
wire n_338;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_7464;
wire n_4260;
wire n_903;
wire n_7626;
wire n_3348;
wire n_239;
wire n_3261;
wire n_1761;
wire n_7965;
wire n_7368;
wire n_1690;
wire n_2807;
wire n_6664;
wire n_7562;
wire n_7534;
wire n_1018;
wire n_7428;
wire n_4512;
wire n_6190;
wire n_4132;
wire n_1364;
wire n_7373;
wire n_2390;
wire n_8068;
wire n_6891;
wire n_4500;
wire n_625;
wire n_2322;
wire n_1107;
wire n_331;
wire n_559;
wire n_2663;
wire n_8097;
wire n_5481;
wire n_6539;
wire n_495;
wire n_8114;
wire n_4824;
wire n_7467;
wire n_350;
wire n_8126;
wire n_381;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_1428;
wire n_1284;
wire n_7526;
wire n_1241;
wire n_4741;
wire n_561;
wire n_4143;
wire n_4273;
wire n_507;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_786;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_6197;
wire n_7200;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_277;
wire n_5691;
wire n_7937;
wire n_3482;
wire n_7490;
wire n_6295;
wire n_5403;
wire n_823;
wire n_1900;
wire n_620;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_587;
wire n_863;
wire n_6992;
wire n_303;
wire n_3960;
wire n_2433;
wire n_352;
wire n_899;
wire n_3975;
wire n_8035;
wire n_5830;
wire n_365;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_334;
wire n_192;
wire n_3325;
wire n_6681;
wire n_661;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_533;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_6542;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_273;
wire n_4505;
wire n_6452;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_7306;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_579;
wire n_7507;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_7215;
wire n_149;
wire n_1213;
wire n_2382;
wire n_7441;
wire n_7379;
wire n_237;
wire n_780;
wire n_5292;
wire n_1918;
wire n_7438;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_3458;
wire n_570;
wire n_5843;
wire n_7874;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_490;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_575;
wire n_7695;
wire n_6156;
wire n_1216;
wire n_4908;
wire n_8098;
wire n_3754;
wire n_5060;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_7331;
wire n_5913;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_7944;
wire n_3841;
wire n_5249;
wire n_249;
wire n_851;
wire n_123;
wire n_444;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_6872;
wire n_6644;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_7607;
wire n_7642;
wire n_1386;
wire n_6236;
wire n_7104;
wire n_8147;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_1842;
wire n_4993;
wire n_7397;
wire n_3678;
wire n_7205;
wire n_366;
wire n_2791;
wire n_1661;
wire n_555;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_7461;
wire n_1692;
wire n_2611;
wire n_8075;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_7638;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_7224;
wire n_6966;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_7259;
wire n_7838;
wire n_5984;
wire n_5204;
wire n_6705;
wire n_6724;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_203;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_150;
wire n_2930;
wire n_7840;
wire n_2745;
wire n_2087;
wire n_619;
wire n_2161;
wire n_746;
wire n_6624;
wire n_1357;
wire n_7888;
wire n_292;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_8108;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_6553;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_6261;
wire n_6659;
wire n_428;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_7583;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_542;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_1087;
wire n_632;
wire n_2388;
wire n_2273;
wire n_8130;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_7488;
wire n_3700;
wire n_7690;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_6206;
wire n_7893;
wire n_2954;
wire n_382;
wire n_489;
wire n_4438;
wire n_6538;
wire n_7966;
wire n_251;
wire n_974;
wire n_506;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_7599;
wire n_7231;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_1447;
wire n_1220;
wire n_7900;
wire n_2019;
wire n_5708;
wire n_8123;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_124;
wire n_5454;
wire n_307;
wire n_1209;
wire n_4254;
wire n_646;
wire n_3438;
wire n_404;
wire n_2625;
wire n_5373;
wire n_7403;
wire n_1578;
wire n_6665;
wire n_3147;
wire n_299;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_133;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_1247;
wire n_6860;
wire n_522;
wire n_1568;
wire n_2919;
wire n_7322;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_367;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_424;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_7963;
wire n_6382;
wire n_670;
wire n_2677;
wire n_4296;
wire n_379;
wire n_138;
wire n_162;
wire n_2483;
wire n_7938;
wire n_5088;
wire n_6615;
wire n_441;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_207;
wire n_720;
wire n_6263;
wire n_1943;
wire n_6731;
wire n_5138;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_194;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_6234;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_5230;
wire n_4555;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_7202;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_5985;
wire n_604;
wire n_478;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_7868;
wire n_3370;
wire n_874;
wire n_7654;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_129;
wire n_126;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_6366;
wire n_1015;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_688;
wire n_7176;
wire n_636;
wire n_1490;
wire n_5552;
wire n_6074;
wire n_7547;
wire n_442;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_8030;
wire n_887;
wire n_2125;
wire n_1156;
wire n_5123;
wire n_4974;
wire n_6689;
wire n_2861;
wire n_7942;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_7527;
wire n_4856;
wire n_2618;
wire n_7948;
wire n_7096;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_5596;
wire n_6482;
wire n_8106;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_616;
wire n_7293;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_7144;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_7316;
wire n_7508;
wire n_3070;
wire n_1005;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_7869;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_6631;
wire n_5889;
wire n_7151;
wire n_3944;
wire n_7762;
wire n_5632;
wire n_4729;
wire n_8002;
wire n_6728;
wire n_1793;
wire n_4446;
wire n_5613;
wire n_4662;
wire n_7472;
wire n_4800;
wire n_1373;
wire n_7075;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_7611;
wire n_7796;
wire n_6508;
wire n_832;
wire n_7989;
wire n_8047;
wire n_744;
wire n_2821;
wire n_3696;
wire n_7936;
wire n_215;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_655;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_2211;
wire n_951;
wire n_8039;
wire n_7546;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_6456;
wire n_5108;
wire n_722;
wire n_7407;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_7481;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_5435;
wire n_6484;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_5476;
wire n_5483;
wire n_7605;
wire n_8090;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_6639;
wire n_358;
wire n_608;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_317;
wire n_3197;
wire n_7423;
wire n_3256;
wire n_1878;
wire n_7375;
wire n_7076;
wire n_7689;
wire n_6344;
wire n_266;
wire n_7736;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_7419;
wire n_811;
wire n_6600;
wire n_7010;
wire n_791;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_480;
wire n_7918;
wire n_642;
wire n_1406;
wire n_5073;
wire n_6555;
wire n_6360;
wire n_4306;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_474;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_386;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_197;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_7346;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_6102;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_6650;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_7385;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_1330;
wire n_906;
wire n_6204;
wire n_2295;
wire n_5225;
wire n_283;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_7148;
wire n_3142;
wire n_7169;
wire n_3129;
wire n_374;
wire n_3495;
wire n_3843;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_7600;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_6946;
wire n_7947;
wire n_5931;
wire n_8146;
wire n_1829;
wire n_4635;
wire n_7847;
wire n_1450;
wire n_5532;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_8027;
wire n_7807;
wire n_1493;
wire n_2911;
wire n_515;
wire n_8063;
wire n_3313;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_7660;
wire n_5365;
wire n_1256;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_6442;
wire n_140;
wire n_6188;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_230;
wire n_3548;
wire n_4906;
wire n_6846;
wire n_4630;
wire n_6840;
wire n_142;
wire n_6645;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_7831;
wire n_8138;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_7455;
wire n_1397;
wire n_5921;
wire n_6247;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_7509;
wire n_6205;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_7497;
wire n_7315;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_7887;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_426;
wire n_6706;
wire n_7431;
wire n_8140;
wire n_398;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_166;
wire n_8117;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_7521;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_8129;
wire n_1291;
wire n_7253;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_7569;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_6551;
wire n_3386;
wire n_400;
wire n_7972;
wire n_7505;
wire n_3921;
wire n_282;
wire n_467;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_7524;
wire n_4196;
wire n_1197;
wire n_7318;
wire n_2613;
wire n_7411;
wire n_7326;
wire n_5667;
wire n_168;
wire n_1517;
wire n_2647;
wire n_8005;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_7573;
wire n_6630;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_6798;
wire n_5999;
wire n_1504;
wire n_2110;
wire n_7498;
wire n_7895;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_3822;
wire n_889;
wire n_7453;
wire n_4355;
wire n_3818;
wire n_7932;
wire n_7890;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6403;
wire n_3497;
wire n_6395;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_565;
wire n_3927;
wire n_6141;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_452;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_6944;
wire n_4452;
wire n_284;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_7240;
wire n_409;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_1056;
wire n_526;
wire n_5584;
wire n_674;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_6559;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_6248;
wire n_6541;
wire n_848;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_629;
wire n_4733;
wire n_7927;
wire n_161;
wire n_1814;
wire n_7219;
wire n_2441;
wire n_8081;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_216;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_7402;
wire n_6351;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_7382;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_7767;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_7510;
wire n_3786;
wire n_875;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_7434;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_7691;
wire n_296;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_6744;
wire n_3645;
wire n_793;
wire n_5705;
wire n_6927;
wire n_7335;
wire n_132;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_7735;
wire n_6116;
wire n_8074;
wire n_494;
wire n_3550;
wire n_7956;
wire n_5510;
wire n_7495;
wire n_7651;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_185;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_972;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_164;
wire n_2843;
wire n_3714;
wire n_184;
wire n_7671;
wire n_4832;
wire n_8033;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_118;
wire n_1679;
wire n_5834;
wire n_7926;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_6495;
wire n_7528;
wire n_6209;
wire n_4672;
wire n_8094;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_7413;
wire n_7993;
wire n_7821;
wire n_160;
wire n_7620;
wire n_119;
wire n_1008;
wire n_3963;
wire n_581;
wire n_3091;
wire n_6274;
wire n_1024;
wire n_176;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_6237;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_7343;
wire n_5982;
wire n_1775;
wire n_908;
wire n_1036;
wire n_7109;
wire n_8028;
wire n_341;
wire n_4083;
wire n_1270;
wire n_109;
wire n_1272;
wire n_549;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_6809;
wire n_6099;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_244;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_6716;
wire n_3565;
wire n_7885;
wire n_6905;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_5824;
wire n_8025;
wire n_5354;
wire n_2453;
wire n_7898;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_3040;
wire n_4230;
wire n_6899;
wire n_7980;
wire n_7817;
wire n_6413;
wire n_445;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_7299;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_8029;
wire n_2215;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_1261;
wire n_7249;
wire n_5763;
wire n_3633;
wire n_857;
wire n_363;
wire n_6061;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_5701;
wire n_7002;
wire n_1064;
wire n_633;
wire n_1446;
wire n_1701;
wire n_6273;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_731;
wire n_1813;
wire n_315;
wire n_2997;
wire n_7018;
wire n_1573;
wire n_6746;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_6174;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_5907;
wire n_784;
wire n_4339;
wire n_7297;
wire n_7730;
wire n_8134;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4169;
wire n_4024;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_3632;
wire n_309;
wire n_1344;
wire n_115;
wire n_485;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_435;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_840;
wire n_2324;
wire n_6575;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_2139;
wire n_7613;
wire n_7995;
wire n_8113;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_7140;
wire n_614;
wire n_4066;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_3303;
wire n_7910;
wire n_6592;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_248;
wire n_7741;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_228;
wire n_6668;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_7698;
wire n_1875;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_1150;
wire n_7800;
wire n_6336;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_7835;
wire n_1136;
wire n_458;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_7415;
wire n_5399;
wire n_658;
wire n_362;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_8016;
wire n_3872;
wire n_5760;
wire n_7747;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_7552;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_5844;
wire n_6298;
wire n_8132;
wire n_7650;
wire n_3441;
wire n_199;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_708;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_7635;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_6525;
wire n_3555;
wire n_5938;
wire n_7274;
wire n_3534;
wire n_450;
wire n_4548;
wire n_7819;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_7788;
wire n_6974;
wire n_1168;
wire n_4663;
wire n_219;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_415;
wire n_4686;
wire n_2384;
wire n_7794;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_7630;
wire n_4161;
wire n_110;
wire n_304;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6951;
wire n_6963;
wire n_1581;
wire n_946;
wire n_757;
wire n_5355;
wire n_2047;
wire n_3058;
wire n_375;
wire n_113;
wire n_1655;
wire n_3398;
wire n_1146;
wire n_3709;
wire n_6284;
wire n_998;
wire n_3592;
wire n_5321;
wire n_7454;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_5915;
wire n_7276;
wire n_174;
wire n_6379;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_925;
wire n_7753;
wire n_6834;
wire n_2880;
wire n_1313;
wire n_3722;
wire n_1001;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_719;
wire n_7541;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_7913;
wire n_8020;
wire n_7946;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_6471;
wire n_6949;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_6760;
wire n_2940;
wire n_548;
wire n_3427;
wire n_3162;
wire n_5966;
wire n_5569;
wire n_4591;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_2491;
wire n_7920;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_1820;
wire n_7841;
wire n_7160;
wire n_7324;
wire n_6046;
wire n_7054;
wire n_1233;
wire n_4493;
wire n_6055;
wire n_7161;
wire n_1808;
wire n_6364;
wire n_6091;
wire n_6348;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_8041;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_886;
wire n_7837;
wire n_359;
wire n_6788;
wire n_1308;
wire n_6144;
wire n_1451;
wire n_1487;
wire n_675;
wire n_5528;
wire n_7806;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_8076;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_7676;
wire n_2334;
wire n_5467;
wire n_7241;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_6285;
wire n_610;
wire n_7644;
wire n_4602;
wire n_1713;
wire n_7816;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_7430;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_7269;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_214;
wire n_4103;
wire n_2529;
wire n_8101;
wire n_2374;
wire n_5439;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_137;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_7879;
wire n_6607;
wire n_4439;
wire n_520;
wire n_870;
wire n_4985;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_2844;
wire n_402;
wire n_1979;
wire n_6616;
wire n_6719;
wire n_829;
wire n_4814;
wire n_8019;
wire n_339;
wire n_6178;
wire n_6677;
wire n_2221;
wire n_7875;
wire n_5502;
wire n_1283;
wire n_7550;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_2442;
wire n_7238;
wire n_6862;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_7292;
wire n_242;
wire n_645;
wire n_7804;
wire n_5098;
wire n_721;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_6443;
wire n_1276;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_7248;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_8040;
wire n_5466;
wire n_1528;
wire n_6941;
wire n_7239;
wire n_6552;
wire n_7826;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_8102;
wire n_3999;
wire n_518;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_7971;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_6531;
wire n_3571;
wire n_238;
wire n_4576;
wire n_7577;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_8144;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_7513;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_7812;
wire n_5330;
wire n_6935;
wire n_1560;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_8058;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_6386;
wire n_2722;
wire n_3728;
wire n_6596;
wire n_612;
wire n_333;
wire n_5107;
wire n_7165;
wire n_512;
wire n_5067;
wire n_4680;
wire n_6830;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_6510;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_6781;
wire n_7667;
wire n_4593;
wire n_8024;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_461;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_8107;
wire n_2981;
wire n_225;
wire n_1006;
wire n_546;
wire n_4995;
wire n_1159;
wire n_5873;
wire n_6514;
wire n_4498;
wire n_772;
wire n_6741;
wire n_1245;
wire n_6434;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_6593;
wire n_676;
wire n_7827;
wire n_3758;
wire n_7631;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_212;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_8122;
wire n_2426;
wire n_652;
wire n_6947;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_798;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_912;
wire n_6375;
wire n_460;
wire n_7781;
wire n_4786;
wire n_6042;
wire n_5203;
wire n_7908;
wire n_7091;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_3159;
wire n_6315;
wire n_7855;
wire n_2855;
wire n_794;
wire n_2848;
wire n_7886;
wire n_7675;
wire n_6775;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_288;
wire n_1292;
wire n_7774;
wire n_6970;
wire n_1026;
wire n_6948;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_306;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_7381;
wire n_5804;
wire n_3240;
wire n_7999;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_7873;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_5992;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_5684;
wire n_1399;
wire n_7228;
wire n_5981;
wire n_7784;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_7713;
wire n_6623;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_1226;
wire n_2224;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_5444;
wire n_3980;
wire n_8031;
wire n_3257;
wire n_5737;
wire n_8015;
wire n_425;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_6390;
wire n_7640;
wire n_2302;
wire n_6799;
wire n_3014;
wire n_7912;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_397;
wire n_3375;
wire n_2768;
wire n_351;
wire n_155;
wire n_5661;
wire n_3760;
wire n_7641;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_7949;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_1020;
wire n_7764;
wire n_172;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_8128;
wire n_7520;
wire n_5314;
wire n_7616;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_6271;
wire n_7235;
wire n_2511;
wire n_564;
wire n_6572;
wire n_3981;
wire n_7271;
wire n_2681;
wire n_7222;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_345;
wire n_6930;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_130;
wire n_6387;
wire n_466;
wire n_4201;
wire n_346;
wire n_6470;
wire n_7206;
wire n_552;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_264;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_7383;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_6826;
wire n_1217;
wire n_327;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_7854;
wire n_926;
wire n_2296;
wire n_5735;
wire n_7959;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_7897;
wire n_186;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_6865;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_7132;
wire n_1570;
wire n_7533;
wire n_3377;
wire n_6722;
wire n_1518;
wire n_6420;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_855;
wire n_2059;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_1287;
wire n_1611;
wire n_120;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_6981;
wire n_4870;
wire n_7776;
wire n_4818;
wire n_8001;
wire n_7436;
wire n_7020;
wire n_5935;
wire n_8064;
wire n_6696;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_529;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_7978;
wire n_5488;
wire n_1105;
wire n_6900;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_8131;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_7694;
wire n_5832;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_983;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_699;
wire n_3542;
wire n_301;
wire n_3263;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_325;
wire n_1740;
wire n_5016;
wire n_6011;
wire n_4616;
wire n_7465;
wire n_5470;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_729;
wire n_6222;
wire n_2218;
wire n_1122;
wire n_7760;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_6969;
wire n_390;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_6587;
wire n_6688;
wire n_6505;
wire n_5362;
wire n_388;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_7629;
wire n_6987;
wire n_877;
wire n_3995;
wire n_7567;
wire n_3908;
wire n_6453;
wire n_6308;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_7449;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_6187;
wire n_735;
wire n_6597;
wire n_4844;
wire n_6220;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_7479;
wire n_7882;
wire n_1649;
wire n_2470;
wire n_7517;
wire n_1297;
wire n_3551;
wire n_417;
wire n_1708;
wire n_5037;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_8070;
wire n_4525;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_7878;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_278;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_842;
wire n_148;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_6547;
wire n_7177;
wire n_7902;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_476;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_8054;
wire n_982;
wire n_3791;
wire n_915;
wire n_6478;
wire n_2008;
wire n_454;
wire n_298;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_6906;
wire n_403;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_606;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_7818;
wire n_509;
wire n_7645;
wire n_5385;
wire n_7482;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_7907;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_521;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_7862;
wire n_3735;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_1513;
wire n_1527;
wire n_3656;
wire n_7721;
wire n_4524;
wire n_8061;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_6999;
wire n_8086;
wire n_8072;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_7539;
wire n_6440;
wire n_4977;
wire n_2492;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_241;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_5936;
wire n_595;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_7830;
wire n_8050;
wire n_3124;
wire n_3811;
wire n_295;
wire n_4200;
wire n_190;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_463;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_469;
wire n_726;
wire n_5504;
wire n_878;
wire n_7348;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_8010;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_6464;
wire n_5129;
wire n_806;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_1616;
wire n_7935;
wire n_2416;
wire n_8143;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_7933;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_349;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_6850;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_7743;
wire n_5389;
wire n_4764;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_6550;
wire n_6656;
wire n_6972;
wire n_3591;
wire n_198;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_7043;
wire n_7986;
wire n_3317;
wire n_8049;
wire n_7266;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_554;
wire n_4420;
wire n_7996;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_354;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_594;
wire n_7035;
wire n_4173;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_422;
wire n_1269;
wire n_7442;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_6258;
wire n_1288;
wire n_7939;
wire n_7715;
wire n_2173;
wire n_3982;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_1143;
wire n_3973;
wire n_8052;
wire n_4799;
wire n_8082;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_7699;
wire n_1153;
wire n_271;
wire n_465;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_562;
wire n_2020;
wire n_7580;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_510;
wire n_5911;
wire n_7340;
wire n_8080;
wire n_256;
wire n_3600;
wire n_7303;
wire n_1023;
wire n_914;
wire n_7870;
wire n_689;
wire n_6139;
wire n_7568;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_497;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_455;
wire n_588;
wire n_638;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_7207;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_5841;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_413;
wire n_2935;
wire n_4246;
wire n_715;
wire n_7618;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_617;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_8008;
wire n_7633;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_2592;
wire n_3490;
wire n_7280;
wire n_962;
wire n_5043;
wire n_7339;
wire n_7597;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_7768;
wire n_918;
wire n_1968;
wire n_5645;
wire n_639;
wire n_6455;
wire n_673;
wire n_5020;
wire n_2842;
wire n_7615;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_6183;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_6003;
wire n_5443;
wire n_8133;
wire n_7612;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_5631;
wire n_3481;
wire n_280;
wire n_6994;
wire n_7401;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_6185;
wire n_692;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_223;
wire n_2150;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_6695;
wire n_7529;
wire n_3354;
wire n_5608;
wire n_6501;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_6467;
wire n_2231;
wire n_4212;
wire n_622;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_8088;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_792;
wire n_1262;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_6213;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_229;
wire n_923;
wire n_1124;
wire n_7872;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_7958;
wire n_2282;
wire n_4605;
wire n_8118;
wire n_981;
wire n_4649;
wire n_3873;
wire n_5747;
wire n_7101;
wire n_1204;
wire n_7843;
wire n_994;
wire n_2428;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_7578;
wire n_3410;
wire n_5415;
wire n_856;
wire n_7261;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_6993;
wire n_508;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_8100;
wire n_1858;
wire n_353;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_6767;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6558;
wire n_6755;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_7263;
wire n_3782;
wire n_1317;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_7688;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7925;
wire n_7310;
wire n_294;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_7585;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_7772;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_679;
wire n_220;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_7514;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_6105;
wire n_387;
wire n_826;
wire n_5512;
wire n_7738;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_7609;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_607;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_7282;
wire n_372;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_7921;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_7489;
wire n_6331;
wire n_5308;
wire n_311;
wire n_4434;
wire n_5068;
wire n_7863;
wire n_6493;
wire n_7363;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_7968;
wire n_6023;
wire n_7820;
wire n_269;
wire n_816;
wire n_7833;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_7750;
wire n_5057;
wire n_446;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_7588;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_7697;
wire n_5887;
wire n_7808;
wire n_3068;
wire n_1629;
wire n_7603;
wire n_1094;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_3002;
wire n_7192;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_8012;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_7988;
wire n_550;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_6450;
wire n_1152;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_671;
wire n_8105;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_7943;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_7377;
wire n_4392;
wire n_3103;
wire n_488;
wire n_6064;
wire n_505;
wire n_2048;
wire n_7723;
wire n_498;
wire n_3028;
wire n_4691;
wire n_7904;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_684;
wire n_5461;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_6164;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_6330;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_838;
wire n_1941;
wire n_7045;
wire n_175;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_7777;
wire n_4258;
wire n_5756;
wire n_310;
wire n_7693;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_8078;
wire n_2097;
wire n_662;
wire n_3461;
wire n_7682;
wire n_7300;
wire n_1410;
wire n_939;
wire n_2297;
wire n_6861;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_7558;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_572;
wire n_8103;
wire n_1983;
wire n_7798;
wire n_4767;
wire n_4569;
wire n_948;
wire n_448;
wire n_6528;
wire n_5144;
wire n_3820;
wire n_6895;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_6472;
wire n_3763;
wire n_933;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_492;
wire n_252;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_7672;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_389;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_5751;
wire n_626;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_7712;
wire n_6885;
wire n_7681;
wire n_5039;
wire n_1818;
wire n_6580;
wire n_6613;
wire n_4265;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_7491;
wire n_265;
wire n_1583;
wire n_4612;
wire n_5997;
wire n_5375;
wire n_5438;
wire n_7150;
wire n_7954;
wire n_7974;
wire n_1264;
wire n_6530;
wire n_6602;
wire n_7915;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_6135;
wire n_246;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_6942;
wire n_7860;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_7357;
wire n_8112;
wire n_8060;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_8096;
wire n_7336;
wire n_5932;
wire n_289;
wire n_112;
wire n_6598;
wire n_6795;
wire n_6121;
wire n_457;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_6001;
wire n_411;
wire n_4971;
wire n_2095;
wire n_7493;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_357;
wire n_3041;
wire n_412;
wire n_5823;
wire n_1421;
wire n_2423;
wire n_2208;
wire n_5422;
wire n_5944;
wire n_6989;
wire n_8145;
wire n_6299;
wire n_7424;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_573;
wire n_2823;
wire n_7273;
wire n_7901;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_7149;
wire n_589;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_1383;
wire n_603;
wire n_8055;
wire n_373;
wire n_4259;
wire n_5870;
wire n_7909;
wire n_2030;
wire n_6053;
wire n_850;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_245;
wire n_319;
wire n_6758;
wire n_2407;
wire n_690;
wire n_5367;
wire n_525;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_5601;
wire n_4965;
wire n_7601;
wire n_3742;
wire n_1837;
wire n_7033;
wire n_6010;
wire n_4178;
wire n_189;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_7596;
wire n_5294;
wire n_5570;
wire n_6411;
wire n_2731;
wire n_3703;
wire n_5670;
wire n_5411;
wire n_1246;
wire n_5265;
wire n_5955;
wire n_7549;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_3435;
wire n_410;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_6918;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_568;
wire n_4796;
wire n_1088;
wire n_7138;
wire n_766;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_7976;
wire n_377;
wire n_2750;
wire n_2547;
wire n_7617;
wire n_279;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_8062;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_7700;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_500;
wire n_665;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_5575;
wire n_6654;
wire n_7661;
wire n_672;
wire n_4968;
wire n_7801;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_4038;
wire n_3856;
wire n_5316;
wire n_7876;
wire n_2735;
wire n_953;
wire n_4214;
wire n_143;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_557;
wire n_3419;
wire n_7323;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_6517;
wire n_795;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_8048;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_7929;
wire n_486;
wire n_2782;
wire n_569;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_7755;
wire n_6504;
wire n_4176;
wire n_7556;
wire n_222;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_7216;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_8043;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_5845;
wire n_4608;
wire n_6691;
wire n_432;
wire n_293;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_206;
wire n_2332;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_611;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_136;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_300;
wire n_6025;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_7962;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_376;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_6771;
wire n_7905;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_7476;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_209;
wire n_5503;
wire n_5718;
wire n_1461;
wire n_5240;
wire n_7208;
wire n_7718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_6567;
wire n_503;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_380;
wire n_3119;
wire n_6671;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_7632;
wire n_4394;
wire n_257;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_475;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_8073;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_577;
wire n_5610;
wire n_407;
wire n_916;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_7265;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_5808;
wire n_1182;
wire n_6527;
wire n_4594;
wire n_8045;
wire n_7289;
wire n_7538;
wire n_2748;
wire n_4642;
wire n_6913;
wire n_1376;
wire n_7473;
wire n_7242;
wire n_6533;
wire n_513;
wire n_179;
wire n_7164;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_8022;
wire n_3544;
wire n_6845;
wire n_5300;
wire n_7853;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_436;
wire n_5770;
wire n_7483;
wire n_5710;
wire n_324;
wire n_1491;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_111;
wire n_274;
wire n_1083;
wire n_5799;
wire n_5333;
wire n_6265;
wire n_4914;
wire n_3510;
wire n_7046;
wire n_7834;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_563;
wire n_2219;
wire n_6148;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_990;
wire n_6357;
wire n_867;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_7811;
wire n_4285;
wire n_7097;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_7880;
wire n_712;
wire n_909;
wire n_6713;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_7851;
wire n_2220;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_6108;
wire n_7664;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_7332;
wire n_5862;
wire n_471;
wire n_7477;
wire n_1914;
wire n_2253;
wire n_7468;
wire n_5886;
wire n_7714;
wire n_7899;
wire n_6415;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_7845;
wire n_347;
wire n_2434;
wire n_183;
wire n_1234;
wire n_3936;
wire n_479;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_7858;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_6513;
wire n_6392;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_6720;
wire n_5883;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_370;
wire n_7680;
wire n_5630;
wire n_6666;
wire n_286;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_6815;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_7710;
wire n_5394;
wire n_4751;
wire n_5975;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_7061;
wire n_8104;
wire n_7066;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_8014;
wire n_4122;
wire n_6661;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_4952;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_7783;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_487;
wire n_4728;
wire n_7171;
wire n_7990;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_7003;
wire n_8137;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_6302;
wire n_3863;
wire n_2327;
wire n_158;
wire n_3882;
wire n_3916;
wire n_6922;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_405;
wire n_3332;
wire n_8069;
wire n_7501;
wire n_320;
wire n_6432;
wire n_7984;
wire n_2055;
wire n_2998;
wire n_7366;
wire n_1423;
wire n_4359;
wire n_481;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_7589;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_218;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_1798;
wire n_8091;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_6699;
wire n_547;
wire n_439;
wire n_677;
wire n_3983;
wire n_703;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_7511;
wire n_326;
wire n_227;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_6957;
wire n_5074;
wire n_7917;
wire n_3788;
wire n_3939;
wire n_727;
wire n_590;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_6694;
wire n_545;
wire n_2496;
wire n_3260;
wire n_536;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_1602;
wire n_7422;
wire n_3139;
wire n_427;
wire n_3801;
wire n_5681;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_7621;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_163;
wire n_2716;
wire n_6441;
wire n_7158;
wire n_7572;
wire n_314;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_7500;
wire n_1202;
wire n_4084;
wire n_627;
wire n_7985;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_233;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_321;
wire n_6662;
wire n_7494;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_6433;
wire n_1763;
wire n_6200;
wire n_5641;
wire n_8071;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_5657;
wire n_297;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_178;
wire n_551;
wire n_4521;
wire n_6956;
wire n_7587;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_7704;
wire n_5420;
wire n_6497;
wire n_7865;
wire n_2283;
wire n_5206;
wire n_582;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_534;
wire n_2508;
wire n_3186;
wire n_6701;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_560;
wire n_890;
wire n_3626;
wire n_451;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_7881;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_535;
wire n_4565;
wire n_7032;
wire n_3392;
wire n_1800;
wire n_7198;
wire n_6884;
wire n_7752;
wire n_5081;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_7953;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_8046;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_6362;
wire n_4328;
wire n_1854;
wire n_666;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_7126;
wire n_5867;
wire n_456;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_7496;
wire n_6430;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_342;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_7196;
wire n_2614;
wire n_7360;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_6678;
wire n_7982;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_6385;
wire n_1668;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_8032;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_8036;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_618;
wire n_1191;
wire n_4535;
wire n_7518;
wire n_4385;
wire n_7779;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_7575;
wire n_2337;
wire n_7073;
wire n_8092;
wire n_1786;
wire n_6309;
wire n_3732;
wire n_211;
wire n_1804;
wire n_408;
wire n_8135;
wire n_6519;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_5989;
wire n_4766;
wire n_592;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_7349;
wire n_1929;
wire n_4319;
wire n_6585;
wire n_7786;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_7579;
wire n_7122;
wire n_4874;
wire n_180;
wire n_2656;
wire n_4904;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_640;
wire n_1733;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_7624;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_7828;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_7543;
wire n_5475;
wire n_8042;
wire n_7727;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_5431;
wire n_643;
wire n_8034;
wire n_226;
wire n_7778;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_7019;
wire n_682;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_7702;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_686;
wire n_1154;
wire n_584;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_6685;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_7952;
wire n_7347;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_7791;
wire n_6971;
wire n_3336;
wire n_7739;
wire n_396;
wire n_7945;
wire n_7656;
wire n_5903;
wire n_7199;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_6549;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_6683;
wire n_3067;
wire n_154;
wire n_3809;
wire n_4921;
wire n_473;
wire n_1852;
wire n_801;
wire n_5912;
wire n_5745;
wire n_7923;
wire n_6086;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_272;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_7610;
wire n_7107;
wire n_4561;
wire n_1541;
wire n_597;
wire n_3291;
wire n_7456;
wire n_8095;
wire n_7369;
wire n_1472;
wire n_1050;
wire n_7548;
wire n_2578;
wire n_152;
wire n_1201;
wire n_7598;
wire n_1185;
wire n_2475;
wire n_7250;
wire n_7823;
wire n_4715;
wire n_6157;
wire n_2715;
wire n_335;
wire n_2665;
wire n_4879;
wire n_344;
wire n_5044;
wire n_210;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_6676;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_224;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_7525;
wire n_4418;
wire n_7924;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_276;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_6923;
wire n_7649;
wire n_843;
wire n_8009;
wire n_3358;
wire n_6704;
wire n_7634;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_7406;
wire n_4682;
wire n_1128;
wire n_6673;
wire n_2419;
wire n_2330;
wire n_6534;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_1440;
wire n_6246;
wire n_1370;
wire n_305;
wire n_5005;
wire n_6126;
wire n_7372;
wire n_1549;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_7844;
wire n_5207;
wire n_7934;
wire n_361;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_5474;
wire n_2767;
wire n_7009;
wire n_3376;
wire n_181;
wire n_7371;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_683;
wire n_7463;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_5700;
wire n_5755;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_660;
wire n_464;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_6723;
wire n_7398;
wire n_1038;
wire n_3723;
wire n_7941;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_414;
wire n_571;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_613;
wire n_1022;
wire n_5465;
wire n_171;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_6184;
wire n_8018;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_7083;
wire n_316;
wire n_125;
wire n_1973;
wire n_1444;
wire n_820;
wire n_254;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_7701;
wire n_7969;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_6312;
wire n_4577;
wire n_7683;
wire n_532;
wire n_2154;
wire n_7669;
wire n_1986;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_8023;
wire n_7330;
wire n_6007;
wire n_621;
wire n_6734;
wire n_6535;
wire n_8053;
wire n_8059;
wire n_1772;
wire n_6879;
wire n_493;
wire n_1311;
wire n_3106;
wire n_6208;
wire n_7190;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_7692;
wire n_697;
wire n_4620;
wire n_5397;
wire n_6255;
wire n_6457;
wire n_4924;
wire n_4044;
wire n_6270;
wire n_2305;
wire n_5996;
wire n_880;
wire n_5566;
wire n_3304;
wire n_7288;
wire n_4388;
wire n_7362;
wire n_7237;
wire n_7082;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_739;
wire n_1028;
wire n_530;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_7042;
wire n_2809;
wire n_5652;
wire n_975;
wire n_1645;
wire n_5805;
wire n_7304;
wire n_932;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_8077;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_7754;
wire n_3178;
wire n_268;
wire n_7023;
wire n_2251;
wire n_5842;
wire n_5758;
wire n_3100;
wire n_3721;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_7981;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_191;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_8109;
wire n_116;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_7378;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_7877;
wire n_7787;
wire n_7836;
wire n_8007;
wire n_2387;
wire n_4318;
wire n_332;
wire n_5227;
wire n_830;
wire n_5902;
wire n_987;
wire n_2510;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_6764;
wire n_7871;
wire n_541;
wire n_499;
wire n_2639;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_6215;
wire n_4554;
wire n_7571;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_6955;
wire n_7563;
wire n_5952;
wire n_7180;
wire n_2086;
wire n_1926;
wire n_6569;
wire n_1630;
wire n_7919;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_443;
wire n_3431;
wire n_3355;
wire n_7031;
wire n_1738;
wire n_5716;
wire n_406;
wire n_3897;
wire n_7103;
wire n_139;
wire n_6605;
wire n_1735;
wire n_391;
wire n_5888;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_6832;
wire n_5980;
wire n_956;
wire n_765;
wire n_4092;
wire n_122;
wire n_4875;
wire n_7771;
wire n_4255;
wire n_2758;
wire n_385;
wire n_6544;
wire n_6469;
wire n_5036;
wire n_1271;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_399;
wire n_7130;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_2471;
wire n_7134;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_1551;
wire n_5271;
wire n_4849;
wire n_2039;
wire n_7133;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_6289;
wire n_6651;
wire n_3838;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_8067;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_7706;
wire n_7813;
wire n_8142;
wire n_2420;
wire n_7992;
wire n_7643;
wire n_153;
wire n_648;
wire n_6836;
wire n_3273;
wire n_2918;
wire n_6595;
wire n_835;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_401;
wire n_7628;
wire n_1792;
wire n_5628;
wire n_504;
wire n_5245;
wire n_2062;
wire n_483;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_6035;
wire n_839;
wire n_1754;
wire n_7236;
wire n_4833;
wire n_3394;
wire n_6405;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_6786;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_8110;
wire n_5072;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_2260;
wire n_323;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_7519;
wire n_7802;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_7457;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_6416;
wire n_654;
wire n_2933;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_6214;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_7049;
wire n_7884;
wire n_6945;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_7749;
wire n_7592;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_539;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_7914;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_4390;
wire n_459;
wire n_1782;
wire n_7892;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4609;
wire n_4361;
wire n_7325;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_723;
wire n_1393;
wire n_7674;
wire n_6175;
wire n_6445;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_6198;
wire n_5172;
wire n_881;
wire n_1019;
wire n_1477;
wire n_6499;
wire n_1982;
wire n_7983;
wire n_641;
wire n_5311;
wire n_910;
wire n_290;
wire n_5164;
wire n_4964;
wire n_6842;
wire n_4700;
wire n_4002;
wire n_217;
wire n_7361;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_201;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_1043;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_255;
wire n_2869;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_1613;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_196;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_231;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_664;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_6732;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_544;
wire n_7646;
wire n_3779;
wire n_599;
wire n_6982;
wire n_537;
wire n_1063;
wire n_7291;
wire n_991;
wire n_2275;
wire n_7668;
wire n_7435;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_583;
wire n_1000;
wire n_313;
wire n_4868;
wire n_7017;
wire n_378;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_4465;
wire n_8127;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_7861;
wire n_472;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_7889;
wire n_208;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_7554;
wire n_275;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_7648;
wire n_147;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_7653;
wire n_6400;
wire n_1644;
wire n_7846;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_131;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_250;
wire n_773;
wire n_5135;
wire n_7551;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_718;
wire n_1434;
wire n_8093;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_7737;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_523;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_6621;
wire n_6851;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_7606;
wire n_7420;
wire n_8115;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_484;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_796;
wire n_127;
wire n_531;
wire n_1374;
wire n_2089;
wire n_7896;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_5900;
wire n_7319;
wire n_1486;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_6819;
wire n_6122;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_423;
wire n_4085;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_5851;
wire n_7516;
wire n_6317;
wire n_6928;
wire n_6707;
wire n_7244;
wire n_187;
wire n_1463;
wire n_4626;
wire n_7625;
wire n_4997;
wire n_5065;
wire n_6806;
wire n_924;
wire n_7991;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_7857;
wire n_7970;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_117;
wire n_7154;
wire n_524;
wire n_634;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_5173;
wire n_4683;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_7175;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_7163;
wire n_3797;
wire n_1836;
wire n_7027;
wire n_3416;
wire n_5861;
wire n_4600;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_7964;
wire n_5749;
wire n_6320;
wire n_6316;
wire n_419;
wire n_7068;
wire n_2908;
wire n_270;
wire n_4106;
wire n_285;
wire n_2156;
wire n_1184;
wire n_202;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_7327;
wire n_1277;
wire n_1746;
wire n_6610;
wire n_1062;
wire n_5998;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_167;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_6752;
wire n_6959;
wire n_6250;
wire n_3283;
wire n_259;
wire n_7317;
wire n_4331;
wire n_4159;
wire n_7864;
wire n_3451;
wire n_8051;
wire n_4734;
wire n_6675;
wire n_7955;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_7384;
wire n_267;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_5678;
wire n_6561;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_7512;
wire n_1718;
wire n_7814;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_200;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_7152;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_7223;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_7761;
wire n_8141;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_8004;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_7437;
wire n_6489;
wire n_5310;
wire n_2769;
wire n_438;
wire n_1548;
wire n_4987;
wire n_6714;
wire n_440;
wire n_7849;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_7417;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_1544;
wire n_6620;
wire n_6791;
wire n_4540;
wire n_6821;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_1354;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_7859;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_491;
wire n_1595;
wire n_8017;
wire n_1142;
wire n_5477;
wire n_260;
wire n_2727;
wire n_942;
wire n_7523;
wire n_5234;
wire n_1416;
wire n_6890;
wire n_7559;
wire n_7576;
wire n_6988;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_8000;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_7769;
wire n_7257;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_287;
wire n_3191;
wire n_1716;
wire n_302;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_7081;
wire n_7742;
wire n_5253;
wire n_3588;
wire n_355;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_135;
wire n_3095;
wire n_947;
wire n_7341;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_6256;
wire n_4775;
wire n_482;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_7264;
wire n_7842;
wire n_2499;
wire n_2549;
wire n_6648;
wire n_7492;
wire n_804;
wire n_6649;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_3885;
wire n_955;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_514;
wire n_6431;
wire n_418;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_669;
wire n_5580;
wire n_5215;
wire n_337;
wire n_437;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_615;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_517;
wire n_8124;
wire n_3604;
wire n_5430;
wire n_6041;
wire n_824;
wire n_159;
wire n_7997;
wire n_5659;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_144;
wire n_3792;
wire n_7950;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_7793;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_470;
wire n_3021;
wire n_7746;
wire n_477;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_7570;
wire n_2898;
wire n_1825;
wire n_6912;
wire n_3567;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_1731;
wire n_799;
wire n_7894;
wire n_1147;
wire n_7957;
wire n_2378;
wire n_5530;
wire n_6718;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_7121;
wire n_7531;
wire n_6410;
wire n_356;
wire n_6473;
wire n_8087;
wire n_4056;
wire n_4806;
wire n_7961;
wire n_1674;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_6857;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_6975;
wire n_7763;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_205;
wire n_7703;
wire n_7928;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_713;
wire n_3179;
wire n_598;
wire n_6622;
wire n_5522;
wire n_7665;
wire n_4836;
wire n_7677;
wire n_5262;
wire n_3889;
wire n_3262;
wire n_5319;
wire n_927;
wire n_7469;
wire n_261;
wire n_3699;
wire n_6118;
wire n_706;
wire n_2120;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_1419;
wire n_3816;
wire n_8099;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_4207;
wire n_8085;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_348;
wire n_2312;
wire n_7203;
wire n_7797;
wire n_1826;
wire n_5943;
wire n_6556;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_7128;
wire n_5335;
wire n_1259;
wire n_6365;
wire n_7111;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_7057;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_6167;
wire n_3200;
wire n_3642;
wire n_145;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_7278;
wire n_6772;
wire n_7088;
wire n_7799;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_7048;
wire n_7979;
wire n_6617;
wire n_553;
wire n_7725;
wire n_814;
wire n_578;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_647;
wire n_2027;
wire n_2932;
wire n_6217;
wire n_600;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_5455;
wire n_2195;
wire n_3922;
wire n_502;
wire n_6777;
wire n_6742;
wire n_1467;
wire n_7447;
wire n_5209;
wire n_247;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_6479;
wire n_5099;
wire n_681;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_7365;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_5022;
wire n_8089;
wire n_6370;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_3009;
wire n_777;
wire n_7095;
wire n_7390;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_1132;
wire n_8125;
wire n_501;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_6712;
wire n_7530;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_7471;
wire n_6465;
wire n_221;
wire n_5673;
wire n_861;
wire n_5814;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_8011;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_281;
wire n_3326;
wire n_262;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_8065;
wire n_527;
wire n_2949;
wire n_7008;
wire n_6468;
wire n_7709;
wire n_4269;
wire n_1927;
wire n_7540;
wire n_7581;
wire n_343;
wire n_1222;
wire n_7139;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_7782;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_6483;
wire n_1572;
wire n_7770;
wire n_4463;
wire n_5357;
wire n_7173;
wire n_3648;
wire n_6576;
wire n_6810;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_8026;
wire n_6667;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_6305;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_7751;
wire n_7951;
wire n_657;
wire n_7060;
wire n_3924;
wire n_3997;
wire n_7591;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_6750;
wire n_7444;
wire n_7911;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_2306;
wire n_7790;
wire n_2071;
wire n_7426;
wire n_430;
wire n_3953;
wire n_7502;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_6855;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_5768;
wire n_1342;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_8120;
wire n_852;
wire n_2916;
wire n_7252;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_4192;
wire n_8003;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_7065;
wire n_1466;
wire n_8083;
wire n_6177;
wire n_8057;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_7367;
wire n_7267;
wire n_7405;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_6825;
wire n_7614;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_134;
wire n_4035;
wire n_6952;
wire n_1480;
wire n_3670;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_6218;
wire n_7685;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_157;
wire n_7619;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_624;
wire n_5577;
wire n_876;
wire n_5872;
wire n_7883;
wire n_6692;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_602;
wire n_854;
wire n_2091;
wire n_393;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_7270;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_7731;
wire n_6626;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_7034;
wire n_3694;
wire n_6854;
wire n_7940;
wire n_771;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_421;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_7537;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_7458;
wire n_1824;
wire n_7740;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_819;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_3543;
wire n_7179;
wire n_1776;
wire n_3448;
wire n_7433;
wire n_4279;
wire n_605;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_6334;
wire n_6257;
wire n_4152;
wire n_6874;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_7987;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_6377;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_7272;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_151;
wire n_7906;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_7765;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_6511;
wire n_7815;
wire n_1052;
wire n_4732;
wire n_2203;
wire n_2076;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_4969;
wire n_8121;
wire n_5252;
wire n_5777;
wire n_7785;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_566;
wire n_7728;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_169;
wire n_7181;
wire n_173;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_2136;
wire n_433;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_253;
wire n_928;
wire n_3769;
wire n_7825;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_128;
wire n_7916;
wire n_3055;
wire n_420;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_748;
wire n_7903;
wire n_7089;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_7604;
wire n_7647;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_330;
wire n_5868;
wire n_6417;
wire n_328;
wire n_368;
wire n_7145;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_7803;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_5104;
wire n_6961;
wire n_576;
wire n_511;
wire n_7622;
wire n_429;
wire n_7839;
wire n_6792;
wire n_7720;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_8136;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_141;
wire n_4430;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_1356;
wire n_6831;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_312;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_7809;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_623;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_453;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_543;
wire n_6986;
wire n_3456;
wire n_4532;
wire n_236;
wire n_601;
wire n_7564;
wire n_628;
wire n_5863;
wire n_6633;
wire n_3790;
wire n_7775;
wire n_907;
wire n_7118;
wire n_7960;
wire n_6152;
wire n_5734;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_7636;
wire n_4341;
wire n_1694;
wire n_6925;
wire n_7186;
wire n_593;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_5480;
wire n_4650;
wire n_6428;
wire n_609;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_8066;
wire n_7666;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_7967;
wire n_5977;
wire n_519;
wire n_384;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_7301;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_7262;
wire n_234;
wire n_5959;
wire n_8056;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_7584;
wire n_7748;
wire n_1789;
wire n_763;
wire n_6301;
wire n_2174;
wire n_540;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_1687;
wire n_4703;
wire n_6282;
wire n_4934;
wire n_7686;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_395;
wire n_6737;
wire n_1587;
wire n_213;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_6459;
wire n_1427;
wire n_7670;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_114;
wire n_5228;
wire n_1100;
wire n_585;
wire n_1617;
wire n_2600;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_6448;
wire n_5186;
wire n_7930;
wire n_7487;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_580;
wire n_3664;
wire n_4218;
wire n_434;
wire n_4687;
wire n_7077;
wire n_394;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_5604;
wire n_3470;
wire n_243;
wire n_7663;
wire n_5221;
wire n_7024;
wire n_1407;
wire n_8148;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_7214;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_7977;
wire n_121;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_3989;
wire n_7652;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_7566;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_322;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_558;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_653;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_556;
wire n_170;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_1471;
wire n_6212;
wire n_3440;
wire n_6816;
wire n_3658;
wire n_7374;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_7678;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_7975;
wire n_6089;
wire n_591;
wire n_5634;
wire n_5133;
wire n_7553;
wire n_5990;
wire n_5305;
wire n_2175;
wire n_1625;
wire n_7086;
wire n_5689;
wire n_7732;
wire n_7891;
wire n_4578;
wire n_318;
wire n_5644;
wire n_3644;
wire n_8038;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_528;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_7038;
wire n_7994;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_8111;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_7345;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_631;
wire n_8021;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_7041;
wire n_6717;
wire n_7593;
wire n_898;
wire n_6881;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_6672;
wire n_5343;
wire n_7757;
wire n_1093;
wire n_7866;
wire n_6518;
wire n_7334;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_6242;
wire n_336;
wire n_6601;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_668;
wire n_2111;
wire n_3743;
wire n_8079;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_7758;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_291;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_7705;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_369;
wire n_240;
wire n_7333;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_8006;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_7337;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_7439;
wire n_4371;
wire n_188;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_7210;
wire n_7744;
wire n_3898;
wire n_694;
wire n_6228;
wire n_6702;
wire n_7358;
wire n_4749;
wire n_7707;
wire n_5924;
wire n_1845;
wire n_7733;
wire n_921;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_7684;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_6997;
wire n_6371;
wire n_4238;
wire n_904;
wire n_7673;
wire n_2005;
wire n_1696;
wire n_7187;
wire n_8013;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_7313;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_3203;
wire n_383;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_6264;
wire n_5782;
wire n_8119;
wire n_630;
wire n_4168;
wire n_1369;
wire n_7036;
wire n_4298;
wire n_7370;
wire n_7931;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_8044;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_235;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_7480;
wire n_371;
wire n_5185;
wire n_2964;
wire n_308;
wire n_5032;
wire n_6990;
wire n_865;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_6288;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_7380;
wire n_2839;
wire n_3237;
wire n_7708;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_6277;
wire n_5115;
wire n_7376;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_596;
wire n_6409;
wire n_4095;
wire n_1310;
wire n_5927;
wire n_4485;
wire n_7657;
wire n_6388;
wire n_574;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_6864;
wire n_1516;
wire n_4890;
wire n_8084;
wire n_2485;
wire n_6679;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_5507;
wire n_195;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_7504;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1631;
wire n_7602;
wire n_156;
wire n_6566;
wire n_1794;
wire n_5696;
wire n_7998;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_204;
wire n_7557;
wire n_3772;
wire n_7408;
wire n_2891;
wire n_496;
wire n_7026;
wire n_4335;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_7394;
wire n_263;
wire n_4516;
wire n_5235;
wire n_360;
wire n_1129;
wire n_7627;
wire n_6436;
wire n_1464;
wire n_7719;
wire n_2798;
wire n_7450;
wire n_165;
wire n_3217;
wire n_6081;
wire n_1249;
wire n_329;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_340;
wire n_3201;
wire n_7462;
wire n_7780;
wire n_3503;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_177;
wire n_364;
wire n_258;
wire n_7582;
wire n_5521;
wire n_431;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_7555;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_447;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_841;
wire n_3204;
wire n_7451;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_18),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_58),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_50),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_59),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_7),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_28),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_40),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_38),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_32),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_64),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_13),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_23),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_17),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_2),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_28),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_52),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_2),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_85),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_45),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_10),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_23),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_22),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_67),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_20),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_10),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_71),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_17),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_22),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_49),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_20),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_14),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_93),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_0),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_14),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_55),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_18),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_24),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_32),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_43),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_40),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_30),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_15),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_34),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_90),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_68),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_98),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_76),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_39),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_35),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_72),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_12),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_83),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_24),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_42),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_100),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_86),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_36),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_4),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_37),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_19),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_97),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_80),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_6),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_41),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_11),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_82),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_60),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_84),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_39),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_77),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_5),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_75),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_3),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_33),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_4),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_0),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_88),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_57),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_35),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_94),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_19),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_27),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_66),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_37),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_56),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_145),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_122),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_153),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_153),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_122),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_122),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_136),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_152),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_116),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

INVx4_ASAP7_75t_R g233 ( 
.A(n_119),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_118),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_124),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_109),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_119),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_109),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_112),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

INVxp33_ASAP7_75t_SL g243 ( 
.A(n_111),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_128),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_128),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_117),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_237),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_235),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_235),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_236),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_236),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_110),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_219),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_239),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_239),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_220),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_246),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_224),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_219),
.B(n_224),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_225),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_225),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_222),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_223),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_217),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_223),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_243),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_246),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_219),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_262),
.B(n_243),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_274),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_257),
.A2(n_245),
.B(n_247),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

AND2x6_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_160),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_250),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_276),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_253),
.A2(n_229),
.B1(n_129),
.B2(n_189),
.Y(n_305)
);

AND2x6_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_160),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_255),
.A2(n_229),
.B1(n_190),
.B2(n_147),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_280),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_262),
.A2(n_186),
.B1(n_206),
.B2(n_203),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_248),
.B(n_226),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_252),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_277),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_259),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_258),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_249),
.B(n_237),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_226),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_260),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_241),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_254),
.Y(n_325)
);

BUFx8_ASAP7_75t_L g326 ( 
.A(n_256),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_272),
.B(n_245),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_254),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_266),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_263),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_266),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_265),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_267),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_261),
.B(n_200),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_267),
.B(n_111),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_269),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_270),
.B(n_143),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_270),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_271),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_271),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_278),
.B(n_112),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_279),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_279),
.Y(n_346)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_250),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_273),
.B(n_143),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_249),
.B(n_113),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_253),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_281),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_257),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_285),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_249),
.B(n_113),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_257),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_248),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_285),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_273),
.B(n_159),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_257),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_285),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_274),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_257),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_274),
.Y(n_367)
);

NOR2x1_ASAP7_75t_L g368 ( 
.A(n_275),
.B(n_126),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_257),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_281),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_285),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_281),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_285),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_273),
.B(n_227),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_281),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_285),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_285),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_274),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_285),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_257),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_249),
.B(n_114),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_249),
.B(n_114),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_273),
.B(n_227),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_257),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_275),
.B(n_127),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_262),
.A2(n_121),
.B1(n_120),
.B2(n_215),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_272),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_250),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_253),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_285),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_274),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_257),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_285),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_249),
.B(n_115),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_249),
.B(n_115),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_285),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_R g397 ( 
.A(n_259),
.B(n_123),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_257),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_257),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_295),
.B(n_123),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_295),
.B(n_184),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_295),
.B(n_184),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_307),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_307),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_286),
.B(n_228),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_290),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_291),
.Y(n_407)
);

AND3x2_ASAP7_75t_L g408 ( 
.A(n_317),
.B(n_137),
.C(n_130),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_291),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_316),
.Y(n_410)
);

CKINVDCx6p67_ASAP7_75t_R g411 ( 
.A(n_333),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_290),
.Y(n_412)
);

NAND2xp33_ASAP7_75t_L g413 ( 
.A(n_368),
.B(n_397),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_300),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_291),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_309),
.B(n_120),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_286),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_300),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_316),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_325),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_289),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_294),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_325),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_352),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

BUFx6f_ASAP7_75t_SL g427 ( 
.A(n_360),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_336),
.B(n_193),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_354),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_357),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_362),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_347),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_315),
.B(n_358),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_387),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_385),
.B(n_193),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_362),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_335),
.B(n_196),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_346),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_366),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_348),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_348),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_387),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_366),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_369),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_399),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_369),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_330),
.B(n_121),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_352),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_306),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_399),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_330),
.B(n_196),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_380),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_392),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_315),
.B(n_228),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_398),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_360),
.B(n_319),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_328),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_331),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_347),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_374),
.B(n_231),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_387),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_360),
.B(n_197),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_329),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_331),
.Y(n_470)
);

CKINVDCx6p67_ASAP7_75t_R g471 ( 
.A(n_320),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_331),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_314),
.B(n_185),
.C(n_186),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_331),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_319),
.B(n_197),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_331),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_347),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_337),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_334),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_334),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_338),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_341),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_334),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_288),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_306),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_334),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_334),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_297),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_355),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_323),
.B(n_198),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_342),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_359),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_322),
.B(n_198),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_342),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_305),
.B(n_185),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_322),
.B(n_202),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_287),
.B(n_203),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_324),
.B(n_204),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_361),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_363),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_342),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_342),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_323),
.B(n_202),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_324),
.B(n_296),
.Y(n_504)
);

AOI21x1_ASAP7_75t_L g505 ( 
.A1(n_327),
.A2(n_132),
.B(n_209),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_365),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_289),
.B(n_214),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_371),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_342),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_304),
.B(n_214),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_373),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_376),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_304),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_343),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_343),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_343),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_377),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_343),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_299),
.B(n_204),
.Y(n_519)
);

BUFx6f_ASAP7_75t_SL g520 ( 
.A(n_350),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_313),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_374),
.B(n_231),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_308),
.B(n_206),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_343),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_364),
.B(n_216),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_347),
.Y(n_526)
);

AOI21x1_ASAP7_75t_L g527 ( 
.A1(n_303),
.A2(n_142),
.B(n_194),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_311),
.B(n_212),
.Y(n_528)
);

INVxp33_ASAP7_75t_SL g529 ( 
.A(n_364),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_379),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_390),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_393),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_345),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_345),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_294),
.B(n_216),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_345),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_350),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_396),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_345),
.Y(n_539)
);

NAND3xp33_ASAP7_75t_L g540 ( 
.A(n_386),
.B(n_212),
.C(n_215),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_345),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_303),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_367),
.B(n_133),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_310),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_310),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_294),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_383),
.B(n_159),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_367),
.B(n_134),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_350),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_298),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_340),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_378),
.B(n_391),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_294),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_378),
.B(n_139),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_313),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_294),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_321),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_383),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_301),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_391),
.B(n_146),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_332),
.B(n_150),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_298),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_301),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_301),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_339),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_339),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_301),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_301),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_302),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_389),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_389),
.Y(n_571)
);

AO22x2_ASAP7_75t_L g572 ( 
.A1(n_339),
.A2(n_165),
.B1(n_213),
.B2(n_210),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_302),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_302),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_317),
.B(n_232),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_293),
.B(n_155),
.Y(n_576)
);

NAND3xp33_ASAP7_75t_L g577 ( 
.A(n_351),
.B(n_168),
.C(n_156),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_318),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_302),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_302),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_353),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_356),
.B(n_158),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_353),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_353),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_349),
.B(n_163),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_353),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_388),
.B(n_232),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_353),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_370),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_370),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_381),
.B(n_238),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_370),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_370),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_370),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_372),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_372),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_372),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_382),
.B(n_394),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_372),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_395),
.B(n_176),
.C(n_177),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_372),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_375),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_375),
.Y(n_603)
);

BUFx6f_ASAP7_75t_SL g604 ( 
.A(n_306),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_318),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_375),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_344),
.B(n_125),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_375),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_292),
.A2(n_131),
.B1(n_211),
.B2(n_208),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_375),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_292),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_312),
.B(n_238),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_326),
.B(n_138),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_292),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_292),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_292),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_292),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_306),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_306),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_306),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_326),
.Y(n_621)
);

BUFx10_ASAP7_75t_L g622 ( 
.A(n_326),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_295),
.B(n_140),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_298),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_307),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_295),
.B(n_141),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_307),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_352),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_291),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_286),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_295),
.B(n_151),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_290),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_L g633 ( 
.A(n_385),
.B(n_162),
.C(n_149),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_290),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_290),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_290),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_295),
.B(n_154),
.Y(n_637)
);

AND3x2_ASAP7_75t_L g638 ( 
.A(n_317),
.B(n_188),
.C(n_167),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_290),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_300),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_309),
.B(n_207),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_291),
.Y(n_642)
);

INVxp67_ASAP7_75t_R g643 ( 
.A(n_293),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_319),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_307),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_286),
.B(n_244),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_290),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_291),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_295),
.B(n_174),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_307),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_385),
.B(n_164),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_286),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_307),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_290),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_300),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_291),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_504),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_403),
.B(n_165),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_450),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_403),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_474),
.B(n_135),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_427),
.A2(n_175),
.B1(n_157),
.B2(n_161),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_450),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_414),
.Y(n_664)
);

OR2x2_ASAP7_75t_SL g665 ( 
.A(n_621),
.B(n_187),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_414),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_474),
.B(n_135),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_414),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_422),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_422),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_404),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_425),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_417),
.B(n_169),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_605),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_570),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_558),
.B(n_244),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_449),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_417),
.B(n_205),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_404),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_630),
.B(n_171),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_513),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_630),
.B(n_181),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_474),
.B(n_135),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_625),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_570),
.Y(n_685)
);

BUFx4f_ASAP7_75t_L g686 ( 
.A(n_411),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_625),
.Y(n_687)
);

BUFx8_ASAP7_75t_SL g688 ( 
.A(n_644),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_504),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_543),
.B(n_199),
.C(n_201),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_434),
.B(n_242),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_627),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_627),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_427),
.A2(n_558),
.B1(n_520),
.B2(n_549),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_571),
.Y(n_695)
);

INVx5_ASAP7_75t_L g696 ( 
.A(n_450),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_622),
.Y(n_697)
);

NAND2x1p5_ASAP7_75t_L g698 ( 
.A(n_550),
.B(n_242),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_537),
.B(n_1),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_652),
.B(n_166),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_645),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_645),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_450),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_520),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_650),
.B(n_148),
.Y(n_705)
);

BUFx10_ASAP7_75t_L g706 ( 
.A(n_554),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_437),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_652),
.B(n_170),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_598),
.B(n_3),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_462),
.B(n_5),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_474),
.B(n_135),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_466),
.B(n_522),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_529),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_437),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_650),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_653),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_571),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_653),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_463),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_437),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_463),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_440),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_622),
.Y(n_723)
);

AND2x6_ASAP7_75t_L g724 ( 
.A(n_618),
.B(n_148),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_628),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_466),
.B(n_172),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_411),
.B(n_178),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_440),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_483),
.B(n_135),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_440),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_622),
.Y(n_731)
);

CKINVDCx11_ASAP7_75t_R g732 ( 
.A(n_421),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_444),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_469),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_469),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_444),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_550),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_478),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_485),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_427),
.B(n_6),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_427),
.B(n_7),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_522),
.B(n_173),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_434),
.B(n_8),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_537),
.B(n_8),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_421),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_628),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_478),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_549),
.B(n_9),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_421),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_483),
.B(n_135),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_498),
.B(n_11),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_444),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_485),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_405),
.B(n_180),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_445),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_483),
.B(n_135),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_422),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_575),
.B(n_12),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_422),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_485),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_405),
.B(n_182),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_481),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_575),
.B(n_13),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_618),
.B(n_148),
.Y(n_764)
);

NAND2x1p5_ASAP7_75t_L g765 ( 
.A(n_550),
.B(n_148),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_445),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_646),
.B(n_183),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_481),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_621),
.B(n_15),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_422),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_483),
.B(n_516),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_482),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_445),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_482),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_646),
.B(n_16),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_516),
.B(n_148),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_436),
.B(n_16),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_520),
.Y(n_778)
);

INVx4_ASAP7_75t_L g779 ( 
.A(n_520),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_521),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_551),
.B(n_21),
.Y(n_781)
);

CKINVDCx16_ASAP7_75t_R g782 ( 
.A(n_622),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_551),
.B(n_21),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_621),
.B(n_25),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_422),
.B(n_144),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_484),
.Y(n_786)
);

AND2x6_ASAP7_75t_L g787 ( 
.A(n_618),
.B(n_611),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_484),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_565),
.B(n_25),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_556),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_468),
.B(n_26),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_447),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_578),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_498),
.B(n_26),
.Y(n_794)
);

BUFx10_ASAP7_75t_L g795 ( 
.A(n_576),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_624),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_555),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_488),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_488),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_572),
.A2(n_144),
.B1(n_233),
.B2(n_30),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_489),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_516),
.B(n_144),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_651),
.B(n_27),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_565),
.B(n_29),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_489),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_447),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_447),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_453),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_SL g809 ( 
.A(n_471),
.B(n_421),
.Y(n_809)
);

BUFx6f_ASAP7_75t_SL g810 ( 
.A(n_471),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_492),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_572),
.A2(n_144),
.B1(n_233),
.B2(n_33),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_516),
.B(n_144),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_587),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_587),
.B(n_29),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_438),
.B(n_31),
.Y(n_816)
);

NAND2x1p5_ASAP7_75t_L g817 ( 
.A(n_624),
.B(n_54),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_572),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_582),
.B(n_38),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_416),
.B(n_44),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_497),
.B(n_46),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_453),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_524),
.B(n_47),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_524),
.B(n_48),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_453),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_524),
.B(n_464),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_492),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_499),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_572),
.Y(n_829)
);

CKINVDCx11_ASAP7_75t_R g830 ( 
.A(n_643),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_624),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_499),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_500),
.Y(n_833)
);

AND2x2_ASAP7_75t_SL g834 ( 
.A(n_609),
.B(n_62),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_556),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_591),
.B(n_63),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_500),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_524),
.B(n_73),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_591),
.B(n_493),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_454),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_556),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_454),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_464),
.B(n_78),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_562),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_556),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_454),
.Y(n_846)
);

NAND3x1_ASAP7_75t_L g847 ( 
.A(n_609),
.B(n_96),
.C(n_99),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_556),
.B(n_103),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_506),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_506),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_556),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_643),
.B(n_448),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_508),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_455),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_455),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_508),
.A2(n_538),
.B1(n_532),
.B2(n_531),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_496),
.B(n_459),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_566),
.B(n_459),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_559),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_511),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_566),
.B(n_433),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_562),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_511),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_464),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_433),
.B(n_465),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_455),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_512),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_559),
.Y(n_868)
);

INVx6_ASAP7_75t_L g869 ( 
.A(n_559),
.Y(n_869)
);

OR2x2_ASAP7_75t_SL g870 ( 
.A(n_473),
.B(n_540),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_408),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_559),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_512),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_517),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_517),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_607),
.B(n_557),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_465),
.B(n_477),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_641),
.B(n_585),
.Y(n_878)
);

BUFx10_ASAP7_75t_L g879 ( 
.A(n_519),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_638),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_523),
.B(n_528),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_456),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_495),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_559),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_530),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_470),
.B(n_480),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_477),
.B(n_526),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_456),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_552),
.B(n_547),
.Y(n_889)
);

AND2x6_ASAP7_75t_L g890 ( 
.A(n_611),
.B(n_619),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_456),
.Y(n_891)
);

NAND2x1p5_ASAP7_75t_L g892 ( 
.A(n_526),
.B(n_470),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_470),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_557),
.B(n_530),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_531),
.Y(n_895)
);

OAI21xp33_ASAP7_75t_SL g896 ( 
.A1(n_532),
.A2(n_538),
.B(n_428),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_446),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_446),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_480),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_451),
.Y(n_900)
);

XOR2xp5_ASAP7_75t_L g901 ( 
.A(n_495),
.B(n_612),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_612),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_633),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_559),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_451),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_457),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_410),
.B(n_419),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_410),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_419),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_457),
.Y(n_910)
);

OR2x2_ASAP7_75t_SL g911 ( 
.A(n_577),
.B(n_600),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_561),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_613),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_457),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_593),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_593),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_SL g917 ( 
.A(n_604),
.B(n_616),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_452),
.B(n_400),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_420),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_475),
.B(n_490),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_420),
.B(n_424),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_480),
.B(n_486),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_548),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_424),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_426),
.B(n_439),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_426),
.B(n_439),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_441),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_458),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_593),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_503),
.B(n_507),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_486),
.B(n_487),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_401),
.B(n_402),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_442),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_560),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_442),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_418),
.Y(n_936)
);

AND2x2_ASAP7_75t_SL g937 ( 
.A(n_486),
.B(n_487),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_593),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_458),
.Y(n_939)
);

INVx6_ASAP7_75t_L g940 ( 
.A(n_593),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_510),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_413),
.B(n_407),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_458),
.Y(n_943)
);

NAND2xp33_ASAP7_75t_L g944 ( 
.A(n_593),
.B(n_594),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_487),
.B(n_491),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_594),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_491),
.B(n_494),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_594),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_460),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_460),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_491),
.B(n_494),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_418),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_460),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_461),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_525),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_494),
.B(n_501),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_594),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_623),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_501),
.B(n_502),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_594),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_423),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_626),
.B(n_631),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_461),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_501),
.B(n_502),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_423),
.Y(n_965)
);

AND2x6_ASAP7_75t_L g966 ( 
.A(n_611),
.B(n_619),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_461),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_429),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_637),
.B(n_649),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_407),
.B(n_409),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_502),
.B(n_509),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_509),
.Y(n_972)
);

AND2x6_ASAP7_75t_L g973 ( 
.A(n_620),
.B(n_614),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_429),
.B(n_430),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_937),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_669),
.Y(n_976)
);

OAI21xp33_ASAP7_75t_L g977 ( 
.A1(n_878),
.A2(n_535),
.B(n_407),
.Y(n_977)
);

INVx8_ASAP7_75t_L g978 ( 
.A(n_696),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_907),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_921),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_L g981 ( 
.A(n_696),
.B(n_594),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_664),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_664),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_657),
.B(n_509),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_881),
.B(n_514),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_666),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_712),
.B(n_514),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_879),
.B(n_514),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_689),
.B(n_515),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_839),
.B(n_515),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_L g991 ( 
.A(n_696),
.B(n_407),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_925),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_793),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_937),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_876),
.B(n_515),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_672),
.Y(n_996)
);

INVxp67_ASAP7_75t_L g997 ( 
.A(n_725),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_857),
.B(n_518),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_814),
.B(n_518),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_834),
.A2(n_430),
.B1(n_432),
.B2(n_655),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_696),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_746),
.B(n_518),
.Y(n_1002)
);

OAI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_727),
.A2(n_539),
.B1(n_541),
.B2(n_536),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_926),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_660),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_709),
.B(n_533),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_709),
.B(n_533),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_666),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_879),
.B(n_533),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_858),
.B(n_534),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_706),
.B(n_534),
.Y(n_1011)
);

NOR2xp67_ASAP7_75t_L g1012 ( 
.A(n_796),
.B(n_534),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_858),
.B(n_536),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_858),
.B(n_536),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_835),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_869),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_691),
.B(n_539),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_879),
.B(n_539),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_758),
.B(n_541),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_763),
.B(n_541),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_671),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_668),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_894),
.B(n_472),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_706),
.B(n_573),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_668),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_707),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_743),
.B(n_719),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_679),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_706),
.B(n_573),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_L g1030 ( 
.A(n_821),
.B(n_479),
.C(n_476),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_834),
.A2(n_640),
.B1(n_655),
.B2(n_431),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_721),
.B(n_479),
.Y(n_1032)
);

INVx8_ASAP7_75t_L g1033 ( 
.A(n_931),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_695),
.B(n_588),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_901),
.A2(n_640),
.B1(n_432),
.B2(n_431),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_795),
.B(n_472),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_717),
.B(n_595),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_677),
.B(n_595),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_707),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_734),
.B(n_476),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_797),
.B(n_601),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_735),
.B(n_656),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_SL g1043 ( 
.A(n_681),
.B(n_604),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_889),
.B(n_601),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_688),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_795),
.B(n_656),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_795),
.B(n_656),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_713),
.B(n_599),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_686),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_684),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_687),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_821),
.A2(n_588),
.B1(n_597),
.B2(n_599),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_692),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_686),
.B(n_656),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_856),
.A2(n_642),
.B1(n_409),
.B2(n_648),
.Y(n_1055)
);

AO22x2_ASAP7_75t_L g1056 ( 
.A1(n_699),
.A2(n_744),
.B1(n_784),
.B2(n_769),
.Y(n_1056)
);

OAI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_751),
.A2(n_467),
.B1(n_409),
.B2(n_648),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_713),
.B(n_597),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_714),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_829),
.A2(n_545),
.B1(n_544),
.B2(n_542),
.Y(n_1060)
);

OAI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_815),
.A2(n_467),
.B1(n_409),
.B2(n_648),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_697),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_704),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_852),
.B(n_467),
.Y(n_1064)
);

AND2x6_ASAP7_75t_SL g1065 ( 
.A(n_688),
.B(n_617),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_681),
.B(n_467),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_720),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_738),
.B(n_629),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_710),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_747),
.B(n_629),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_720),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_675),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_693),
.Y(n_1073)
);

OAI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_690),
.A2(n_642),
.B1(n_648),
.B2(n_415),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_762),
.B(n_768),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_745),
.B(n_749),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_869),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_745),
.B(n_443),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_780),
.B(n_603),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_869),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_722),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_772),
.B(n_443),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_749),
.B(n_443),
.Y(n_1083)
);

BUFx5_ASAP7_75t_L g1084 ( 
.A(n_787),
.Y(n_1084)
);

NOR2xp67_ASAP7_75t_SL g1085 ( 
.A(n_669),
.B(n_642),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_774),
.B(n_443),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_722),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_701),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_728),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_702),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_710),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_786),
.B(n_642),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_674),
.B(n_629),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_728),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_941),
.B(n_629),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_715),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_730),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_730),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_733),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_788),
.B(n_415),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_798),
.B(n_799),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_716),
.Y(n_1102)
);

O2A1O1Ixp5_ASAP7_75t_L g1103 ( 
.A1(n_819),
.A2(n_584),
.B(n_596),
.C(n_602),
.Y(n_1103)
);

OAI221xp5_ASAP7_75t_L g1104 ( 
.A1(n_791),
.A2(n_415),
.B1(n_435),
.B2(n_617),
.C(n_615),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_941),
.B(n_415),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_801),
.B(n_805),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_819),
.A2(n_603),
.B1(n_615),
.B2(n_614),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_718),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_733),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_811),
.B(n_435),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_809),
.B(n_435),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_934),
.B(n_435),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_816),
.A2(n_820),
.B(n_791),
.C(n_783),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_736),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_934),
.B(n_584),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_789),
.B(n_584),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_897),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_898),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_940),
.Y(n_1119)
);

INVxp67_ASAP7_75t_L g1120 ( 
.A(n_685),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_789),
.B(n_804),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_736),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_900),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_827),
.B(n_828),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_781),
.Y(n_1125)
);

INVxp33_ASAP7_75t_L g1126 ( 
.A(n_830),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_832),
.B(n_545),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_905),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_833),
.B(n_544),
.Y(n_1129)
);

OAI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_803),
.A2(n_580),
.B1(n_592),
.B2(n_610),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_789),
.B(n_584),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_816),
.A2(n_592),
.B(n_606),
.C(n_610),
.Y(n_1132)
);

NOR3xp33_ASAP7_75t_L g1133 ( 
.A(n_932),
.B(n_918),
.C(n_958),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_804),
.B(n_602),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_804),
.B(n_602),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_918),
.A2(n_592),
.B1(n_606),
.B2(n_610),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_913),
.B(n_581),
.Y(n_1137)
);

NAND2xp33_ASAP7_75t_L g1138 ( 
.A(n_669),
.B(n_581),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_752),
.Y(n_1139)
);

BUFx4_ASAP7_75t_L g1140 ( 
.A(n_810),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_752),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_837),
.B(n_545),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_849),
.B(n_544),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_850),
.B(n_542),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_781),
.A2(n_580),
.B1(n_579),
.B2(n_608),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_853),
.B(n_860),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_932),
.B(n_606),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_863),
.B(n_542),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_867),
.B(n_546),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_912),
.B(n_580),
.Y(n_1150)
);

NAND2xp33_ASAP7_75t_L g1151 ( 
.A(n_669),
.B(n_602),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_873),
.B(n_581),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_913),
.B(n_581),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_755),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_SL g1155 ( 
.A(n_670),
.B(n_757),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_908),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_874),
.B(n_875),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_SL g1158 ( 
.A(n_697),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_955),
.B(n_596),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_704),
.B(n_620),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_755),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_885),
.B(n_596),
.Y(n_1162)
);

NOR2xp67_ASAP7_75t_L g1163 ( 
.A(n_796),
.B(n_596),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_766),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_766),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_835),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_909),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_903),
.B(n_579),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_895),
.B(n_579),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_676),
.B(n_574),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_940),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_919),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_676),
.B(n_783),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_773),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_676),
.B(n_574),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_794),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_769),
.B(n_574),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_769),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_970),
.A2(n_546),
.B(n_608),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_673),
.B(n_546),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_670),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_673),
.B(n_680),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_835),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_680),
.B(n_608),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_682),
.B(n_586),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_784),
.B(n_586),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_784),
.B(n_583),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_740),
.A2(n_583),
.B1(n_569),
.B2(n_590),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_682),
.B(n_589),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_726),
.B(n_589),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_938),
.Y(n_1191)
);

INVxp33_ASAP7_75t_L g1192 ( 
.A(n_830),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_773),
.Y(n_1193)
);

AND2x2_ASAP7_75t_SL g1194 ( 
.A(n_800),
.B(n_569),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_944),
.A2(n_590),
.B(n_568),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_923),
.B(n_865),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_777),
.A2(n_568),
.B(n_567),
.C(n_564),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_792),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_865),
.B(n_567),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_865),
.B(n_563),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_792),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_877),
.B(n_563),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_806),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_SL g1204 ( 
.A(n_818),
.B(n_564),
.C(n_553),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_806),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_807),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_924),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_723),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_920),
.B(n_930),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_775),
.B(n_553),
.Y(n_1210)
);

BUFx8_ASAP7_75t_L g1211 ( 
.A(n_810),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_807),
.Y(n_1212)
);

NAND2x1_ASAP7_75t_L g1213 ( 
.A(n_940),
.B(n_406),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_742),
.B(n_406),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_754),
.B(n_406),
.Y(n_1215)
);

INVxp67_ASAP7_75t_SL g1216 ( 
.A(n_944),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_808),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_808),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_822),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_761),
.B(n_767),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_699),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_740),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_870),
.B(n_505),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_741),
.A2(n_604),
.B1(n_634),
.B2(n_635),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_927),
.B(n_654),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_933),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_822),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_748),
.B(n_654),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_962),
.B(n_505),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_704),
.B(n_412),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_969),
.B(n_604),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_877),
.B(n_412),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_935),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_748),
.B(n_654),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_877),
.B(n_412),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_678),
.B(n_647),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_974),
.Y(n_1237)
);

OAI221xp5_ASAP7_75t_L g1238 ( 
.A1(n_812),
.A2(n_741),
.B1(n_880),
.B2(n_871),
.C(n_896),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_902),
.A2(n_632),
.B1(n_634),
.B2(n_635),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_861),
.B(n_647),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_861),
.B(n_647),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_887),
.B(n_796),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_861),
.B(n_632),
.Y(n_1243)
);

INVxp67_ASAP7_75t_L g1244 ( 
.A(n_883),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_825),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_699),
.B(n_632),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_744),
.B(n_639),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_942),
.B(n_665),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_968),
.Y(n_1249)
);

O2A1O1Ixp5_ASAP7_75t_L g1250 ( 
.A1(n_661),
.A2(n_634),
.B(n_635),
.C(n_636),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_825),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_902),
.A2(n_636),
.B1(n_639),
.B2(n_527),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_968),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_744),
.B(n_636),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_887),
.B(n_639),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_887),
.B(n_527),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_670),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_945),
.B(n_956),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_936),
.Y(n_1259)
);

NAND2xp33_ASAP7_75t_L g1260 ( 
.A(n_670),
.B(n_757),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_840),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_945),
.B(n_956),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_945),
.B(n_956),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_844),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_778),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_840),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_757),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_842),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_842),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_959),
.B(n_964),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_959),
.B(n_964),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_959),
.B(n_964),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_658),
.A2(n_662),
.B1(n_931),
.B2(n_844),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_732),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_864),
.B(n_893),
.Y(n_1275)
);

AND2x6_ASAP7_75t_L g1276 ( 
.A(n_659),
.B(n_663),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_782),
.B(n_732),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_911),
.B(n_723),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_700),
.A2(n_708),
.B(n_771),
.C(n_826),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_731),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_864),
.B(n_893),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_778),
.B(n_779),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_931),
.B(n_694),
.Y(n_1283)
);

INVxp33_ASAP7_75t_L g1284 ( 
.A(n_698),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_831),
.B(n_737),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_846),
.Y(n_1286)
);

INVx4_ASAP7_75t_L g1287 ( 
.A(n_778),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_846),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_952),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_899),
.B(n_972),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_938),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_862),
.A2(n_779),
.B1(n_965),
.B2(n_961),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_854),
.Y(n_1293)
);

INVxp67_ASAP7_75t_L g1294 ( 
.A(n_862),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_899),
.B(n_972),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_731),
.B(n_771),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_854),
.B(n_855),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_855),
.B(n_866),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_826),
.B(n_836),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_866),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_882),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_882),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_888),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_888),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_891),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_886),
.B(n_922),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_970),
.A2(n_957),
.B(n_659),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_886),
.B(n_922),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_891),
.B(n_906),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_931),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_658),
.A2(n_847),
.B1(n_698),
.B2(n_848),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_779),
.B(n_831),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_957),
.A2(n_760),
.B(n_659),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_906),
.B(n_910),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_831),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_910),
.B(n_914),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_947),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_737),
.B(n_757),
.Y(n_1318)
);

OR2x6_ASAP7_75t_L g1319 ( 
.A(n_663),
.B(n_703),
.Y(n_1319)
);

OAI221xp5_ASAP7_75t_L g1320 ( 
.A1(n_951),
.A2(n_971),
.B1(n_848),
.B2(n_892),
.C(n_947),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_914),
.B(n_954),
.Y(n_1321)
);

AND2x4_ASAP7_75t_SL g1322 ( 
.A(n_938),
.B(n_904),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_663),
.A2(n_753),
.B1(n_760),
.B2(n_739),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_928),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_939),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_951),
.B(n_971),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_943),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_943),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_949),
.B(n_967),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_892),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_658),
.Y(n_1331)
);

BUFx8_ASAP7_75t_L g1332 ( 
.A(n_658),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_759),
.B(n_851),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_949),
.B(n_967),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_658),
.A2(n_963),
.B1(n_954),
.B2(n_953),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_950),
.B(n_963),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_950),
.B(n_845),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_973),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_841),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_973),
.A2(n_966),
.B1(n_890),
.B2(n_787),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_759),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_703),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_759),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_973),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_759),
.Y(n_1345)
);

OR2x6_ASAP7_75t_L g1346 ( 
.A(n_703),
.B(n_760),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_841),
.B(n_845),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_739),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_841),
.B(n_872),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_973),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_845),
.B(n_859),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_770),
.B(n_851),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_859),
.B(n_872),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_859),
.B(n_872),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_770),
.B(n_915),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_884),
.B(n_929),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_884),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_770),
.B(n_915),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_884),
.B(n_929),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_929),
.B(n_946),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_973),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_946),
.B(n_851),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_770),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_890),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_790),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_790),
.B(n_851),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_SL g1367 ( 
.A(n_705),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_890),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_790),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_787),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_787),
.A2(n_966),
.B1(n_890),
.B2(n_847),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_966),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_868),
.B(n_904),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_966),
.Y(n_1374)
);

INVx5_ASAP7_75t_L g1375 ( 
.A(n_868),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_868),
.B(n_904),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_868),
.B(n_904),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_966),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_960),
.B(n_948),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_915),
.B(n_960),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_915),
.B(n_960),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_916),
.B(n_960),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_916),
.B(n_948),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_916),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_948),
.B(n_917),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_948),
.B(n_661),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_776),
.A2(n_813),
.B1(n_802),
.B2(n_785),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_765),
.B(n_724),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_667),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_765),
.B(n_724),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_724),
.B(n_764),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_817),
.B(n_838),
.Y(n_1392)
);

NAND2xp33_ASAP7_75t_L g1393 ( 
.A(n_817),
.B(n_838),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_667),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_823),
.A2(n_824),
.B(n_813),
.C(n_802),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_724),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_683),
.B(n_756),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_724),
.B(n_764),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_683),
.A2(n_756),
.B1(n_711),
.B2(n_729),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_823),
.B(n_843),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_764),
.B(n_785),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_764),
.B(n_776),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_711),
.B(n_729),
.C(n_750),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_750),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_764),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_843),
.B(n_705),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_705),
.B(n_448),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_705),
.A2(n_878),
.B1(n_323),
.B2(n_319),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_705),
.B(n_878),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_664),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_878),
.B(n_881),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_878),
.B(n_881),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_878),
.B(n_330),
.Y(n_1413)
);

OAI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_878),
.A2(n_448),
.B1(n_324),
.B2(n_504),
.C(n_881),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_878),
.A2(n_323),
.B1(n_319),
.B2(n_834),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_664),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_878),
.B(n_881),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_978),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1056),
.B(n_1033),
.Y(n_1419)
);

NAND2x1p5_ASAP7_75t_L g1420 ( 
.A(n_1375),
.B(n_1230),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1415),
.A2(n_1414),
.B1(n_1182),
.B2(n_1113),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1225),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1225),
.Y(n_1423)
);

OR2x6_ASAP7_75t_L g1424 ( 
.A(n_1056),
.B(n_1033),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1301),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_993),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1408),
.B(n_1222),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_982),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1125),
.B(n_1069),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1417),
.B(n_1413),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1315),
.Y(n_1432)
);

NOR2xp67_ASAP7_75t_L g1433 ( 
.A(n_1375),
.B(n_1365),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1091),
.B(n_1244),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1044),
.B(n_1124),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1301),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1124),
.B(n_1209),
.Y(n_1437)
);

AND2x6_ASAP7_75t_SL g1438 ( 
.A(n_1277),
.B(n_1278),
.Y(n_1438)
);

NOR2xp67_ASAP7_75t_L g1439 ( 
.A(n_1375),
.B(n_1365),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_997),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_982),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1057),
.A2(n_1061),
.B1(n_1176),
.B2(n_1220),
.C(n_1074),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1033),
.Y(n_1443)
);

INVx6_ASAP7_75t_L g1444 ( 
.A(n_1033),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_978),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1002),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1303),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1173),
.B(n_1248),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1041),
.B(n_1133),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1315),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1056),
.B(n_1149),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1375),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1303),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1048),
.B(n_1058),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_984),
.B(n_979),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1002),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1056),
.A2(n_1121),
.B1(n_1027),
.B2(n_1052),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1304),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_989),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_979),
.B(n_980),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1375),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_978),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_991),
.A2(n_1216),
.B(n_1393),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_983),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_980),
.B(n_992),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_978),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_992),
.B(n_1004),
.Y(n_1469)
);

AND2x6_ASAP7_75t_L g1470 ( 
.A(n_1371),
.B(n_1311),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1001),
.Y(n_1471)
);

INVx5_ASAP7_75t_L g1472 ( 
.A(n_1396),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1004),
.B(n_1147),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1120),
.B(n_1072),
.Y(n_1474)
);

BUFx8_ASAP7_75t_L g1475 ( 
.A(n_1158),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1001),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1049),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_976),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1238),
.A2(n_1035),
.B1(n_1283),
.B2(n_1221),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_985),
.B(n_989),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_996),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1168),
.A2(n_1043),
.B1(n_1194),
.B2(n_1178),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_SL g1483 ( 
.A1(n_1085),
.A2(n_1223),
.B(n_1299),
.C(n_1347),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1264),
.B(n_1294),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1049),
.Y(n_1485)
);

BUFx4f_ASAP7_75t_L g1486 ( 
.A(n_1396),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1038),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1024),
.B(n_1029),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1075),
.B(n_1101),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_986),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1126),
.A2(n_1192),
.B1(n_1274),
.B2(n_1045),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1062),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1106),
.B(n_1146),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1079),
.B(n_1076),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1001),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1011),
.B(n_1273),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1157),
.B(n_1150),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1373),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1324),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_976),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_986),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1005),
.B(n_1021),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1005),
.B(n_1021),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1324),
.Y(n_1504)
);

AND2x6_ASAP7_75t_L g1505 ( 
.A(n_1311),
.B(n_1396),
.Y(n_1505)
);

OR2x6_ASAP7_75t_L g1506 ( 
.A(n_1283),
.B(n_1177),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1095),
.B(n_1105),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1332),
.A2(n_1194),
.B1(n_1231),
.B2(n_1367),
.Y(n_1508)
);

BUFx8_ASAP7_75t_L g1509 ( 
.A(n_1158),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_976),
.Y(n_1510)
);

NOR3xp33_ASAP7_75t_L g1511 ( 
.A(n_1112),
.B(n_1153),
.C(n_1137),
.Y(n_1511)
);

AND2x2_ASAP7_75t_SL g1512 ( 
.A(n_1393),
.B(n_1224),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1062),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1249),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1008),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_991),
.A2(n_981),
.B(n_1228),
.Y(n_1516)
);

A2O1A1Ixp33_ASAP7_75t_L g1517 ( 
.A1(n_1229),
.A2(n_1279),
.B(n_977),
.C(n_1030),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1249),
.Y(n_1518)
);

A2O1A1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1180),
.A2(n_1184),
.B(n_1189),
.C(n_1185),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1028),
.B(n_1050),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1022),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_981),
.A2(n_1234),
.B(n_1400),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1230),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1103),
.A2(n_1007),
.B(n_1006),
.Y(n_1525)
);

NAND2x1_ASAP7_75t_L g1526 ( 
.A(n_1155),
.B(n_1276),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1022),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1253),
.Y(n_1528)
);

NOR2x1p5_ASAP7_75t_L g1529 ( 
.A(n_1280),
.B(n_1208),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1025),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1253),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1259),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_976),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1034),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_976),
.Y(n_1535)
);

INVx5_ASAP7_75t_L g1536 ( 
.A(n_1396),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1208),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1025),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1356),
.B(n_1063),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1028),
.B(n_1050),
.Y(n_1540)
);

NOR2x1_ASAP7_75t_L g1541 ( 
.A(n_1063),
.B(n_1287),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1149),
.B(n_1129),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1409),
.B(n_1280),
.Y(n_1543)
);

INVx5_ASAP7_75t_L g1544 ( 
.A(n_1396),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1026),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1126),
.A2(n_1192),
.B1(n_1045),
.B2(n_1239),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1037),
.A2(n_1104),
.B1(n_1053),
.B2(n_1073),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1259),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1332),
.A2(n_1367),
.B1(n_975),
.B2(n_994),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1051),
.B(n_1073),
.Y(n_1550)
);

INVx4_ASAP7_75t_L g1551 ( 
.A(n_1276),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1356),
.B(n_1063),
.Y(n_1552)
);

AND2x2_ASAP7_75t_SL g1553 ( 
.A(n_1405),
.B(n_1340),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1129),
.B(n_1143),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1026),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1332),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1211),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1289),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1003),
.B(n_1356),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1039),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_975),
.A2(n_994),
.B1(n_1237),
.B2(n_1289),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1284),
.B(n_1296),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1416),
.Y(n_1563)
);

NAND2x2_ASAP7_75t_L g1564 ( 
.A(n_1343),
.B(n_1363),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1088),
.A2(n_1090),
.B1(n_1102),
.B2(n_1096),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1416),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1088),
.B(n_1090),
.Y(n_1567)
);

INVxp67_ASAP7_75t_SL g1568 ( 
.A(n_1246),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1284),
.B(n_1170),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1410),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1196),
.B(n_1064),
.Y(n_1571)
);

NOR2x1p5_ASAP7_75t_L g1572 ( 
.A(n_1287),
.B(n_1010),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1039),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1175),
.B(n_1017),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1013),
.B(n_1014),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1258),
.B(n_1262),
.Y(n_1576)
);

INVx6_ASAP7_75t_L g1577 ( 
.A(n_1287),
.Y(n_1577)
);

INVx5_ASAP7_75t_L g1578 ( 
.A(n_1405),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1373),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1116),
.A2(n_1134),
.B1(n_1135),
.B2(n_1131),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1322),
.B(n_1160),
.Y(n_1581)
);

INVx5_ASAP7_75t_L g1582 ( 
.A(n_1405),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1204),
.A2(n_1031),
.B1(n_1000),
.B2(n_1407),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1276),
.Y(n_1584)
);

NOR2x2_ASAP7_75t_L g1585 ( 
.A(n_1140),
.B(n_1065),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1181),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1096),
.B(n_1102),
.Y(n_1587)
);

AND2x6_ASAP7_75t_L g1588 ( 
.A(n_1405),
.B(n_1370),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1143),
.B(n_1237),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1322),
.B(n_1160),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_987),
.B(n_995),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_990),
.B(n_1181),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1059),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1186),
.A2(n_1187),
.B1(n_1270),
.B2(n_1263),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1271),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1059),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1108),
.A2(n_1118),
.B1(n_1123),
.B2(n_1117),
.Y(n_1597)
);

AO22x1_ASAP7_75t_L g1598 ( 
.A1(n_1405),
.A2(n_1265),
.B1(n_1310),
.B2(n_1331),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1181),
.B(n_1267),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1181),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1067),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1267),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1267),
.B(n_1345),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1108),
.A2(n_1118),
.B1(n_1123),
.B2(n_1117),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_998),
.B(n_1272),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1019),
.A2(n_1020),
.B1(n_1128),
.B2(n_1156),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1071),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1071),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1128),
.B(n_1156),
.Y(n_1609)
);

NOR2x2_ASAP7_75t_L g1610 ( 
.A(n_1140),
.B(n_1211),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1247),
.B(n_1254),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1267),
.B(n_1345),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1240),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1345),
.B(n_1369),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1343),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1241),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1345),
.B(n_1369),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1167),
.B(n_1172),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1345),
.B(n_1369),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1081),
.Y(n_1620)
);

NAND3xp33_ASAP7_75t_SL g1621 ( 
.A(n_1115),
.B(n_1066),
.C(n_1093),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1081),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1087),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1160),
.B(n_1363),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1369),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1087),
.Y(n_1626)
);

BUFx12f_ASAP7_75t_SL g1627 ( 
.A(n_1319),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1159),
.B(n_999),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1158),
.B(n_1207),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1243),
.Y(n_1630)
);

INVx3_ASAP7_75t_L g1631 ( 
.A(n_1369),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1226),
.A2(n_1233),
.B1(n_1111),
.B2(n_1107),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1188),
.B(n_1292),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1233),
.B(n_1353),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1089),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1089),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1023),
.B(n_1353),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1306),
.A2(n_1308),
.B1(n_1326),
.B2(n_1242),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1094),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1330),
.B(n_1169),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1160),
.B(n_1265),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1046),
.B(n_1047),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1379),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1379),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1190),
.A2(n_1060),
.B1(n_1261),
.B2(n_1325),
.Y(n_1645)
);

NAND3xp33_ASAP7_75t_SL g1646 ( 
.A(n_1054),
.B(n_1083),
.C(n_1078),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1382),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_1319),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1032),
.B(n_1040),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1097),
.A2(n_1302),
.B1(n_1300),
.B2(n_1293),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1097),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1382),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1275),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1136),
.B(n_1281),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1098),
.B(n_1099),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1109),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1109),
.B(n_1114),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_SL g1658 ( 
.A(n_1395),
.B(n_1036),
.C(n_1145),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1015),
.B(n_1166),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1114),
.Y(n_1660)
);

NAND2x1p5_ASAP7_75t_L g1661 ( 
.A(n_1155),
.B(n_1015),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1122),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1290),
.B(n_1295),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1211),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1055),
.A2(n_1200),
.B1(n_1199),
.B2(n_1202),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1015),
.B(n_1166),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1139),
.A2(n_1293),
.B1(n_1305),
.B2(n_1302),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1016),
.B(n_1077),
.Y(n_1668)
);

AND2x4_ASAP7_75t_SL g1669 ( 
.A(n_1319),
.B(n_1346),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1141),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1339),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1141),
.Y(n_1672)
);

INVx4_ASAP7_75t_L g1673 ( 
.A(n_1276),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1154),
.A2(n_1198),
.B1(n_1218),
.B2(n_1305),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1255),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1317),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1154),
.Y(n_1677)
);

NAND2x1p5_ASAP7_75t_L g1678 ( 
.A(n_1166),
.B(n_1183),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1339),
.Y(n_1679)
);

AND2x2_ASAP7_75t_SL g1680 ( 
.A(n_1260),
.B(n_1406),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1357),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_988),
.B(n_1009),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1404),
.A2(n_1397),
.B1(n_1086),
.B2(n_1092),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1084),
.Y(n_1684)
);

OR2x6_ASAP7_75t_L g1685 ( 
.A(n_1370),
.B(n_1378),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1161),
.A2(n_1206),
.B1(n_1325),
.B2(n_1327),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1357),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1161),
.B(n_1164),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1384),
.Y(n_1689)
);

NOR2x1p5_ASAP7_75t_L g1690 ( 
.A(n_1183),
.B(n_1191),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1165),
.B(n_1174),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1183),
.B(n_1191),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1236),
.A2(n_1210),
.B1(n_1214),
.B2(n_1215),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1193),
.B(n_1198),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1201),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1201),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1203),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1016),
.B(n_1077),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1392),
.A2(n_1403),
.B(n_1252),
.C(n_1386),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1203),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1080),
.B(n_1119),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1205),
.B(n_1206),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1191),
.B(n_1291),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1205),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1212),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1212),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1217),
.B(n_1218),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1080),
.B(n_1119),
.Y(n_1708)
);

NAND2x1p5_ASAP7_75t_L g1709 ( 
.A(n_1291),
.B(n_1378),
.Y(n_1709)
);

O2A1O1Ixp5_ASAP7_75t_L g1710 ( 
.A1(n_1213),
.A2(n_1130),
.B(n_1018),
.C(n_1132),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1384),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1127),
.B(n_1142),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1217),
.A2(n_1245),
.B1(n_1327),
.B2(n_1328),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1291),
.B(n_1163),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1219),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1219),
.B(n_1227),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1227),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_SL g1718 ( 
.A1(n_1367),
.A2(n_1084),
.B1(n_1406),
.B2(n_1344),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1144),
.B(n_1148),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1245),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1362),
.B(n_1171),
.Y(n_1721)
);

OR2x6_ASAP7_75t_L g1722 ( 
.A(n_1338),
.B(n_1344),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1349),
.B(n_1351),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1084),
.Y(n_1724)
);

INVx5_ASAP7_75t_L g1725 ( 
.A(n_1276),
.Y(n_1725)
);

AND2x6_ASAP7_75t_SL g1726 ( 
.A(n_1152),
.B(n_1162),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1276),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1383),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1354),
.B(n_1359),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1257),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1251),
.B(n_1261),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1251),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1266),
.B(n_1268),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1266),
.Y(n_1734)
);

INVx2_ASAP7_75t_SL g1735 ( 
.A(n_1321),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1268),
.Y(n_1736)
);

BUFx12f_ASAP7_75t_L g1737 ( 
.A(n_1210),
.Y(n_1737)
);

AND2x2_ASAP7_75t_SL g1738 ( 
.A(n_1138),
.B(n_1151),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1269),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1269),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1286),
.B(n_1288),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1300),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1163),
.B(n_1342),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1328),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1319),
.Y(n_1745)
);

BUFx8_ASAP7_75t_L g1746 ( 
.A(n_1084),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1321),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1297),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1042),
.B(n_1068),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1250),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1070),
.A2(n_1110),
.B1(n_1082),
.B2(n_1100),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1298),
.Y(n_1752)
);

BUFx6f_ASAP7_75t_L g1753 ( 
.A(n_1346),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1389),
.A2(n_1394),
.B1(n_1335),
.B2(n_1350),
.Y(n_1754)
);

NOR2x1p5_ASAP7_75t_L g1755 ( 
.A(n_1341),
.B(n_1368),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1309),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1342),
.B(n_1348),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1179),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1314),
.B(n_1329),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1316),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_SL g1761 ( 
.A(n_1346),
.Y(n_1761)
);

INVx5_ASAP7_75t_L g1762 ( 
.A(n_1346),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1360),
.B(n_1348),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1334),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1342),
.B(n_1348),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1336),
.B(n_1337),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1385),
.B(n_1085),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1389),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1394),
.B(n_1012),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1364),
.Y(n_1770)
);

NAND2x1p5_ASAP7_75t_L g1771 ( 
.A(n_1364),
.B(n_1374),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1318),
.B(n_1372),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1012),
.B(n_1372),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1368),
.B(n_1374),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1232),
.Y(n_1775)
);

BUFx8_ASAP7_75t_L g1776 ( 
.A(n_1084),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1235),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1338),
.B(n_1361),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1256),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1350),
.B(n_1361),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1402),
.Y(n_1781)
);

BUFx8_ASAP7_75t_L g1782 ( 
.A(n_1320),
.Y(n_1782)
);

AND2x4_ASAP7_75t_SL g1783 ( 
.A(n_1387),
.B(n_1213),
.Y(n_1783)
);

INVx4_ASAP7_75t_L g1784 ( 
.A(n_1323),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1333),
.B(n_1376),
.Y(n_1785)
);

BUFx8_ASAP7_75t_L g1786 ( 
.A(n_1352),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1399),
.A2(n_1398),
.B1(n_1391),
.B2(n_1401),
.Y(n_1787)
);

NOR2xp67_ASAP7_75t_L g1788 ( 
.A(n_1355),
.B(n_1366),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1307),
.B(n_1313),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1358),
.B(n_1380),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1377),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1381),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1285),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1388),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1197),
.Y(n_1795)
);

BUFx6f_ASAP7_75t_L g1796 ( 
.A(n_1390),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1195),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1413),
.B(n_330),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1225),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1415),
.A2(n_834),
.B1(n_878),
.B2(n_881),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1225),
.Y(n_1801)
);

INVxp67_ASAP7_75t_SL g1802 ( 
.A(n_1056),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1413),
.B(n_330),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1414),
.A2(n_305),
.B1(n_312),
.B2(n_901),
.Y(n_1804)
);

INVx2_ASAP7_75t_SL g1805 ( 
.A(n_1033),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1225),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1113),
.A2(n_1182),
.B1(n_1415),
.B2(n_834),
.Y(n_1808)
);

NAND3xp33_ASAP7_75t_SL g1809 ( 
.A(n_1415),
.B(n_323),
.C(n_319),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_993),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_978),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1225),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1225),
.Y(n_1813)
);

INVx5_ASAP7_75t_L g1814 ( 
.A(n_978),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1225),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_993),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1225),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_979),
.B(n_980),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1819)
);

BUFx6f_ASAP7_75t_L g1820 ( 
.A(n_978),
.Y(n_1820)
);

NOR3xp33_ASAP7_75t_SL g1821 ( 
.A(n_1045),
.B(n_644),
.C(n_513),
.Y(n_1821)
);

OR2x4_ASAP7_75t_L g1822 ( 
.A(n_1277),
.B(n_1024),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_1211),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1045),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1225),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1056),
.B(n_1124),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_SL g1828 ( 
.A1(n_1414),
.A2(n_1415),
.B1(n_1125),
.B2(n_1069),
.Y(n_1828)
);

INVxp67_ASAP7_75t_SL g1829 ( 
.A(n_1056),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1225),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1833)
);

OR2x6_ASAP7_75t_L g1834 ( 
.A(n_1056),
.B(n_1033),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1033),
.Y(n_1835)
);

INVx2_ASAP7_75t_SL g1836 ( 
.A(n_1033),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1225),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1173),
.B(n_1182),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1033),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1225),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1033),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_978),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1225),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_993),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1225),
.Y(n_1851)
);

BUFx8_ASAP7_75t_L g1852 ( 
.A(n_1158),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1413),
.B(n_330),
.Y(n_1853)
);

BUFx4f_ASAP7_75t_L g1854 ( 
.A(n_978),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1033),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1225),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1225),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1414),
.A2(n_305),
.B1(n_312),
.B2(n_901),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1315),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_993),
.Y(n_1860)
);

NAND3xp33_ASAP7_75t_SL g1861 ( 
.A(n_1415),
.B(n_323),
.C(n_319),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1862)
);

AOI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1415),
.A2(n_834),
.B1(n_878),
.B2(n_881),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1225),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1225),
.Y(n_1865)
);

NOR2xp67_ASAP7_75t_L g1866 ( 
.A(n_1375),
.B(n_1365),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1225),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1415),
.A2(n_834),
.B1(n_878),
.B2(n_881),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1225),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1225),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1415),
.A2(n_834),
.B1(n_878),
.B2(n_881),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1315),
.Y(n_1874)
);

NAND2x1p5_ASAP7_75t_L g1875 ( 
.A(n_1375),
.B(n_696),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1056),
.B(n_1124),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1225),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_SL g1879 ( 
.A1(n_1414),
.A2(n_1415),
.B1(n_1125),
.B2(n_1069),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_993),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1225),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1413),
.B(n_330),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1056),
.B(n_1124),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1415),
.A2(n_834),
.B1(n_878),
.B2(n_881),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1225),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1225),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1889)
);

NOR2xp67_ASAP7_75t_L g1890 ( 
.A(n_1375),
.B(n_1365),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1225),
.Y(n_1891)
);

INVx1_ASAP7_75t_SL g1892 ( 
.A(n_1002),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1225),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1225),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_L g1898 ( 
.A(n_978),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_979),
.B(n_980),
.Y(n_1899)
);

INVx2_ASAP7_75t_SL g1900 ( 
.A(n_1033),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1225),
.Y(n_1901)
);

INVx5_ASAP7_75t_L g1902 ( 
.A(n_978),
.Y(n_1902)
);

OR2x2_ASAP7_75t_SL g1903 ( 
.A(n_1182),
.B(n_782),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1225),
.Y(n_1904)
);

INVx2_ASAP7_75t_SL g1905 ( 
.A(n_1033),
.Y(n_1905)
);

BUFx4f_ASAP7_75t_L g1906 ( 
.A(n_978),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_979),
.B(n_980),
.Y(n_1907)
);

OR2x6_ASAP7_75t_L g1908 ( 
.A(n_1056),
.B(n_1033),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_978),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1912)
);

INVxp67_ASAP7_75t_SL g1913 ( 
.A(n_1056),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1414),
.A2(n_305),
.B1(n_312),
.B2(n_901),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1415),
.A2(n_834),
.B1(n_878),
.B2(n_881),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1225),
.Y(n_1919)
);

OAI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1113),
.A2(n_1182),
.B1(n_1415),
.B2(n_834),
.Y(n_1920)
);

INVx3_ASAP7_75t_L g1921 ( 
.A(n_978),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1413),
.B(n_330),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1225),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1414),
.A2(n_305),
.B1(n_312),
.B2(n_901),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1225),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1225),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1113),
.A2(n_709),
.B(n_821),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1413),
.B(n_330),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1414),
.A2(n_305),
.B1(n_312),
.B2(n_901),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1225),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_R g1936 ( 
.A(n_1045),
.B(n_681),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_978),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_978),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1225),
.Y(n_1943)
);

INVx2_ASAP7_75t_SL g1944 ( 
.A(n_1033),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1225),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1225),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1225),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1225),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1045),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1282),
.B(n_1312),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_993),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1225),
.Y(n_1953)
);

INVx4_ASAP7_75t_L g1954 ( 
.A(n_1033),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1415),
.A2(n_834),
.B1(n_878),
.B2(n_881),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1225),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1415),
.A2(n_834),
.B1(n_878),
.B2(n_881),
.Y(n_1957)
);

INVx3_ASAP7_75t_L g1958 ( 
.A(n_978),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1225),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_1033),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1961)
);

BUFx3_ASAP7_75t_L g1962 ( 
.A(n_1315),
.Y(n_1962)
);

INVx5_ASAP7_75t_L g1963 ( 
.A(n_978),
.Y(n_1963)
);

OR2x6_ASAP7_75t_L g1964 ( 
.A(n_1056),
.B(n_1033),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1414),
.A2(n_305),
.B1(n_312),
.B2(n_901),
.Y(n_1966)
);

BUFx8_ASAP7_75t_L g1967 ( 
.A(n_1158),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1225),
.Y(n_1968)
);

INVxp67_ASAP7_75t_SL g1969 ( 
.A(n_1056),
.Y(n_1969)
);

INVx1_ASAP7_75t_SL g1970 ( 
.A(n_1002),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1413),
.B(n_330),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1972)
);

OAI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1415),
.A2(n_1414),
.B1(n_1182),
.B2(n_448),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1413),
.B(n_330),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1413),
.B(n_330),
.Y(n_1976)
);

NOR2xp67_ASAP7_75t_L g1977 ( 
.A(n_1375),
.B(n_1365),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1225),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1182),
.B(n_1415),
.Y(n_1980)
);

NAND3xp33_ASAP7_75t_SL g1981 ( 
.A(n_1415),
.B(n_323),
.C(n_319),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1315),
.Y(n_1983)
);

CKINVDCx6p67_ASAP7_75t_R g1984 ( 
.A(n_1049),
.Y(n_1984)
);

INVx2_ASAP7_75t_SL g1985 ( 
.A(n_1033),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1225),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_993),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1056),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1225),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1225),
.Y(n_1990)
);

AOI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1415),
.A2(n_834),
.B1(n_878),
.B2(n_881),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1225),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1225),
.Y(n_1994)
);

INVx3_ASAP7_75t_L g1995 ( 
.A(n_978),
.Y(n_1995)
);

NAND2xp33_ASAP7_75t_L g1996 ( 
.A(n_1113),
.B(n_513),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1411),
.B(n_1412),
.Y(n_1997)
);

INVxp67_ASAP7_75t_L g1998 ( 
.A(n_996),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_979),
.B(n_980),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1045),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1804),
.A2(n_1858),
.B1(n_1924),
.B2(n_1914),
.Y(n_2001)
);

XOR2xp5_ASAP7_75t_L g2002 ( 
.A(n_1934),
.B(n_1966),
.Y(n_2002)
);

AND2x6_ASAP7_75t_L g2003 ( 
.A(n_1727),
.B(n_1581),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1454),
.B(n_1993),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1931),
.A2(n_1465),
.B(n_1516),
.Y(n_2005)
);

OAI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1800),
.A2(n_1868),
.B1(n_1872),
.B2(n_1863),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1429),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1997),
.B(n_1427),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1481),
.Y(n_2009)
);

A2O1A1Ixp33_ASAP7_75t_L g2010 ( 
.A1(n_1931),
.A2(n_1800),
.B(n_1868),
.C(n_1863),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1872),
.A2(n_1886),
.B1(n_1955),
.B2(n_1917),
.Y(n_2011)
);

OAI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1808),
.A2(n_1920),
.B(n_1917),
.Y(n_2012)
);

BUFx12f_ASAP7_75t_L g2013 ( 
.A(n_1557),
.Y(n_2013)
);

OR2x6_ASAP7_75t_L g2014 ( 
.A(n_1419),
.B(n_1424),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1831),
.B(n_1833),
.Y(n_2015)
);

O2A1O1Ixp33_ASAP7_75t_SL g2016 ( 
.A1(n_1808),
.A2(n_1920),
.B(n_1819),
.C(n_1889),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1838),
.B(n_1841),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1886),
.A2(n_1957),
.B1(n_1991),
.B2(n_1955),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1429),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1844),
.B(n_1846),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1957),
.A2(n_1991),
.B1(n_1421),
.B2(n_1879),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1429),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1936),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1828),
.A2(n_1879),
.B1(n_1973),
.B2(n_1470),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1849),
.B(n_1873),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1768),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_R g2027 ( 
.A(n_1823),
.B(n_1824),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1878),
.B(n_1883),
.Y(n_2028)
);

A2O1A1Ixp33_ASAP7_75t_L g2029 ( 
.A1(n_1421),
.A2(n_1996),
.B(n_1894),
.C(n_1909),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1458),
.B(n_1460),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1526),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1738),
.A2(n_1526),
.B(n_1522),
.Y(n_2032)
);

OAI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1826),
.A2(n_1916),
.B(n_1915),
.Y(n_2033)
);

AO21x1_ASAP7_75t_L g2034 ( 
.A1(n_1457),
.A2(n_1933),
.B(n_1928),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1828),
.A2(n_1940),
.B1(n_1972),
.B2(n_1946),
.Y(n_2035)
);

OAI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1980),
.A2(n_1534),
.B(n_1449),
.Y(n_2036)
);

HB1xp67_ASAP7_75t_L g2037 ( 
.A(n_1440),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1885),
.B(n_1893),
.Y(n_2038)
);

CKINVDCx20_ASAP7_75t_R g2039 ( 
.A(n_1950),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_1738),
.A2(n_1512),
.B(n_1725),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1497),
.B(n_1473),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1982),
.B(n_1896),
.Y(n_2042)
);

A2O1A1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_1512),
.A2(n_1583),
.B(n_1482),
.C(n_1699),
.Y(n_2043)
);

AOI21x1_ASAP7_75t_L g2044 ( 
.A1(n_1789),
.A2(n_1797),
.B(n_1795),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1441),
.Y(n_2045)
);

BUFx12f_ASAP7_75t_L g2046 ( 
.A(n_2000),
.Y(n_2046)
);

OAI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1798),
.A2(n_1853),
.B(n_1803),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1882),
.B(n_1922),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1470),
.A2(n_1988),
.B1(n_1508),
.B2(n_1479),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_1431),
.A2(n_1457),
.B1(n_1547),
.B2(n_1437),
.Y(n_2050)
);

AOI21x1_ASAP7_75t_L g2051 ( 
.A1(n_1797),
.A2(n_1795),
.B(n_1654),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1738),
.A2(n_1512),
.B(n_1725),
.Y(n_2052)
);

O2A1O1Ixp33_ASAP7_75t_L g2053 ( 
.A1(n_1428),
.A2(n_1861),
.B(n_1981),
.C(n_1809),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1912),
.B(n_1918),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_SL g2055 ( 
.A(n_1782),
.B(n_1551),
.Y(n_2055)
);

OAI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_1494),
.A2(n_1971),
.B1(n_1974),
.B2(n_1932),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1768),
.Y(n_2057)
);

BUFx6f_ASAP7_75t_L g2058 ( 
.A(n_1486),
.Y(n_2058)
);

BUFx2_ASAP7_75t_L g2059 ( 
.A(n_1779),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_1976),
.A2(n_1435),
.B1(n_1927),
.B2(n_1925),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_1475),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1937),
.B(n_1938),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1441),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1487),
.B(n_1455),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1942),
.B(n_1961),
.Y(n_2065)
);

BUFx10_ASAP7_75t_L g2066 ( 
.A(n_1474),
.Y(n_2066)
);

AO21x1_ASAP7_75t_L g2067 ( 
.A1(n_1693),
.A2(n_1633),
.B(n_1496),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1965),
.B(n_1975),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1441),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1978),
.B(n_1840),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1725),
.A2(n_1584),
.B(n_1551),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_1426),
.Y(n_2072)
);

NAND2x1p5_ASAP7_75t_L g2073 ( 
.A(n_1725),
.B(n_1762),
.Y(n_2073)
);

O2A1O1Ixp33_ASAP7_75t_L g2074 ( 
.A1(n_1430),
.A2(n_1483),
.B(n_1488),
.C(n_1810),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1466),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1486),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_L g2077 ( 
.A(n_1822),
.B(n_1903),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1466),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1840),
.B(n_1448),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1784),
.A2(n_1903),
.B1(n_1434),
.B2(n_1638),
.Y(n_2080)
);

AOI21xp5_ASAP7_75t_L g2081 ( 
.A1(n_1673),
.A2(n_1784),
.B(n_1525),
.Y(n_2081)
);

OAI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1517),
.A2(n_1606),
.B(n_1525),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1638),
.B(n_1728),
.Y(n_2083)
);

OAI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_1784),
.A2(n_1547),
.B1(n_1822),
.B2(n_1489),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1493),
.B(n_1446),
.Y(n_2085)
);

NAND2x1p5_ASAP7_75t_L g2086 ( 
.A(n_1762),
.B(n_1673),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1779),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1827),
.B(n_1876),
.Y(n_2088)
);

OAI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1784),
.A2(n_1822),
.B1(n_1683),
.B2(n_1580),
.Y(n_2089)
);

A2O1A1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_1583),
.A2(n_1482),
.B(n_1629),
.C(n_1571),
.Y(n_2090)
);

O2A1O1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_1816),
.A2(n_1850),
.B(n_1880),
.C(n_1860),
.Y(n_2091)
);

NOR2xp67_ASAP7_75t_L g2092 ( 
.A(n_1673),
.B(n_1762),
.Y(n_2092)
);

AO32x1_ASAP7_75t_L g2093 ( 
.A1(n_1750),
.A2(n_1797),
.A3(n_1597),
.B1(n_1604),
.B2(n_1565),
.Y(n_2093)
);

CKINVDCx8_ASAP7_75t_R g2094 ( 
.A(n_1438),
.Y(n_2094)
);

OAI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1683),
.A2(n_1580),
.B1(n_1507),
.B2(n_1606),
.Y(n_2095)
);

AOI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_1749),
.A2(n_1591),
.B(n_1519),
.Y(n_2096)
);

AOI21xp5_ASAP7_75t_L g2097 ( 
.A1(n_1712),
.A2(n_1719),
.B(n_1661),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1456),
.B(n_1462),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_1432),
.A2(n_1859),
.B1(n_1874),
.B2(n_1450),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1467),
.B(n_1469),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1425),
.Y(n_2101)
);

INVx4_ASAP7_75t_L g2102 ( 
.A(n_1814),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1589),
.B(n_1818),
.Y(n_2103)
);

BUFx3_ASAP7_75t_L g2104 ( 
.A(n_1475),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1589),
.B(n_1818),
.Y(n_2105)
);

BUFx4f_ASAP7_75t_L g2106 ( 
.A(n_1418),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1899),
.B(n_1907),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_1712),
.A2(n_1719),
.B(n_1661),
.Y(n_2108)
);

OAI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_1751),
.A2(n_1442),
.B(n_1723),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1899),
.B(n_1907),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1999),
.B(n_1892),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1999),
.B(n_1892),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1970),
.B(n_1634),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_1827),
.B(n_1876),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_1432),
.B(n_1450),
.Y(n_2115)
);

INVx11_ASAP7_75t_L g2116 ( 
.A(n_1475),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1970),
.B(n_1634),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1609),
.B(n_1618),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_1727),
.A2(n_1658),
.B(n_1669),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_L g2120 ( 
.A(n_1432),
.B(n_1450),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1859),
.A2(n_1962),
.B1(n_1983),
.B2(n_1874),
.Y(n_2121)
);

OAI21xp33_ASAP7_75t_L g2122 ( 
.A1(n_1632),
.A2(n_1751),
.B(n_1729),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1609),
.B(n_1618),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1554),
.B(n_1542),
.Y(n_2124)
);

AOI21xp5_ASAP7_75t_L g2125 ( 
.A1(n_1727),
.A2(n_1669),
.B(n_1649),
.Y(n_2125)
);

BUFx12f_ASAP7_75t_L g2126 ( 
.A(n_1475),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_1669),
.A2(n_1750),
.B(n_1710),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1554),
.B(n_1542),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_1783),
.A2(n_1603),
.B(n_1599),
.Y(n_2129)
);

O2A1O1Ixp33_ASAP7_75t_L g2130 ( 
.A1(n_1952),
.A2(n_1987),
.B(n_1562),
.C(n_1597),
.Y(n_2130)
);

OR2x2_ASAP7_75t_L g2131 ( 
.A(n_1884),
.B(n_1988),
.Y(n_2131)
);

O2A1O1Ixp33_ASAP7_75t_L g2132 ( 
.A1(n_1565),
.A2(n_1604),
.B(n_1484),
.C(n_1621),
.Y(n_2132)
);

NOR2xp33_ASAP7_75t_L g2133 ( 
.A(n_1859),
.B(n_1874),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_1962),
.B(n_1983),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1595),
.B(n_1461),
.Y(n_2135)
);

O2A1O1Ixp33_ASAP7_75t_SL g2136 ( 
.A1(n_1646),
.A2(n_1743),
.B(n_1765),
.C(n_1757),
.Y(n_2136)
);

BUFx4f_ASAP7_75t_L g2137 ( 
.A(n_1418),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1425),
.Y(n_2138)
);

AOI22xp5_ASAP7_75t_L g2139 ( 
.A1(n_1470),
.A2(n_1632),
.B1(n_1442),
.B2(n_1737),
.Y(n_2139)
);

O2A1O1Ixp33_ASAP7_75t_L g2140 ( 
.A1(n_1511),
.A2(n_1698),
.B(n_1701),
.C(n_1668),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_1962),
.B(n_1983),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1461),
.B(n_1480),
.Y(n_2142)
);

CKINVDCx6p67_ASAP7_75t_R g2143 ( 
.A(n_1984),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1884),
.B(n_1451),
.Y(n_2144)
);

AO21x1_ASAP7_75t_L g2145 ( 
.A1(n_1559),
.A2(n_1592),
.B(n_1767),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1998),
.B(n_1605),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_1783),
.A2(n_1614),
.B(n_1612),
.Y(n_2147)
);

A2O1A1Ixp33_ASAP7_75t_L g2148 ( 
.A1(n_1628),
.A2(n_1665),
.B(n_1758),
.C(n_1778),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1605),
.B(n_1576),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1576),
.B(n_1502),
.Y(n_2150)
);

XOR2xp5_ASAP7_75t_L g2151 ( 
.A(n_1491),
.B(n_1546),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1470),
.A2(n_1737),
.B1(n_1546),
.B2(n_1505),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1436),
.Y(n_2153)
);

AOI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_1617),
.A2(n_1619),
.B(n_1854),
.Y(n_2154)
);

NOR2xp33_ASAP7_75t_L g2155 ( 
.A(n_1984),
.B(n_1477),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_SL g2156 ( 
.A(n_1648),
.B(n_1753),
.Y(n_2156)
);

OAI22xp5_ASAP7_75t_L g2157 ( 
.A1(n_1529),
.A2(n_1665),
.B1(n_1690),
.B2(n_1642),
.Y(n_2157)
);

AOI21xp5_ASAP7_75t_L g2158 ( 
.A1(n_1854),
.A2(n_1906),
.B(n_1637),
.Y(n_2158)
);

AOI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_1470),
.A2(n_1737),
.B1(n_1505),
.B2(n_1761),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_1477),
.B(n_1438),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_1477),
.B(n_1485),
.Y(n_2161)
);

INVx4_ASAP7_75t_L g2162 ( 
.A(n_1814),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_1485),
.B(n_1491),
.Y(n_2163)
);

NOR2xp67_ASAP7_75t_SL g2164 ( 
.A(n_1814),
.B(n_1902),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_1906),
.A2(n_1637),
.B(n_1520),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1503),
.B(n_1540),
.Y(n_2166)
);

INVxp67_ASAP7_75t_L g2167 ( 
.A(n_1653),
.Y(n_2167)
);

CKINVDCx20_ASAP7_75t_R g2168 ( 
.A(n_1821),
.Y(n_2168)
);

A2O1A1Ixp33_ASAP7_75t_L g2169 ( 
.A1(n_1758),
.A2(n_1772),
.B(n_1682),
.C(n_1550),
.Y(n_2169)
);

OAI21xp33_ASAP7_75t_L g2170 ( 
.A1(n_1763),
.A2(n_1587),
.B(n_1567),
.Y(n_2170)
);

AOI21x1_ASAP7_75t_L g2171 ( 
.A1(n_1598),
.A2(n_1769),
.B(n_1773),
.Y(n_2171)
);

NOR3xp33_ASAP7_75t_L g2172 ( 
.A(n_1543),
.B(n_1708),
.C(n_1785),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1747),
.B(n_1640),
.Y(n_2173)
);

AOI22xp33_ASAP7_75t_L g2174 ( 
.A1(n_1470),
.A2(n_1505),
.B1(n_1782),
.B2(n_1506),
.Y(n_2174)
);

AOI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_1762),
.A2(n_1666),
.B(n_1659),
.Y(n_2175)
);

NAND2x1p5_ASAP7_75t_L g2176 ( 
.A(n_1762),
.B(n_1472),
.Y(n_2176)
);

AOI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_1762),
.A2(n_1666),
.B(n_1659),
.Y(n_2177)
);

INVx4_ASAP7_75t_L g2178 ( 
.A(n_1814),
.Y(n_2178)
);

CKINVDCx20_ASAP7_75t_R g2179 ( 
.A(n_1509),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1451),
.B(n_1422),
.Y(n_2180)
);

AOI21xp5_ASAP7_75t_L g2181 ( 
.A1(n_1659),
.A2(n_1692),
.B(n_1666),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1747),
.B(n_1735),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_1470),
.A2(n_1505),
.B1(n_1782),
.B2(n_1506),
.Y(n_2183)
);

BUFx8_ASAP7_75t_L g2184 ( 
.A(n_1664),
.Y(n_2184)
);

AOI21x1_ASAP7_75t_L g2185 ( 
.A1(n_1598),
.A2(n_1788),
.B(n_1663),
.Y(n_2185)
);

AND2x4_ASAP7_75t_L g2186 ( 
.A(n_1458),
.B(n_1460),
.Y(n_2186)
);

AOI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_1659),
.A2(n_1692),
.B(n_1666),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1422),
.B(n_1423),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1735),
.B(n_1532),
.Y(n_2189)
);

OAI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_1788),
.A2(n_1790),
.B(n_1721),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1436),
.Y(n_2191)
);

OAI21x1_ASAP7_75t_L g2192 ( 
.A1(n_1771),
.A2(n_1709),
.B(n_1787),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1532),
.B(n_1548),
.Y(n_2193)
);

OAI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_1574),
.A2(n_1792),
.B(n_1791),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1548),
.B(n_1558),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1558),
.B(n_1611),
.Y(n_2196)
);

NAND3xp33_ASAP7_75t_L g2197 ( 
.A(n_1754),
.B(n_1777),
.C(n_1775),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1611),
.B(n_1676),
.Y(n_2198)
);

O2A1O1Ixp33_ASAP7_75t_L g2199 ( 
.A1(n_1569),
.A2(n_1664),
.B(n_1793),
.C(n_1513),
.Y(n_2199)
);

CKINVDCx11_ASAP7_75t_R g2200 ( 
.A(n_1726),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1447),
.Y(n_2201)
);

AND2x4_ASAP7_75t_L g2202 ( 
.A(n_1458),
.B(n_1460),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1498),
.B(n_1579),
.Y(n_2203)
);

OAI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_1529),
.A2(n_1690),
.B1(n_1594),
.B2(n_1561),
.Y(n_2204)
);

HB1xp67_ASAP7_75t_L g2205 ( 
.A(n_1647),
.Y(n_2205)
);

A2O1A1Ixp33_ASAP7_75t_L g2206 ( 
.A1(n_1568),
.A2(n_1777),
.B(n_1775),
.C(n_1572),
.Y(n_2206)
);

AOI21xp5_ASAP7_75t_L g2207 ( 
.A1(n_1692),
.A2(n_1703),
.B(n_1766),
.Y(n_2207)
);

AOI21x1_ASAP7_75t_L g2208 ( 
.A1(n_1780),
.A2(n_1774),
.B(n_1722),
.Y(n_2208)
);

BUFx6f_ASAP7_75t_L g2209 ( 
.A(n_1472),
.Y(n_2209)
);

BUFx4f_ASAP7_75t_L g2210 ( 
.A(n_1418),
.Y(n_2210)
);

OAI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_1791),
.A2(n_1792),
.B(n_1541),
.Y(n_2211)
);

AOI21x1_ASAP7_75t_L g2212 ( 
.A1(n_1722),
.A2(n_1439),
.B(n_1433),
.Y(n_2212)
);

NAND2xp33_ASAP7_75t_L g2213 ( 
.A(n_1470),
.B(n_1505),
.Y(n_2213)
);

NOR3xp33_ASAP7_75t_L g2214 ( 
.A(n_1793),
.B(n_1513),
.C(n_1492),
.Y(n_2214)
);

AOI21x1_ASAP7_75t_L g2215 ( 
.A1(n_1722),
.A2(n_1439),
.B(n_1433),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1447),
.Y(n_2216)
);

OAI22xp33_ASAP7_75t_L g2217 ( 
.A1(n_1506),
.A2(n_1556),
.B1(n_1564),
.B2(n_1424),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1648),
.B(n_1753),
.Y(n_2218)
);

NOR2xp33_ASAP7_75t_L g2219 ( 
.A(n_1492),
.B(n_1537),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_1703),
.A2(n_1541),
.B(n_1714),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1498),
.B(n_1579),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_1761),
.A2(n_1745),
.B1(n_1572),
.B2(n_1799),
.Y(n_2222)
);

AOI21xp5_ASAP7_75t_L g2223 ( 
.A1(n_1703),
.A2(n_1714),
.B(n_1552),
.Y(n_2223)
);

AO21x1_ASAP7_75t_L g2224 ( 
.A1(n_1799),
.A2(n_1812),
.B(n_1807),
.Y(n_2224)
);

INVx3_ASAP7_75t_L g2225 ( 
.A(n_1478),
.Y(n_2225)
);

NAND3xp33_ASAP7_75t_L g2226 ( 
.A(n_1782),
.B(n_1812),
.C(n_1807),
.Y(n_2226)
);

AOI21xp5_ASAP7_75t_L g2227 ( 
.A1(n_1714),
.A2(n_1552),
.B(n_1539),
.Y(n_2227)
);

OAI21xp5_ASAP7_75t_L g2228 ( 
.A1(n_1575),
.A2(n_1792),
.B(n_1791),
.Y(n_2228)
);

OAI21xp5_ASAP7_75t_L g2229 ( 
.A1(n_1681),
.A2(n_1817),
.B(n_1813),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1422),
.B(n_1423),
.Y(n_2230)
);

NAND2x1p5_ASAP7_75t_L g2231 ( 
.A(n_1472),
.B(n_1536),
.Y(n_2231)
);

INVx5_ASAP7_75t_L g2232 ( 
.A(n_1505),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_1423),
.B(n_1801),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1613),
.B(n_1616),
.Y(n_2234)
);

CKINVDCx8_ASAP7_75t_R g2235 ( 
.A(n_1726),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1453),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_R g2237 ( 
.A(n_1509),
.B(n_1852),
.Y(n_2237)
);

OAI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_1761),
.A2(n_1745),
.B1(n_1817),
.B2(n_1813),
.Y(n_2238)
);

HB1xp67_ASAP7_75t_L g2239 ( 
.A(n_1647),
.Y(n_2239)
);

NOR2x1_ASAP7_75t_L g2240 ( 
.A(n_1714),
.B(n_1755),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_1801),
.B(n_1815),
.Y(n_2241)
);

AOI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_1505),
.A2(n_1761),
.B1(n_1506),
.B2(n_1553),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_1613),
.B(n_1616),
.Y(n_2243)
);

O2A1O1Ixp33_ASAP7_75t_L g2244 ( 
.A1(n_1537),
.A2(n_1832),
.B(n_1843),
.C(n_1825),
.Y(n_2244)
);

A2O1A1Ixp33_ASAP7_75t_L g2245 ( 
.A1(n_1553),
.A2(n_1829),
.B(n_1913),
.C(n_1802),
.Y(n_2245)
);

NAND3xp33_ASAP7_75t_L g2246 ( 
.A(n_1825),
.B(n_1843),
.C(n_1832),
.Y(n_2246)
);

NOR3xp33_ASAP7_75t_L g2247 ( 
.A(n_1745),
.B(n_1615),
.C(n_1510),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_1478),
.Y(n_2248)
);

INVxp67_ASAP7_75t_L g2249 ( 
.A(n_1644),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_1472),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_1505),
.A2(n_1506),
.B1(n_1553),
.B2(n_1460),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_L g2252 ( 
.A(n_1509),
.B(n_1852),
.Y(n_2252)
);

OAI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_1745),
.A2(n_1848),
.B1(n_1865),
.B2(n_1856),
.Y(n_2253)
);

NOR3xp33_ASAP7_75t_L g2254 ( 
.A(n_1615),
.B(n_1510),
.C(n_1500),
.Y(n_2254)
);

AOI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_1539),
.A2(n_1552),
.B(n_1875),
.Y(n_2255)
);

O2A1O1Ixp33_ASAP7_75t_L g2256 ( 
.A1(n_1848),
.A2(n_1856),
.B(n_1867),
.C(n_1865),
.Y(n_2256)
);

AO21x2_ASAP7_75t_L g2257 ( 
.A1(n_1514),
.A2(n_1528),
.B(n_1518),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_1630),
.B(n_1675),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_1801),
.B(n_1815),
.Y(n_2259)
);

AOI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_1458),
.A2(n_1806),
.B1(n_1830),
.B2(n_1524),
.Y(n_2260)
);

AOI33xp33_ASAP7_75t_L g2261 ( 
.A1(n_1867),
.A2(n_1871),
.A3(n_1953),
.B1(n_1992),
.B2(n_1990),
.B3(n_1948),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1630),
.B(n_1675),
.Y(n_2262)
);

AOI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_1524),
.A2(n_1830),
.B1(n_1837),
.B2(n_1806),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_1539),
.A2(n_1552),
.B(n_1875),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1644),
.B(n_1815),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_1839),
.B(n_1851),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_1509),
.B(n_1852),
.Y(n_2267)
);

OAI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_1871),
.A2(n_1877),
.B1(n_1888),
.B2(n_1887),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1839),
.B(n_1851),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_1852),
.B(n_1967),
.Y(n_2270)
);

NOR2xp33_ASAP7_75t_L g2271 ( 
.A(n_1967),
.B(n_1539),
.Y(n_2271)
);

A2O1A1Ixp33_ASAP7_75t_L g2272 ( 
.A1(n_1969),
.A2(n_1556),
.B(n_1755),
.C(n_1770),
.Y(n_2272)
);

AO22x1_ASAP7_75t_L g2273 ( 
.A1(n_1967),
.A2(n_1556),
.B1(n_1776),
.B2(n_1746),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1839),
.B(n_1851),
.Y(n_2274)
);

A2O1A1Ixp33_ASAP7_75t_L g2275 ( 
.A1(n_1770),
.A2(n_1877),
.B(n_1888),
.C(n_1887),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1857),
.B(n_1864),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_1524),
.B(n_1806),
.Y(n_2277)
);

O2A1O1Ixp33_ASAP7_75t_L g2278 ( 
.A1(n_1895),
.A2(n_1901),
.B(n_1923),
.C(n_1919),
.Y(n_2278)
);

INVx5_ASAP7_75t_L g2279 ( 
.A(n_1419),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1857),
.B(n_1864),
.Y(n_2280)
);

AOI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_1875),
.A2(n_1678),
.B(n_1680),
.Y(n_2281)
);

AOI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_1678),
.A2(n_1680),
.B(n_1684),
.Y(n_2282)
);

AOI22xp33_ASAP7_75t_L g2283 ( 
.A1(n_1419),
.A2(n_1424),
.B1(n_1908),
.B2(n_1834),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_1678),
.A2(n_1680),
.B(n_1684),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1857),
.B(n_1864),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1869),
.B(n_1881),
.Y(n_2286)
);

INVx1_ASAP7_75t_SL g2287 ( 
.A(n_1730),
.Y(n_2287)
);

AO21x1_ASAP7_75t_L g2288 ( 
.A1(n_1895),
.A2(n_1919),
.B(n_1901),
.Y(n_2288)
);

BUFx12f_ASAP7_75t_L g2289 ( 
.A(n_1967),
.Y(n_2289)
);

NAND2xp33_ASAP7_75t_L g2290 ( 
.A(n_1814),
.B(n_1902),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_1524),
.B(n_1806),
.Y(n_2291)
);

NOR2x1_ASAP7_75t_L g2292 ( 
.A(n_1471),
.B(n_1476),
.Y(n_2292)
);

INVxp67_ASAP7_75t_L g2293 ( 
.A(n_1643),
.Y(n_2293)
);

OAI21xp33_ASAP7_75t_L g2294 ( 
.A1(n_1923),
.A2(n_1930),
.B(n_1926),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_1869),
.B(n_1881),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_1830),
.B(n_1837),
.Y(n_2296)
);

AOI21xp5_ASAP7_75t_L g2297 ( 
.A1(n_1724),
.A2(n_1759),
.B(n_1535),
.Y(n_2297)
);

AO21x1_ASAP7_75t_L g2298 ( 
.A1(n_1926),
.A2(n_1935),
.B(n_1930),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1453),
.Y(n_2299)
);

NOR2xp67_ASAP7_75t_L g2300 ( 
.A(n_1472),
.B(n_1536),
.Y(n_2300)
);

BUFx2_ASAP7_75t_L g2301 ( 
.A(n_1722),
.Y(n_2301)
);

INVx4_ASAP7_75t_L g2302 ( 
.A(n_1814),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_1891),
.B(n_1897),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_1891),
.B(n_1897),
.Y(n_2304)
);

INVx4_ASAP7_75t_L g2305 ( 
.A(n_1902),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1490),
.Y(n_2306)
);

A2O1A1Ixp33_ASAP7_75t_L g2307 ( 
.A1(n_1770),
.A2(n_1935),
.B(n_1948),
.C(n_1945),
.Y(n_2307)
);

AOI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_1478),
.A2(n_1625),
.B(n_1535),
.Y(n_2308)
);

AOI21xp5_ASAP7_75t_L g2309 ( 
.A1(n_1478),
.A2(n_1625),
.B(n_1535),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1891),
.B(n_1897),
.Y(n_2310)
);

NOR2xp67_ASAP7_75t_L g2311 ( 
.A(n_1472),
.B(n_1536),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1459),
.Y(n_2312)
);

INVx1_ASAP7_75t_SL g2313 ( 
.A(n_1730),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1904),
.B(n_1943),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_1830),
.B(n_1837),
.Y(n_2315)
);

AOI22xp33_ASAP7_75t_L g2316 ( 
.A1(n_1419),
.A2(n_1424),
.B1(n_1908),
.B2(n_1834),
.Y(n_2316)
);

AOI21xp5_ASAP7_75t_L g2317 ( 
.A1(n_1535),
.A2(n_1625),
.B(n_1495),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_1904),
.B(n_1943),
.Y(n_2318)
);

A2O1A1Ixp33_ASAP7_75t_L g2319 ( 
.A1(n_1945),
.A2(n_1953),
.B(n_1959),
.C(n_1956),
.Y(n_2319)
);

O2A1O1Ixp33_ASAP7_75t_L g2320 ( 
.A1(n_1956),
.A2(n_1968),
.B(n_1979),
.C(n_1959),
.Y(n_2320)
);

BUFx6f_ASAP7_75t_L g2321 ( 
.A(n_1536),
.Y(n_2321)
);

INVx1_ASAP7_75t_SL g2322 ( 
.A(n_1523),
.Y(n_2322)
);

O2A1O1Ixp33_ASAP7_75t_L g2323 ( 
.A1(n_1968),
.A2(n_1986),
.B(n_1990),
.C(n_1979),
.Y(n_2323)
);

NOR2xp67_ASAP7_75t_SL g2324 ( 
.A(n_1902),
.B(n_1963),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1501),
.Y(n_2325)
);

A2O1A1Ixp33_ASAP7_75t_L g2326 ( 
.A1(n_1986),
.A2(n_1992),
.B(n_1523),
.C(n_1994),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_1625),
.A2(n_1495),
.B(n_1862),
.Y(n_2327)
);

AOI21xp5_ASAP7_75t_L g2328 ( 
.A1(n_1495),
.A2(n_1870),
.B(n_1862),
.Y(n_2328)
);

AOI21xp5_ASAP7_75t_L g2329 ( 
.A1(n_1495),
.A2(n_1870),
.B(n_1862),
.Y(n_2329)
);

AOI21xp5_ASAP7_75t_L g2330 ( 
.A1(n_1862),
.A2(n_1910),
.B(n_1870),
.Y(n_2330)
);

AOI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_1870),
.A2(n_1929),
.B(n_1910),
.Y(n_2331)
);

AND2x4_ASAP7_75t_L g2332 ( 
.A(n_1910),
.B(n_1929),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1947),
.B(n_1949),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_1910),
.A2(n_1951),
.B(n_1929),
.Y(n_2334)
);

O2A1O1Ixp33_ASAP7_75t_L g2335 ( 
.A1(n_1995),
.A2(n_1939),
.B(n_1921),
.C(n_1911),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_1947),
.B(n_1949),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1947),
.B(n_1949),
.Y(n_2337)
);

A2O1A1Ixp33_ASAP7_75t_L g2338 ( 
.A1(n_1989),
.A2(n_1994),
.B(n_1781),
.C(n_1794),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_1989),
.B(n_1994),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_1501),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_1929),
.A2(n_1951),
.B(n_1420),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1459),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1501),
.Y(n_2343)
);

BUFx6f_ASAP7_75t_L g2344 ( 
.A(n_1536),
.Y(n_2344)
);

AOI21xp5_ASAP7_75t_L g2345 ( 
.A1(n_1951),
.A2(n_1420),
.B(n_1641),
.Y(n_2345)
);

NAND3xp33_ASAP7_75t_L g2346 ( 
.A(n_1786),
.B(n_1681),
.C(n_1679),
.Y(n_2346)
);

AOI21xp5_ASAP7_75t_L g2347 ( 
.A1(n_1951),
.A2(n_1420),
.B(n_1641),
.Y(n_2347)
);

BUFx6f_ASAP7_75t_L g2348 ( 
.A(n_1536),
.Y(n_2348)
);

AOI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_1641),
.A2(n_1578),
.B(n_1544),
.Y(n_2349)
);

INVxp67_ASAP7_75t_L g2350 ( 
.A(n_1643),
.Y(n_2350)
);

NOR2xp67_ASAP7_75t_SL g2351 ( 
.A(n_1902),
.B(n_1963),
.Y(n_2351)
);

AOI21xp5_ASAP7_75t_L g2352 ( 
.A1(n_1641),
.A2(n_1578),
.B(n_1544),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1499),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_SL g2354 ( 
.A(n_1627),
.B(n_1443),
.Y(n_2354)
);

AOI21xp33_ASAP7_75t_L g2355 ( 
.A1(n_1748),
.A2(n_1756),
.B(n_1752),
.Y(n_2355)
);

AOI22xp33_ASAP7_75t_L g2356 ( 
.A1(n_1419),
.A2(n_1908),
.B1(n_1424),
.B2(n_1834),
.Y(n_2356)
);

O2A1O1Ixp33_ASAP7_75t_L g2357 ( 
.A1(n_1445),
.A2(n_1995),
.B(n_1911),
.C(n_1921),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_1643),
.B(n_1652),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_1652),
.B(n_1504),
.Y(n_2359)
);

OAI22xp5_ASAP7_75t_L g2360 ( 
.A1(n_1577),
.A2(n_1834),
.B1(n_1908),
.B2(n_1964),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_1504),
.B(n_1748),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_1652),
.B(n_1627),
.Y(n_2362)
);

HB1xp67_ASAP7_75t_L g2363 ( 
.A(n_1671),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1752),
.B(n_1756),
.Y(n_2364)
);

OAI22xp5_ASAP7_75t_L g2365 ( 
.A1(n_1577),
.A2(n_1908),
.B1(n_1964),
.B2(n_1834),
.Y(n_2365)
);

BUFx8_ASAP7_75t_L g2366 ( 
.A(n_1418),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1760),
.B(n_1764),
.Y(n_2367)
);

AOI21xp5_ASAP7_75t_L g2368 ( 
.A1(n_1544),
.A2(n_1582),
.B(n_1578),
.Y(n_2368)
);

AOI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_1544),
.A2(n_1582),
.B(n_1578),
.Y(n_2369)
);

INVx1_ASAP7_75t_SL g2370 ( 
.A(n_1781),
.Y(n_2370)
);

NOR2xp33_ASAP7_75t_L g2371 ( 
.A(n_1627),
.B(n_1586),
.Y(n_2371)
);

AOI21x1_ASAP7_75t_L g2372 ( 
.A1(n_1722),
.A2(n_1890),
.B(n_1866),
.Y(n_2372)
);

OAI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_1577),
.A2(n_1964),
.B1(n_1564),
.B2(n_1445),
.Y(n_2373)
);

AOI21xp5_ASAP7_75t_L g2374 ( 
.A1(n_1582),
.A2(n_1476),
.B(n_1471),
.Y(n_2374)
);

INVx1_ASAP7_75t_SL g2375 ( 
.A(n_1586),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_1760),
.B(n_1764),
.Y(n_2376)
);

INVx1_ASAP7_75t_SL g2377 ( 
.A(n_1586),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1514),
.B(n_1518),
.Y(n_2378)
);

NOR2x1p5_ASAP7_75t_SL g2379 ( 
.A(n_1528),
.B(n_1531),
.Y(n_2379)
);

HB1xp67_ASAP7_75t_L g2380 ( 
.A(n_1687),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1531),
.B(n_1657),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_1581),
.A2(n_1590),
.B(n_1510),
.Y(n_2382)
);

AOI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_1581),
.A2(n_1590),
.B(n_1533),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1563),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_1515),
.Y(n_2385)
);

INVx5_ASAP7_75t_L g2386 ( 
.A(n_1964),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_1657),
.B(n_1691),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1515),
.Y(n_2388)
);

NOR2xp33_ASAP7_75t_L g2389 ( 
.A(n_1600),
.B(n_1602),
.Y(n_2389)
);

AOI21xp5_ASAP7_75t_L g2390 ( 
.A1(n_1581),
.A2(n_1590),
.B(n_1533),
.Y(n_2390)
);

NAND2x1_ASAP7_75t_L g2391 ( 
.A(n_1577),
.B(n_1500),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_1691),
.B(n_1694),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_1694),
.B(n_1707),
.Y(n_2393)
);

AOI21xp5_ASAP7_75t_L g2394 ( 
.A1(n_1590),
.A2(n_1631),
.B(n_1902),
.Y(n_2394)
);

AOI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_1631),
.A2(n_1963),
.B(n_1452),
.Y(n_2395)
);

AOI21xp5_ASAP7_75t_L g2396 ( 
.A1(n_1631),
.A2(n_1963),
.B(n_1463),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_1707),
.B(n_1716),
.Y(n_2397)
);

AOI22x1_ASAP7_75t_L g2398 ( 
.A1(n_1709),
.A2(n_1771),
.B1(n_1958),
.B2(n_1445),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_1964),
.B(n_1716),
.Y(n_2399)
);

CKINVDCx16_ASAP7_75t_R g2400 ( 
.A(n_1600),
.Y(n_2400)
);

OAI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_1577),
.A2(n_1564),
.B1(n_1921),
.B2(n_1464),
.Y(n_2401)
);

CKINVDCx20_ASAP7_75t_R g2402 ( 
.A(n_1610),
.Y(n_2402)
);

HB1xp67_ASAP7_75t_L g2403 ( 
.A(n_1600),
.Y(n_2403)
);

AOI21xp5_ASAP7_75t_L g2404 ( 
.A1(n_1963),
.A2(n_1977),
.B(n_1890),
.Y(n_2404)
);

INVxp67_ASAP7_75t_L g2405 ( 
.A(n_1689),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_1733),
.B(n_1741),
.Y(n_2406)
);

AOI21xp5_ASAP7_75t_L g2407 ( 
.A1(n_1602),
.A2(n_1709),
.B(n_1624),
.Y(n_2407)
);

AOI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_1624),
.A2(n_1444),
.B1(n_1443),
.B2(n_1954),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_L g2409 ( 
.A(n_1602),
.B(n_1443),
.Y(n_2409)
);

AO21x1_ASAP7_75t_L g2410 ( 
.A1(n_1771),
.A2(n_1624),
.B(n_1702),
.Y(n_2410)
);

NAND2x1p5_ASAP7_75t_L g2411 ( 
.A(n_1624),
.B(n_1443),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1566),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_1566),
.Y(n_2413)
);

OAI22xp5_ASAP7_75t_SL g2414 ( 
.A1(n_1585),
.A2(n_1549),
.B1(n_1718),
.B2(n_1444),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_SL g2415 ( 
.A(n_1820),
.B(n_1847),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1570),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_R g2417 ( 
.A(n_1820),
.B(n_1847),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_1468),
.A2(n_1995),
.B1(n_1958),
.B2(n_1939),
.Y(n_2418)
);

OAI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_1645),
.A2(n_1711),
.B(n_1689),
.Y(n_2419)
);

OA22x2_ASAP7_75t_L g2420 ( 
.A1(n_1685),
.A2(n_1985),
.B1(n_1960),
.B2(n_1805),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_1733),
.B(n_1741),
.Y(n_2421)
);

INVx4_ASAP7_75t_L g2422 ( 
.A(n_1820),
.Y(n_2422)
);

INVxp33_ASAP7_75t_SL g2423 ( 
.A(n_1794),
.Y(n_2423)
);

OAI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_1811),
.A2(n_1958),
.B1(n_1939),
.B2(n_1444),
.Y(n_2424)
);

NAND2x1p5_ASAP7_75t_L g2425 ( 
.A(n_1954),
.B(n_1794),
.Y(n_2425)
);

O2A1O1Ixp33_ASAP7_75t_L g2426 ( 
.A1(n_1958),
.A2(n_1711),
.B(n_1685),
.C(n_1944),
.Y(n_2426)
);

OAI22xp33_ASAP7_75t_L g2427 ( 
.A1(n_1954),
.A2(n_1444),
.B1(n_1985),
.B2(n_1960),
.Y(n_2427)
);

NAND2x1p5_ASAP7_75t_L g2428 ( 
.A(n_1796),
.B(n_1847),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_1521),
.Y(n_2429)
);

AOI21x1_ASAP7_75t_L g2430 ( 
.A1(n_1685),
.A2(n_1655),
.B(n_1731),
.Y(n_2430)
);

O2A1O1Ixp33_ASAP7_75t_L g2431 ( 
.A1(n_1685),
.A2(n_1944),
.B(n_1805),
.C(n_1845),
.Y(n_2431)
);

A2O1A1Ixp33_ASAP7_75t_L g2432 ( 
.A1(n_1835),
.A2(n_1836),
.B(n_1905),
.C(n_1900),
.Y(n_2432)
);

A2O1A1Ixp33_ASAP7_75t_SL g2433 ( 
.A1(n_1521),
.A2(n_1734),
.B(n_1527),
.C(n_1530),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_1593),
.B(n_1596),
.Y(n_2434)
);

OAI22xp5_ASAP7_75t_L g2435 ( 
.A1(n_1444),
.A2(n_1836),
.B1(n_1905),
.B2(n_1900),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_1521),
.Y(n_2436)
);

OAI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_1650),
.A2(n_1686),
.B(n_1674),
.Y(n_2437)
);

BUFx6f_ASAP7_75t_L g2438 ( 
.A(n_1847),
.Y(n_2438)
);

INVx1_ASAP7_75t_SL g2439 ( 
.A(n_1796),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_1596),
.B(n_1742),
.Y(n_2440)
);

OAI22xp5_ASAP7_75t_L g2441 ( 
.A1(n_1835),
.A2(n_1845),
.B1(n_1842),
.B2(n_1855),
.Y(n_2441)
);

A2O1A1Ixp33_ASAP7_75t_L g2442 ( 
.A1(n_1842),
.A2(n_1855),
.B(n_1677),
.C(n_1623),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_1688),
.A2(n_1941),
.B(n_1898),
.Y(n_2443)
);

AOI21xp5_ASAP7_75t_L g2444 ( 
.A1(n_1847),
.A2(n_1941),
.B(n_1898),
.Y(n_2444)
);

INVx4_ASAP7_75t_L g2445 ( 
.A(n_1898),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_1527),
.Y(n_2446)
);

AND2x2_ASAP7_75t_SL g2447 ( 
.A(n_1898),
.B(n_1941),
.Y(n_2447)
);

A2O1A1Ixp33_ASAP7_75t_L g2448 ( 
.A1(n_1608),
.A2(n_1623),
.B(n_1695),
.C(n_1662),
.Y(n_2448)
);

A2O1A1Ixp33_ASAP7_75t_L g2449 ( 
.A1(n_1608),
.A2(n_1622),
.B(n_1662),
.C(n_1742),
.Y(n_2449)
);

AOI221xp5_ASAP7_75t_L g2450 ( 
.A1(n_1620),
.A2(n_1697),
.B1(n_1739),
.B2(n_1732),
.C(n_1720),
.Y(n_2450)
);

O2A1O1Ixp33_ASAP7_75t_L g2451 ( 
.A1(n_1622),
.A2(n_1739),
.B(n_1732),
.C(n_1720),
.Y(n_2451)
);

AOI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_1796),
.A2(n_1527),
.B(n_1530),
.Y(n_2452)
);

O2A1O1Ixp33_ASAP7_75t_L g2453 ( 
.A1(n_1626),
.A2(n_1717),
.B(n_1715),
.C(n_1705),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_SL g2454 ( 
.A(n_1786),
.B(n_1776),
.Y(n_2454)
);

AOI21xp5_ASAP7_75t_L g2455 ( 
.A1(n_1538),
.A2(n_1545),
.B(n_1555),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_1639),
.B(n_1717),
.Y(n_2456)
);

OAI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_1667),
.A2(n_1713),
.B1(n_1670),
.B2(n_1700),
.Y(n_2457)
);

A2O1A1Ixp33_ASAP7_75t_L g2458 ( 
.A1(n_1651),
.A2(n_1700),
.B(n_1697),
.C(n_1660),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_1651),
.B(n_1660),
.Y(n_2459)
);

AOI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_1588),
.A2(n_1786),
.B1(n_1776),
.B2(n_1746),
.Y(n_2460)
);

AOI21xp5_ASAP7_75t_L g2461 ( 
.A1(n_1538),
.A2(n_1545),
.B(n_1555),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_1545),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_1555),
.Y(n_2463)
);

AOI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_1560),
.A2(n_1573),
.B(n_1744),
.Y(n_2464)
);

AOI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_1560),
.A2(n_1573),
.B(n_1744),
.Y(n_2465)
);

OAI21xp5_ASAP7_75t_L g2466 ( 
.A1(n_1588),
.A2(n_1656),
.B(n_1573),
.Y(n_2466)
);

AOI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_1560),
.A2(n_1706),
.B(n_1601),
.Y(n_2467)
);

OAI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_1588),
.A2(n_1601),
.B(n_1607),
.Y(n_2468)
);

O2A1O1Ixp33_ASAP7_75t_L g2469 ( 
.A1(n_1601),
.A2(n_1706),
.B(n_1607),
.C(n_1635),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_1786),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_1588),
.B(n_1607),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_L g2472 ( 
.A(n_1588),
.Y(n_2472)
);

AOI21xp5_ASAP7_75t_L g2473 ( 
.A1(n_1635),
.A2(n_1734),
.B(n_1636),
.Y(n_2473)
);

BUFx12f_ASAP7_75t_L g2474 ( 
.A(n_1588),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_1672),
.B(n_1736),
.Y(n_2475)
);

INVx4_ASAP7_75t_L g2476 ( 
.A(n_1588),
.Y(n_2476)
);

BUFx2_ASAP7_75t_L g2477 ( 
.A(n_1588),
.Y(n_2477)
);

NAND3xp33_ASAP7_75t_L g2478 ( 
.A(n_1746),
.B(n_1776),
.C(n_1704),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_1696),
.B(n_1704),
.Y(n_2479)
);

AOI21xp5_ASAP7_75t_L g2480 ( 
.A1(n_1696),
.A2(n_1706),
.B(n_1740),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_1740),
.Y(n_2481)
);

NAND3xp33_ASAP7_75t_L g2482 ( 
.A(n_1746),
.B(n_1740),
.C(n_1744),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_SL g2483 ( 
.A(n_1454),
.B(n_1931),
.Y(n_2483)
);

OAI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_1800),
.A2(n_1868),
.B1(n_1872),
.B2(n_1863),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_1768),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_1454),
.B(n_1931),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_1454),
.B(n_1427),
.Y(n_2487)
);

OAI21xp5_ASAP7_75t_L g2488 ( 
.A1(n_1931),
.A2(n_1113),
.B(n_1808),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_1454),
.B(n_1427),
.Y(n_2489)
);

AOI21xp5_ASAP7_75t_L g2490 ( 
.A1(n_1931),
.A2(n_1465),
.B(n_1113),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_L g2491 ( 
.A(n_1454),
.B(n_529),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_1429),
.Y(n_2492)
);

NOR2xp67_ASAP7_75t_L g2493 ( 
.A(n_1725),
.B(n_1465),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_1454),
.B(n_1427),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_L g2495 ( 
.A(n_1454),
.B(n_529),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_SL g2496 ( 
.A(n_1454),
.B(n_1931),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_1936),
.Y(n_2497)
);

O2A1O1Ixp33_ASAP7_75t_L g2498 ( 
.A1(n_1931),
.A2(n_1113),
.B(n_878),
.C(n_1973),
.Y(n_2498)
);

AOI21xp5_ASAP7_75t_L g2499 ( 
.A1(n_1931),
.A2(n_1465),
.B(n_1113),
.Y(n_2499)
);

OAI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_1800),
.A2(n_1868),
.B1(n_1872),
.B2(n_1863),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_1454),
.B(n_1427),
.Y(n_2501)
);

OAI21xp5_ASAP7_75t_L g2502 ( 
.A1(n_1931),
.A2(n_1113),
.B(n_1808),
.Y(n_2502)
);

OAI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_1931),
.A2(n_1113),
.B(n_878),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_1454),
.B(n_529),
.Y(n_2504)
);

A2O1A1Ixp33_ASAP7_75t_L g2505 ( 
.A1(n_1931),
.A2(n_1113),
.B(n_821),
.C(n_1800),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_1429),
.Y(n_2506)
);

OAI21xp5_ASAP7_75t_L g2507 ( 
.A1(n_1931),
.A2(n_1113),
.B(n_1808),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_1931),
.A2(n_1465),
.B(n_1113),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_R g2509 ( 
.A(n_1823),
.B(n_681),
.Y(n_2509)
);

AOI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_1800),
.A2(n_1863),
.B1(n_1872),
.B2(n_1868),
.Y(n_2510)
);

AOI22xp33_ASAP7_75t_L g2511 ( 
.A1(n_1804),
.A2(n_1858),
.B1(n_1924),
.B2(n_1914),
.Y(n_2511)
);

AND2x4_ASAP7_75t_L g2512 ( 
.A(n_1458),
.B(n_1460),
.Y(n_2512)
);

OAI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_1800),
.A2(n_1868),
.B1(n_1872),
.B2(n_1863),
.Y(n_2513)
);

INVx11_ASAP7_75t_L g2514 ( 
.A(n_1475),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_1429),
.Y(n_2515)
);

AO32x2_ASAP7_75t_L g2516 ( 
.A1(n_1808),
.A2(n_1920),
.A3(n_1693),
.B1(n_1604),
.B2(n_1597),
.Y(n_2516)
);

OR2x6_ASAP7_75t_L g2517 ( 
.A(n_1419),
.B(n_1424),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_1454),
.B(n_1427),
.Y(n_2518)
);

OAI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_1800),
.A2(n_1868),
.B1(n_1872),
.B2(n_1863),
.Y(n_2519)
);

AOI21xp5_ASAP7_75t_L g2520 ( 
.A1(n_1931),
.A2(n_1465),
.B(n_1113),
.Y(n_2520)
);

AOI21xp5_ASAP7_75t_L g2521 ( 
.A1(n_1931),
.A2(n_1465),
.B(n_1113),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_1768),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_1429),
.Y(n_2523)
);

OAI22xp5_ASAP7_75t_L g2524 ( 
.A1(n_1800),
.A2(n_1868),
.B1(n_1872),
.B2(n_1863),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_1454),
.B(n_1427),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_1454),
.B(n_1427),
.Y(n_2526)
);

AOI22xp33_ASAP7_75t_L g2527 ( 
.A1(n_1804),
.A2(n_1858),
.B1(n_1924),
.B2(n_1914),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_1768),
.Y(n_2528)
);

NAND3xp33_ASAP7_75t_L g2529 ( 
.A(n_1931),
.B(n_1113),
.C(n_1808),
.Y(n_2529)
);

A2O1A1Ixp33_ASAP7_75t_L g2530 ( 
.A1(n_1931),
.A2(n_1113),
.B(n_821),
.C(n_1800),
.Y(n_2530)
);

AOI21xp5_ASAP7_75t_L g2531 ( 
.A1(n_1931),
.A2(n_1465),
.B(n_1113),
.Y(n_2531)
);

AOI22xp33_ASAP7_75t_L g2532 ( 
.A1(n_1804),
.A2(n_1858),
.B1(n_1924),
.B2(n_1914),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_1768),
.Y(n_2533)
);

AOI21xp5_ASAP7_75t_L g2534 ( 
.A1(n_1931),
.A2(n_1465),
.B(n_1113),
.Y(n_2534)
);

AOI22xp33_ASAP7_75t_L g2535 ( 
.A1(n_1804),
.A2(n_1858),
.B1(n_1924),
.B2(n_1914),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_1454),
.B(n_1427),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_1454),
.B(n_1427),
.Y(n_2537)
);

O2A1O1Ixp33_ASAP7_75t_L g2538 ( 
.A1(n_1931),
.A2(n_1113),
.B(n_878),
.C(n_1973),
.Y(n_2538)
);

A2O1A1Ixp33_ASAP7_75t_L g2539 ( 
.A1(n_1931),
.A2(n_1113),
.B(n_821),
.C(n_1800),
.Y(n_2539)
);

BUFx12f_ASAP7_75t_L g2540 ( 
.A(n_1557),
.Y(n_2540)
);

OA21x2_ASAP7_75t_L g2541 ( 
.A1(n_1931),
.A2(n_1517),
.B(n_1525),
.Y(n_2541)
);

A2O1A1Ixp33_ASAP7_75t_L g2542 ( 
.A1(n_2505),
.A2(n_2530),
.B(n_2539),
.C(n_2538),
.Y(n_2542)
);

AOI21xp33_ASAP7_75t_L g2543 ( 
.A1(n_2498),
.A2(n_2067),
.B(n_2034),
.Y(n_2543)
);

INVxp67_ASAP7_75t_L g2544 ( 
.A(n_2198),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2180),
.B(n_2516),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2546)
);

NAND3xp33_ASAP7_75t_SL g2547 ( 
.A(n_2053),
.B(n_2035),
.C(n_2047),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_2490),
.A2(n_2508),
.B(n_2499),
.Y(n_2548)
);

BUFx6f_ASAP7_75t_L g2549 ( 
.A(n_2209),
.Y(n_2549)
);

OAI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2529),
.A2(n_2521),
.B(n_2520),
.Y(n_2550)
);

OAI21xp5_ASAP7_75t_L g2551 ( 
.A1(n_2529),
.A2(n_2534),
.B(n_2531),
.Y(n_2551)
);

OAI22x1_ASAP7_75t_L g2552 ( 
.A1(n_2011),
.A2(n_2510),
.B1(n_2050),
.B2(n_2035),
.Y(n_2552)
);

OAI21xp5_ASAP7_75t_L g2553 ( 
.A1(n_2503),
.A2(n_2502),
.B(n_2488),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2257),
.Y(n_2554)
);

AO21x1_ASAP7_75t_L g2555 ( 
.A1(n_2021),
.A2(n_2018),
.B(n_2006),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2489),
.B(n_2494),
.Y(n_2556)
);

BUFx2_ASAP7_75t_SL g2557 ( 
.A(n_2061),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2501),
.B(n_2518),
.Y(n_2558)
);

OAI21x1_ASAP7_75t_L g2559 ( 
.A1(n_2044),
.A2(n_2051),
.B(n_2071),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2525),
.B(n_2526),
.Y(n_2560)
);

AOI21xp5_ASAP7_75t_L g2561 ( 
.A1(n_2016),
.A2(n_2502),
.B(n_2488),
.Y(n_2561)
);

OAI21xp5_ASAP7_75t_L g2562 ( 
.A1(n_2507),
.A2(n_2029),
.B(n_2122),
.Y(n_2562)
);

A2O1A1Ixp33_ASAP7_75t_L g2563 ( 
.A1(n_2010),
.A2(n_2043),
.B(n_2012),
.C(n_2122),
.Y(n_2563)
);

AO31x2_ASAP7_75t_L g2564 ( 
.A1(n_2034),
.A2(n_2067),
.A3(n_2288),
.B(n_2224),
.Y(n_2564)
);

AOI21x1_ASAP7_75t_L g2565 ( 
.A1(n_2164),
.A2(n_2351),
.B(n_2324),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2536),
.B(n_2537),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2180),
.B(n_2516),
.Y(n_2567)
);

OAI21xp33_ASAP7_75t_L g2568 ( 
.A1(n_2011),
.A2(n_2510),
.B(n_2033),
.Y(n_2568)
);

CKINVDCx20_ASAP7_75t_R g2569 ( 
.A(n_2402),
.Y(n_2569)
);

CKINVDCx16_ASAP7_75t_R g2570 ( 
.A(n_2402),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_SL g2571 ( 
.A(n_2235),
.B(n_2050),
.Y(n_2571)
);

AOI21xp5_ASAP7_75t_L g2572 ( 
.A1(n_2082),
.A2(n_2213),
.B(n_2081),
.Y(n_2572)
);

AO31x2_ASAP7_75t_L g2573 ( 
.A1(n_2224),
.A2(n_2298),
.A3(n_2288),
.B(n_2484),
.Y(n_2573)
);

OAI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2033),
.A2(n_2056),
.B(n_2109),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2070),
.B(n_2079),
.Y(n_2575)
);

BUFx8_ASAP7_75t_L g2576 ( 
.A(n_2126),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2257),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_2509),
.Y(n_2578)
);

NOR2xp33_ASAP7_75t_L g2579 ( 
.A(n_2491),
.B(n_2495),
.Y(n_2579)
);

OAI21x1_ASAP7_75t_L g2580 ( 
.A1(n_2368),
.A2(n_2369),
.B(n_2127),
.Y(n_2580)
);

OR2x6_ASAP7_75t_L g2581 ( 
.A(n_2014),
.B(n_2517),
.Y(n_2581)
);

OAI21x1_ASAP7_75t_L g2582 ( 
.A1(n_2317),
.A2(n_2309),
.B(n_2308),
.Y(n_2582)
);

CKINVDCx20_ASAP7_75t_R g2583 ( 
.A(n_2039),
.Y(n_2583)
);

AO31x2_ASAP7_75t_L g2584 ( 
.A1(n_2298),
.A2(n_2513),
.A3(n_2519),
.B(n_2500),
.Y(n_2584)
);

OAI21x1_ASAP7_75t_L g2585 ( 
.A1(n_2398),
.A2(n_2297),
.B(n_2374),
.Y(n_2585)
);

AOI21xp33_ASAP7_75t_L g2586 ( 
.A1(n_2524),
.A2(n_2024),
.B(n_2002),
.Y(n_2586)
);

AOI221xp5_ASAP7_75t_SL g2587 ( 
.A1(n_2084),
.A2(n_2095),
.B1(n_2132),
.B2(n_2080),
.C(n_2089),
.Y(n_2587)
);

AOI21xp5_ASAP7_75t_L g2588 ( 
.A1(n_2213),
.A2(n_2052),
.B(n_2040),
.Y(n_2588)
);

OAI22x1_ASAP7_75t_L g2589 ( 
.A1(n_2139),
.A2(n_2152),
.B1(n_2151),
.B2(n_2242),
.Y(n_2589)
);

AOI21xp33_ASAP7_75t_L g2590 ( 
.A1(n_2002),
.A2(n_2197),
.B(n_2541),
.Y(n_2590)
);

OA22x2_ASAP7_75t_L g2591 ( 
.A1(n_2152),
.A2(n_2139),
.B1(n_2151),
.B2(n_2251),
.Y(n_2591)
);

INVx2_ASAP7_75t_SL g2592 ( 
.A(n_2287),
.Y(n_2592)
);

AOI21xp33_ASAP7_75t_L g2593 ( 
.A1(n_2197),
.A2(n_2541),
.B(n_2074),
.Y(n_2593)
);

OAI21x1_ASAP7_75t_SL g2594 ( 
.A1(n_2157),
.A2(n_2357),
.B(n_2335),
.Y(n_2594)
);

OAI21xp5_ASAP7_75t_L g2595 ( 
.A1(n_2096),
.A2(n_2148),
.B(n_2036),
.Y(n_2595)
);

AOI21x1_ASAP7_75t_L g2596 ( 
.A1(n_2164),
.A2(n_2351),
.B(n_2324),
.Y(n_2596)
);

NAND2x1p5_ASAP7_75t_L g2597 ( 
.A(n_2232),
.B(n_2476),
.Y(n_2597)
);

AO21x1_ASAP7_75t_L g2598 ( 
.A1(n_2097),
.A2(n_2108),
.B(n_2244),
.Y(n_2598)
);

OAI21x1_ASAP7_75t_L g2599 ( 
.A1(n_2192),
.A2(n_2396),
.B(n_2395),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2146),
.B(n_2060),
.Y(n_2600)
);

INVx2_ASAP7_75t_SL g2601 ( 
.A(n_2287),
.Y(n_2601)
);

O2A1O1Ixp5_ASAP7_75t_L g2602 ( 
.A1(n_2145),
.A2(n_2048),
.B(n_2083),
.C(n_2077),
.Y(n_2602)
);

AND3x4_ASAP7_75t_L g2603 ( 
.A(n_2061),
.B(n_2104),
.C(n_2240),
.Y(n_2603)
);

NAND2x1_ASAP7_75t_L g2604 ( 
.A(n_2031),
.B(n_2003),
.Y(n_2604)
);

A2O1A1Ixp33_ASAP7_75t_L g2605 ( 
.A1(n_2001),
.A2(n_2527),
.B(n_2532),
.C(n_2511),
.Y(n_2605)
);

OAI21x1_ASAP7_75t_SL g2606 ( 
.A1(n_2328),
.A2(n_2329),
.B(n_2223),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2008),
.B(n_2015),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2516),
.B(n_2088),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2257),
.Y(n_2609)
);

OAI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2504),
.A2(n_2235),
.B1(n_2535),
.B2(n_2049),
.Y(n_2610)
);

OAI22x1_ASAP7_75t_L g2611 ( 
.A1(n_2242),
.A2(n_2251),
.B1(n_2159),
.B2(n_2541),
.Y(n_2611)
);

BUFx3_ASAP7_75t_L g2612 ( 
.A(n_2126),
.Y(n_2612)
);

OAI22xp5_ASAP7_75t_L g2613 ( 
.A1(n_2090),
.A2(n_2174),
.B1(n_2183),
.B2(n_2094),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2017),
.B(n_2020),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2025),
.B(n_2028),
.Y(n_2615)
);

OAI22xp5_ASAP7_75t_L g2616 ( 
.A1(n_2094),
.A2(n_2204),
.B1(n_2470),
.B2(n_2541),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2516),
.B(n_2088),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2031),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2038),
.B(n_2042),
.Y(n_2619)
);

AO31x2_ASAP7_75t_L g2620 ( 
.A1(n_2410),
.A2(n_2145),
.A3(n_2449),
.B(n_2448),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2516),
.B(n_2144),
.Y(n_2621)
);

AOI21xp5_ASAP7_75t_L g2622 ( 
.A1(n_2158),
.A2(n_2290),
.B(n_2207),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2054),
.B(n_2062),
.Y(n_2623)
);

BUFx2_ASAP7_75t_L g2624 ( 
.A(n_2313),
.Y(n_2624)
);

OAI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_2470),
.A2(n_2169),
.B1(n_2072),
.B2(n_2143),
.Y(n_2625)
);

OAI21x1_ASAP7_75t_L g2626 ( 
.A1(n_2394),
.A2(n_2352),
.B(n_2349),
.Y(n_2626)
);

OA21x2_ASAP7_75t_L g2627 ( 
.A1(n_2452),
.A2(n_2466),
.B(n_2468),
.Y(n_2627)
);

OAI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2165),
.A2(n_2130),
.B(n_2091),
.Y(n_2628)
);

OAI21x1_ASAP7_75t_SL g2629 ( 
.A1(n_2220),
.A2(n_2187),
.B(n_2181),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2026),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2026),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2057),
.Y(n_2632)
);

A2O1A1Ixp33_ASAP7_75t_L g2633 ( 
.A1(n_2163),
.A2(n_2160),
.B(n_2379),
.C(n_2170),
.Y(n_2633)
);

AOI21xp5_ASAP7_75t_L g2634 ( 
.A1(n_2290),
.A2(n_2493),
.B(n_2327),
.Y(n_2634)
);

OAI21x1_ASAP7_75t_L g2635 ( 
.A1(n_2119),
.A2(n_2231),
.B(n_2443),
.Y(n_2635)
);

INVx3_ASAP7_75t_L g2636 ( 
.A(n_2031),
.Y(n_2636)
);

AO31x2_ASAP7_75t_L g2637 ( 
.A1(n_2410),
.A2(n_2458),
.A3(n_2457),
.B(n_2275),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2144),
.B(n_2359),
.Y(n_2638)
);

AND3x4_ASAP7_75t_L g2639 ( 
.A(n_2104),
.B(n_2240),
.C(n_2172),
.Y(n_2639)
);

INVx1_ASAP7_75t_SL g2640 ( 
.A(n_2313),
.Y(n_2640)
);

AND2x2_ASAP7_75t_SL g2641 ( 
.A(n_2283),
.B(n_2316),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_SL g2642 ( 
.A(n_2474),
.B(n_2055),
.Y(n_2642)
);

OAI21x1_ASAP7_75t_L g2643 ( 
.A1(n_2231),
.A2(n_2086),
.B(n_2129),
.Y(n_2643)
);

OAI21x1_ASAP7_75t_L g2644 ( 
.A1(n_2231),
.A2(n_2086),
.B(n_2147),
.Y(n_2644)
);

OAI21x1_ASAP7_75t_L g2645 ( 
.A1(n_2086),
.A2(n_2125),
.B(n_2073),
.Y(n_2645)
);

INVx6_ASAP7_75t_L g2646 ( 
.A(n_2366),
.Y(n_2646)
);

A2O1A1Ixp33_ASAP7_75t_L g2647 ( 
.A1(n_2379),
.A2(n_2170),
.B(n_2159),
.C(n_2226),
.Y(n_2647)
);

AOI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_2282),
.A2(n_2284),
.B(n_2281),
.Y(n_2648)
);

AOI21x1_ASAP7_75t_L g2649 ( 
.A1(n_2273),
.A2(n_2311),
.B(n_2300),
.Y(n_2649)
);

AOI21xp5_ASAP7_75t_L g2650 ( 
.A1(n_2423),
.A2(n_2227),
.B(n_2136),
.Y(n_2650)
);

AND2x4_ASAP7_75t_L g2651 ( 
.A(n_2232),
.B(n_2477),
.Y(n_2651)
);

AOI21xp33_ASAP7_75t_L g2652 ( 
.A1(n_2433),
.A2(n_2453),
.B(n_2451),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2065),
.B(n_2068),
.Y(n_2653)
);

BUFx6f_ASAP7_75t_SL g2654 ( 
.A(n_2066),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2150),
.B(n_2149),
.Y(n_2655)
);

OAI21x1_ASAP7_75t_L g2656 ( 
.A1(n_2073),
.A2(n_2391),
.B(n_2211),
.Y(n_2656)
);

AOI21xp5_ASAP7_75t_L g2657 ( 
.A1(n_2423),
.A2(n_2264),
.B(n_2255),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_2066),
.B(n_2039),
.Y(n_2658)
);

OAI21x1_ASAP7_75t_L g2659 ( 
.A1(n_2073),
.A2(n_2391),
.B(n_2418),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2100),
.B(n_2103),
.Y(n_2660)
);

AOI21xp5_ASAP7_75t_L g2661 ( 
.A1(n_2330),
.A2(n_2334),
.B(n_2331),
.Y(n_2661)
);

INVx3_ASAP7_75t_L g2662 ( 
.A(n_2225),
.Y(n_2662)
);

AOI21xp5_ASAP7_75t_L g2663 ( 
.A1(n_2175),
.A2(n_2177),
.B(n_2341),
.Y(n_2663)
);

INVx3_ASAP7_75t_L g2664 ( 
.A(n_2225),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2105),
.B(n_2085),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2384),
.Y(n_2666)
);

AOI21xp33_ASAP7_75t_L g2667 ( 
.A1(n_2199),
.A2(n_2419),
.B(n_2431),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2057),
.Y(n_2668)
);

NAND2x1p5_ASAP7_75t_L g2669 ( 
.A(n_2232),
.B(n_2476),
.Y(n_2669)
);

BUFx6f_ASAP7_75t_L g2670 ( 
.A(n_2209),
.Y(n_2670)
);

NAND3xp33_ASAP7_75t_SL g2671 ( 
.A(n_2140),
.B(n_2190),
.C(n_2168),
.Y(n_2671)
);

OR2x6_ASAP7_75t_L g2672 ( 
.A(n_2014),
.B(n_2517),
.Y(n_2672)
);

INVxp67_ASAP7_75t_L g2673 ( 
.A(n_2037),
.Y(n_2673)
);

OAI21x1_ASAP7_75t_L g2674 ( 
.A1(n_2171),
.A2(n_2424),
.B(n_2185),
.Y(n_2674)
);

AOI21xp5_ASAP7_75t_L g2675 ( 
.A1(n_2093),
.A2(n_2154),
.B(n_2442),
.Y(n_2675)
);

A2O1A1Ixp33_ASAP7_75t_L g2676 ( 
.A1(n_2226),
.A2(n_2245),
.B(n_2272),
.C(n_2206),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2041),
.B(n_2124),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2128),
.B(n_2098),
.Y(n_2678)
);

AOI22xp5_ASAP7_75t_L g2679 ( 
.A1(n_2200),
.A2(n_2414),
.B1(n_2064),
.B2(n_2167),
.Y(n_2679)
);

A2O1A1Ixp33_ASAP7_75t_L g2680 ( 
.A1(n_2256),
.A2(n_2320),
.B(n_2323),
.C(n_2278),
.Y(n_2680)
);

NAND2xp33_ASAP7_75t_L g2681 ( 
.A(n_2237),
.B(n_2460),
.Y(n_2681)
);

OAI21x1_ASAP7_75t_L g2682 ( 
.A1(n_2171),
.A2(n_2185),
.B(n_2208),
.Y(n_2682)
);

BUFx3_ASAP7_75t_L g2683 ( 
.A(n_2289),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2107),
.B(n_2110),
.Y(n_2684)
);

AOI21xp5_ASAP7_75t_L g2685 ( 
.A1(n_2093),
.A2(n_2166),
.B(n_2055),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2359),
.B(n_2399),
.Y(n_2686)
);

OR2x2_ASAP7_75t_L g2687 ( 
.A(n_2131),
.B(n_2370),
.Y(n_2687)
);

NAND2x1p5_ASAP7_75t_L g2688 ( 
.A(n_2232),
.B(n_2476),
.Y(n_2688)
);

INVx5_ASAP7_75t_L g2689 ( 
.A(n_2474),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2113),
.B(n_2117),
.Y(n_2690)
);

OAI21x1_ASAP7_75t_L g2691 ( 
.A1(n_2208),
.A2(n_2428),
.B(n_2228),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2118),
.B(n_2123),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2009),
.B(n_2142),
.Y(n_2693)
);

OR2x6_ASAP7_75t_L g2694 ( 
.A(n_2014),
.B(n_2517),
.Y(n_2694)
);

OAI21x1_ASAP7_75t_L g2695 ( 
.A1(n_2428),
.A2(n_2228),
.B(n_2292),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2485),
.Y(n_2696)
);

INVx2_ASAP7_75t_SL g2697 ( 
.A(n_2403),
.Y(n_2697)
);

INVx6_ASAP7_75t_L g2698 ( 
.A(n_2366),
.Y(n_2698)
);

AOI21xp33_ASAP7_75t_L g2699 ( 
.A1(n_2194),
.A2(n_2426),
.B(n_2135),
.Y(n_2699)
);

OAI21x1_ASAP7_75t_L g2700 ( 
.A1(n_2428),
.A2(n_2292),
.B(n_2176),
.Y(n_2700)
);

AOI21x1_ASAP7_75t_SL g2701 ( 
.A1(n_2205),
.A2(n_2239),
.B(n_2168),
.Y(n_2701)
);

OAI21x1_ASAP7_75t_L g2702 ( 
.A1(n_2176),
.A2(n_2407),
.B(n_2444),
.Y(n_2702)
);

AOI21xp5_ASAP7_75t_L g2703 ( 
.A1(n_2093),
.A2(n_2354),
.B(n_2454),
.Y(n_2703)
);

OAI21x1_ASAP7_75t_SL g2704 ( 
.A1(n_2401),
.A2(n_2460),
.B(n_2263),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2196),
.B(n_2111),
.Y(n_2705)
);

AO21x2_ASAP7_75t_L g2706 ( 
.A1(n_2455),
.A2(n_2464),
.B(n_2461),
.Y(n_2706)
);

OAI21xp33_ASAP7_75t_L g2707 ( 
.A1(n_2261),
.A2(n_2294),
.B(n_2246),
.Y(n_2707)
);

AND2x4_ASAP7_75t_L g2708 ( 
.A(n_2232),
.B(n_2477),
.Y(n_2708)
);

AO21x1_ASAP7_75t_L g2709 ( 
.A1(n_2253),
.A2(n_2268),
.B(n_2087),
.Y(n_2709)
);

AOI21x1_ASAP7_75t_SL g2710 ( 
.A1(n_2193),
.A2(n_2195),
.B(n_2143),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2399),
.B(n_2114),
.Y(n_2711)
);

AOI21xp5_ASAP7_75t_L g2712 ( 
.A1(n_2093),
.A2(n_2354),
.B(n_2347),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_L g2713 ( 
.A(n_2066),
.B(n_2200),
.Y(n_2713)
);

AOI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2345),
.A2(n_2254),
.B(n_2137),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2485),
.Y(n_2715)
);

AOI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2106),
.A2(n_2210),
.B(n_2137),
.Y(n_2716)
);

CKINVDCx8_ASAP7_75t_R g2717 ( 
.A(n_2400),
.Y(n_2717)
);

OA21x2_ASAP7_75t_L g2718 ( 
.A1(n_2466),
.A2(n_2468),
.B(n_2338),
.Y(n_2718)
);

AOI21xp5_ASAP7_75t_L g2719 ( 
.A1(n_2106),
.A2(n_2210),
.B(n_2137),
.Y(n_2719)
);

OAI21x1_ASAP7_75t_L g2720 ( 
.A1(n_2176),
.A2(n_2215),
.B(n_2212),
.Y(n_2720)
);

A2O1A1Ixp33_ASAP7_75t_L g2721 ( 
.A1(n_2482),
.A2(n_2271),
.B(n_2346),
.C(n_2155),
.Y(n_2721)
);

OAI22xp33_ASAP7_75t_L g2722 ( 
.A1(n_2260),
.A2(n_2263),
.B1(n_2408),
.B2(n_2289),
.Y(n_2722)
);

INVx1_ASAP7_75t_SL g2723 ( 
.A(n_2370),
.Y(n_2723)
);

NAND2x1p5_ASAP7_75t_L g2724 ( 
.A(n_2279),
.B(n_2386),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2412),
.Y(n_2725)
);

AOI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2106),
.A2(n_2210),
.B(n_2432),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2114),
.B(n_2522),
.Y(n_2727)
);

INVx2_ASAP7_75t_SL g2728 ( 
.A(n_2363),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2413),
.Y(n_2729)
);

AOI21xp5_ASAP7_75t_L g2730 ( 
.A1(n_2415),
.A2(n_2427),
.B(n_2273),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_SL g2731 ( 
.A(n_2414),
.B(n_2214),
.Y(n_2731)
);

OAI21x1_ASAP7_75t_L g2732 ( 
.A1(n_2372),
.A2(n_2248),
.B(n_2225),
.Y(n_2732)
);

OAI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2246),
.A2(n_2326),
.B(n_2346),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2112),
.B(n_2173),
.Y(n_2734)
);

OAI21x1_ASAP7_75t_L g2735 ( 
.A1(n_2248),
.A2(n_2383),
.B(n_2382),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2522),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2528),
.Y(n_2737)
);

INVx5_ASAP7_75t_L g2738 ( 
.A(n_2472),
.Y(n_2738)
);

OAI21xp5_ASAP7_75t_L g2739 ( 
.A1(n_2059),
.A2(n_2405),
.B(n_2087),
.Y(n_2739)
);

NOR2xp67_ASAP7_75t_L g2740 ( 
.A(n_2279),
.B(n_2386),
.Y(n_2740)
);

INVx4_ASAP7_75t_L g2741 ( 
.A(n_2116),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2059),
.Y(n_2742)
);

AOI21xp5_ASAP7_75t_L g2743 ( 
.A1(n_2404),
.A2(n_2478),
.B(n_2377),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2380),
.B(n_2249),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2528),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2234),
.B(n_2243),
.Y(n_2746)
);

AOI21xp5_ASAP7_75t_L g2747 ( 
.A1(n_2478),
.A2(n_2377),
.B(n_2375),
.Y(n_2747)
);

OAI21x1_ASAP7_75t_L g2748 ( 
.A1(n_2248),
.A2(n_2390),
.B(n_2425),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2258),
.B(n_2262),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2533),
.B(n_2101),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_SL g2751 ( 
.A(n_2217),
.B(n_2447),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2189),
.B(n_2182),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2364),
.B(n_2367),
.Y(n_2753)
);

OAI21x1_ASAP7_75t_L g2754 ( 
.A1(n_2425),
.A2(n_2373),
.B(n_2430),
.Y(n_2754)
);

OR2x6_ASAP7_75t_L g2755 ( 
.A(n_2014),
.B(n_2517),
.Y(n_2755)
);

OAI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2219),
.A2(n_2161),
.B(n_2247),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2533),
.B(n_2101),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2138),
.B(n_2153),
.Y(n_2758)
);

AO31x2_ASAP7_75t_L g2759 ( 
.A1(n_2307),
.A2(n_2467),
.A3(n_2473),
.B(n_2465),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2376),
.B(n_2387),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2138),
.B(n_2153),
.Y(n_2761)
);

INVx2_ASAP7_75t_SL g2762 ( 
.A(n_2400),
.Y(n_2762)
);

OAI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_2229),
.A2(n_2319),
.B(n_2482),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2191),
.Y(n_2764)
);

INVx1_ASAP7_75t_SL g2765 ( 
.A(n_2375),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2392),
.B(n_2393),
.Y(n_2766)
);

AOI21x1_ASAP7_75t_L g2767 ( 
.A1(n_2092),
.A2(n_2121),
.B(n_2099),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2413),
.Y(n_2768)
);

AO31x2_ASAP7_75t_L g2769 ( 
.A1(n_2480),
.A2(n_2238),
.A3(n_2007),
.B(n_2523),
.Y(n_2769)
);

OAI21x1_ASAP7_75t_L g2770 ( 
.A1(n_2469),
.A2(n_2092),
.B(n_2420),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2397),
.B(n_2406),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2421),
.B(n_2381),
.Y(n_2772)
);

OAI21x1_ASAP7_75t_L g2773 ( 
.A1(n_2420),
.A2(n_2435),
.B(n_2411),
.Y(n_2773)
);

OAI21x1_ASAP7_75t_L g2774 ( 
.A1(n_2420),
.A2(n_2411),
.B(n_2222),
.Y(n_2774)
);

OAI21xp33_ASAP7_75t_L g2775 ( 
.A1(n_2294),
.A2(n_2229),
.B(n_2201),
.Y(n_2775)
);

BUFx2_ASAP7_75t_L g2776 ( 
.A(n_2301),
.Y(n_2776)
);

BUFx6f_ASAP7_75t_SL g2777 ( 
.A(n_2438),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2188),
.B(n_2230),
.Y(n_2778)
);

AOI21xp5_ASAP7_75t_L g2779 ( 
.A1(n_2030),
.A2(n_2202),
.B(n_2186),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2188),
.B(n_2230),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2250),
.Y(n_2781)
);

AO31x2_ASAP7_75t_L g2782 ( 
.A1(n_2007),
.A2(n_2388),
.A3(n_2523),
.B(n_2019),
.Y(n_2782)
);

O2A1O1Ixp5_ASAP7_75t_L g2783 ( 
.A1(n_2441),
.A2(n_2115),
.B(n_2134),
.C(n_2133),
.Y(n_2783)
);

BUFx3_ASAP7_75t_L g2784 ( 
.A(n_2184),
.Y(n_2784)
);

OAI21x1_ASAP7_75t_L g2785 ( 
.A1(n_2411),
.A2(n_2361),
.B(n_2416),
.Y(n_2785)
);

AOI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_2030),
.A2(n_2202),
.B(n_2186),
.Y(n_2786)
);

OAI21xp33_ASAP7_75t_SL g2787 ( 
.A1(n_2260),
.A2(n_2447),
.B(n_2201),
.Y(n_2787)
);

OAI21xp5_ASAP7_75t_L g2788 ( 
.A1(n_2389),
.A2(n_2322),
.B(n_2293),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2233),
.B(n_2241),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2233),
.B(n_2241),
.Y(n_2790)
);

OAI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2322),
.A2(n_2350),
.B(n_2355),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2191),
.Y(n_2792)
);

OAI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2120),
.A2(n_2141),
.B(n_2409),
.Y(n_2793)
);

OAI21x1_ASAP7_75t_SL g2794 ( 
.A1(n_2422),
.A2(n_2445),
.B(n_2408),
.Y(n_2794)
);

AOI221xp5_ASAP7_75t_L g2795 ( 
.A1(n_2216),
.A2(n_2299),
.B1(n_2236),
.B2(n_2342),
.C(n_2312),
.Y(n_2795)
);

AOI21xp33_ASAP7_75t_L g2796 ( 
.A1(n_2203),
.A2(n_2221),
.B(n_2416),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2259),
.B(n_2266),
.Y(n_2797)
);

AOI21xp5_ASAP7_75t_L g2798 ( 
.A1(n_2277),
.A2(n_2512),
.B(n_2332),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2019),
.Y(n_2799)
);

NAND2x1p5_ASAP7_75t_L g2800 ( 
.A(n_2279),
.B(n_2386),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2216),
.Y(n_2801)
);

AOI21x1_ASAP7_75t_L g2802 ( 
.A1(n_2378),
.A2(n_2299),
.B(n_2236),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2259),
.B(n_2266),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2269),
.B(n_2303),
.Y(n_2804)
);

AOI21xp5_ASAP7_75t_L g2805 ( 
.A1(n_2277),
.A2(n_2332),
.B(n_2512),
.Y(n_2805)
);

NOR2x1_ASAP7_75t_L g2806 ( 
.A(n_2252),
.B(n_2267),
.Y(n_2806)
);

CKINVDCx5p33_ASAP7_75t_R g2807 ( 
.A(n_2027),
.Y(n_2807)
);

OR2x2_ASAP7_75t_L g2808 ( 
.A(n_2131),
.B(n_2301),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2312),
.B(n_2342),
.Y(n_2809)
);

BUFx12f_ASAP7_75t_L g2810 ( 
.A(n_2023),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_2023),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2353),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2358),
.B(n_2269),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2472),
.B(n_2279),
.Y(n_2814)
);

NOR2x1_ASAP7_75t_L g2815 ( 
.A(n_2270),
.B(n_2422),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2434),
.Y(n_2816)
);

BUFx3_ASAP7_75t_L g2817 ( 
.A(n_2184),
.Y(n_2817)
);

NAND2x1_ASAP7_75t_L g2818 ( 
.A(n_2003),
.B(n_2102),
.Y(n_2818)
);

AOI21xp5_ASAP7_75t_L g2819 ( 
.A1(n_2277),
.A2(n_2332),
.B(n_2512),
.Y(n_2819)
);

INVx1_ASAP7_75t_SL g2820 ( 
.A(n_2439),
.Y(n_2820)
);

NOR2xp33_ASAP7_75t_L g2821 ( 
.A(n_2497),
.B(n_2046),
.Y(n_2821)
);

INVxp67_ASAP7_75t_L g2822 ( 
.A(n_2265),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2022),
.Y(n_2823)
);

OR2x2_ASAP7_75t_L g2824 ( 
.A(n_2295),
.B(n_2360),
.Y(n_2824)
);

INVx3_ASAP7_75t_L g2825 ( 
.A(n_2472),
.Y(n_2825)
);

NAND2x1_ASAP7_75t_L g2826 ( 
.A(n_2003),
.B(n_2102),
.Y(n_2826)
);

AOI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2447),
.A2(n_2365),
.B(n_2302),
.Y(n_2827)
);

AO31x2_ASAP7_75t_L g2828 ( 
.A1(n_2022),
.A2(n_2325),
.A3(n_2515),
.B(n_2045),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2303),
.B(n_2291),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2295),
.B(n_2434),
.Y(n_2830)
);

AOI221x1_ASAP7_75t_L g2831 ( 
.A1(n_2437),
.A2(n_2475),
.B1(n_2479),
.B2(n_2318),
.C(n_2339),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2296),
.B(n_2315),
.Y(n_2832)
);

OAI21xp33_ASAP7_75t_L g2833 ( 
.A1(n_2417),
.A2(n_2497),
.B(n_2280),
.Y(n_2833)
);

OAI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2102),
.A2(n_2305),
.B(n_2178),
.Y(n_2834)
);

OAI22x1_ASAP7_75t_L g2835 ( 
.A1(n_2279),
.A2(n_2386),
.B1(n_2439),
.B2(n_2471),
.Y(n_2835)
);

NAND2x1_ASAP7_75t_L g2836 ( 
.A(n_2003),
.B(n_2162),
.Y(n_2836)
);

CKINVDCx8_ASAP7_75t_R g2837 ( 
.A(n_2438),
.Y(n_2837)
);

INVx3_ASAP7_75t_L g2838 ( 
.A(n_2472),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2274),
.B(n_2276),
.Y(n_2839)
);

OAI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2445),
.A2(n_2179),
.B(n_2305),
.Y(n_2840)
);

NAND2x1p5_ASAP7_75t_L g2841 ( 
.A(n_2386),
.B(n_2472),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2440),
.Y(n_2842)
);

OAI21xp5_ASAP7_75t_L g2843 ( 
.A1(n_2162),
.A2(n_2302),
.B(n_2178),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2440),
.Y(n_2844)
);

OAI21x1_ASAP7_75t_SL g2845 ( 
.A1(n_2162),
.A2(n_2178),
.B(n_2302),
.Y(n_2845)
);

INVx2_ASAP7_75t_SL g2846 ( 
.A(n_2116),
.Y(n_2846)
);

OAI21x1_ASAP7_75t_L g2847 ( 
.A1(n_2285),
.A2(n_2336),
.B(n_2337),
.Y(n_2847)
);

AO21x2_ASAP7_75t_L g2848 ( 
.A1(n_2156),
.A2(n_2218),
.B(n_2515),
.Y(n_2848)
);

OA21x2_ASAP7_75t_L g2849 ( 
.A1(n_2450),
.A2(n_2333),
.B(n_2314),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2286),
.B(n_2304),
.Y(n_2850)
);

OAI21xp5_ASAP7_75t_L g2851 ( 
.A1(n_2305),
.A2(n_2371),
.B(n_2310),
.Y(n_2851)
);

INVxp67_ASAP7_75t_SL g2852 ( 
.A(n_2063),
.Y(n_2852)
);

OAI21x1_ASAP7_75t_L g2853 ( 
.A1(n_2063),
.A2(n_2436),
.B(n_2506),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2456),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2456),
.B(n_2459),
.Y(n_2855)
);

AOI21xp5_ASAP7_75t_L g2856 ( 
.A1(n_2321),
.A2(n_2348),
.B(n_2344),
.Y(n_2856)
);

OAI21x1_ASAP7_75t_L g2857 ( 
.A1(n_2069),
.A2(n_2306),
.B(n_2492),
.Y(n_2857)
);

AOI21x1_ASAP7_75t_L g2858 ( 
.A1(n_2471),
.A2(n_2459),
.B(n_2492),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2362),
.B(n_2438),
.Y(n_2859)
);

OAI21x1_ASAP7_75t_L g2860 ( 
.A1(n_2069),
.A2(n_2343),
.B(n_2481),
.Y(n_2860)
);

OAI21x1_ASAP7_75t_L g2861 ( 
.A1(n_2075),
.A2(n_2343),
.B(n_2463),
.Y(n_2861)
);

OAI22xp5_ASAP7_75t_L g2862 ( 
.A1(n_2179),
.A2(n_2514),
.B1(n_2438),
.B2(n_2058),
.Y(n_2862)
);

O2A1O1Ixp5_ASAP7_75t_L g2863 ( 
.A1(n_2471),
.A2(n_2340),
.B(n_2429),
.C(n_2463),
.Y(n_2863)
);

AOI21xp5_ASAP7_75t_L g2864 ( 
.A1(n_2058),
.A2(n_2076),
.B(n_2356),
.Y(n_2864)
);

AOI22xp33_ASAP7_75t_L g2865 ( 
.A1(n_2003),
.A2(n_2325),
.B1(n_2462),
.B2(n_2429),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2184),
.B(n_2003),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2003),
.B(n_2340),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_2078),
.B(n_2385),
.Y(n_2868)
);

OAI22xp5_ASAP7_75t_L g2869 ( 
.A1(n_2514),
.A2(n_2013),
.B1(n_2540),
.B2(n_2046),
.Y(n_2869)
);

BUFx2_ASAP7_75t_L g2870 ( 
.A(n_2366),
.Y(n_2870)
);

OAI21x1_ASAP7_75t_L g2871 ( 
.A1(n_2446),
.A2(n_2013),
.B(n_2540),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2446),
.B(n_2004),
.Y(n_2872)
);

OAI22xp5_ASAP7_75t_L g2873 ( 
.A1(n_2035),
.A2(n_1800),
.B1(n_1868),
.B2(n_1863),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2874)
);

OAI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2875)
);

AOI21x1_ASAP7_75t_L g2876 ( 
.A1(n_2044),
.A2(n_2005),
.B(n_2490),
.Y(n_2876)
);

OAI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2035),
.A2(n_1800),
.B1(n_1868),
.B2(n_1863),
.Y(n_2877)
);

AOI21xp33_ASAP7_75t_L g2878 ( 
.A1(n_2498),
.A2(n_1931),
.B(n_1113),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2180),
.B(n_2516),
.Y(n_2879)
);

AND2x2_ASAP7_75t_L g2880 ( 
.A(n_2180),
.B(n_2516),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2257),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_SL g2882 ( 
.A(n_2235),
.B(n_2035),
.Y(n_2882)
);

AOI21xp5_ASAP7_75t_L g2883 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2883)
);

AOI21xp5_ASAP7_75t_L g2884 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2884)
);

INVx2_ASAP7_75t_SL g2885 ( 
.A(n_2287),
.Y(n_2885)
);

BUFx3_ASAP7_75t_L g2886 ( 
.A(n_2126),
.Y(n_2886)
);

NOR2x1_ASAP7_75t_L g2887 ( 
.A(n_2084),
.B(n_2529),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2888)
);

OAI21xp33_ASAP7_75t_SL g2889 ( 
.A1(n_2488),
.A2(n_1931),
.B(n_2502),
.Y(n_2889)
);

BUFx3_ASAP7_75t_L g2890 ( 
.A(n_2126),
.Y(n_2890)
);

A2O1A1Ixp33_ASAP7_75t_L g2891 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.C(n_2530),
.Y(n_2891)
);

INVx2_ASAP7_75t_SL g2892 ( 
.A(n_2287),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2257),
.Y(n_2894)
);

BUFx3_ASAP7_75t_L g2895 ( 
.A(n_2126),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2180),
.B(n_2516),
.Y(n_2896)
);

AOI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2897)
);

OAI21xp5_ASAP7_75t_L g2898 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2898)
);

NAND2x1p5_ASAP7_75t_L g2899 ( 
.A(n_2232),
.B(n_1725),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2900)
);

AOI21xp5_ASAP7_75t_L g2901 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2901)
);

O2A1O1Ixp33_ASAP7_75t_SL g2902 ( 
.A1(n_2029),
.A2(n_2486),
.B(n_2496),
.C(n_2483),
.Y(n_2902)
);

OAI21x1_ASAP7_75t_SL g2903 ( 
.A1(n_2012),
.A2(n_2502),
.B(n_2488),
.Y(n_2903)
);

HB1xp67_ASAP7_75t_L g2904 ( 
.A(n_2009),
.Y(n_2904)
);

BUFx4f_ASAP7_75t_L g2905 ( 
.A(n_2126),
.Y(n_2905)
);

AOI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2257),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2257),
.Y(n_2908)
);

INVxp67_ASAP7_75t_SL g2909 ( 
.A(n_2423),
.Y(n_2909)
);

OAI21x1_ASAP7_75t_SL g2910 ( 
.A1(n_2012),
.A2(n_2502),
.B(n_2488),
.Y(n_2910)
);

AOI21xp5_ASAP7_75t_L g2911 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2911)
);

NAND2x1_ASAP7_75t_L g2912 ( 
.A(n_2031),
.B(n_2032),
.Y(n_2912)
);

AOI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2913)
);

NOR2x1_ASAP7_75t_SL g2914 ( 
.A(n_2474),
.B(n_2014),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2915)
);

OAI21x1_ASAP7_75t_SL g2916 ( 
.A1(n_2012),
.A2(n_2502),
.B(n_2488),
.Y(n_2916)
);

AOI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2257),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2920)
);

INVx3_ASAP7_75t_L g2921 ( 
.A(n_2031),
.Y(n_2921)
);

A2O1A1Ixp33_ASAP7_75t_L g2922 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.C(n_2530),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2923)
);

NAND2xp33_ASAP7_75t_L g2924 ( 
.A(n_2505),
.B(n_1931),
.Y(n_2924)
);

INVx3_ASAP7_75t_L g2925 ( 
.A(n_2031),
.Y(n_2925)
);

AOI21xp5_ASAP7_75t_L g2926 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2926)
);

AOI21x1_ASAP7_75t_SL g2927 ( 
.A1(n_2004),
.A2(n_969),
.B(n_962),
.Y(n_2927)
);

O2A1O1Ixp33_ASAP7_75t_L g2928 ( 
.A1(n_2503),
.A2(n_1113),
.B(n_1931),
.C(n_1996),
.Y(n_2928)
);

OAI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.Y(n_2929)
);

BUFx2_ASAP7_75t_L g2930 ( 
.A(n_2287),
.Y(n_2930)
);

AOI21xp5_ASAP7_75t_L g2931 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2934)
);

OR2x2_ASAP7_75t_L g2935 ( 
.A(n_2131),
.B(n_2370),
.Y(n_2935)
);

BUFx3_ASAP7_75t_L g2936 ( 
.A(n_2126),
.Y(n_2936)
);

INVx2_ASAP7_75t_SL g2937 ( 
.A(n_2287),
.Y(n_2937)
);

NAND2x1_ASAP7_75t_L g2938 ( 
.A(n_2031),
.B(n_2032),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2939)
);

AO31x2_ASAP7_75t_L g2940 ( 
.A1(n_2505),
.A2(n_2539),
.A3(n_2530),
.B(n_2034),
.Y(n_2940)
);

OAI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2035),
.A2(n_1800),
.B1(n_1868),
.B2(n_1863),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2942)
);

NOR2xp33_ASAP7_75t_L g2943 ( 
.A(n_2491),
.B(n_529),
.Y(n_2943)
);

NAND2x1p5_ASAP7_75t_L g2944 ( 
.A(n_2232),
.B(n_1725),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_2235),
.B(n_2035),
.Y(n_2946)
);

CKINVDCx5p33_ASAP7_75t_R g2947 ( 
.A(n_2509),
.Y(n_2947)
);

OAI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2180),
.B(n_2516),
.Y(n_2949)
);

A2O1A1Ixp33_ASAP7_75t_L g2950 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.C(n_2530),
.Y(n_2950)
);

OAI22x1_ASAP7_75t_L g2951 ( 
.A1(n_2011),
.A2(n_2510),
.B1(n_2050),
.B2(n_2035),
.Y(n_2951)
);

OAI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.Y(n_2952)
);

BUFx4f_ASAP7_75t_L g2953 ( 
.A(n_2126),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2257),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2257),
.Y(n_2955)
);

OAI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2957)
);

O2A1O1Ixp5_ASAP7_75t_L g2958 ( 
.A1(n_2488),
.A2(n_1931),
.B(n_2507),
.C(n_2502),
.Y(n_2958)
);

AOI21x1_ASAP7_75t_L g2959 ( 
.A1(n_2044),
.A2(n_2005),
.B(n_2490),
.Y(n_2959)
);

NOR2xp33_ASAP7_75t_L g2960 ( 
.A(n_2491),
.B(n_529),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2961)
);

AO31x2_ASAP7_75t_L g2962 ( 
.A1(n_2505),
.A2(n_2539),
.A3(n_2530),
.B(n_2034),
.Y(n_2962)
);

NOR2xp33_ASAP7_75t_L g2963 ( 
.A(n_2491),
.B(n_529),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2180),
.B(n_2516),
.Y(n_2964)
);

AOI21xp5_ASAP7_75t_L g2965 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2965)
);

OAI21xp5_ASAP7_75t_SL g2966 ( 
.A1(n_2035),
.A2(n_1863),
.B(n_1800),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2968)
);

AOI22xp5_ASAP7_75t_L g2969 ( 
.A1(n_2021),
.A2(n_1800),
.B1(n_1868),
.B2(n_1863),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2257),
.Y(n_2970)
);

OAI21xp5_ASAP7_75t_L g2971 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_2180),
.B(n_2516),
.Y(n_2974)
);

BUFx6f_ASAP7_75t_L g2975 ( 
.A(n_2209),
.Y(n_2975)
);

OAI21xp5_ASAP7_75t_L g2976 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2257),
.Y(n_2977)
);

AOI21xp5_ASAP7_75t_L g2978 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2180),
.B(n_2516),
.Y(n_2979)
);

OAI21xp5_ASAP7_75t_L g2980 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2980)
);

A2O1A1Ixp33_ASAP7_75t_L g2981 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.C(n_2530),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2983)
);

NOR2x1_ASAP7_75t_L g2984 ( 
.A(n_2084),
.B(n_2529),
.Y(n_2984)
);

AOI21xp5_ASAP7_75t_L g2985 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2985)
);

BUFx8_ASAP7_75t_SL g2986 ( 
.A(n_2402),
.Y(n_2986)
);

A2O1A1Ixp33_ASAP7_75t_L g2987 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.C(n_2530),
.Y(n_2987)
);

AOI21x1_ASAP7_75t_L g2988 ( 
.A1(n_2044),
.A2(n_2005),
.B(n_2490),
.Y(n_2988)
);

OR2x6_ASAP7_75t_L g2989 ( 
.A(n_2014),
.B(n_2517),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2004),
.B(n_2487),
.Y(n_2990)
);

AOI221x1_ASAP7_75t_L g2991 ( 
.A1(n_2505),
.A2(n_1931),
.B1(n_2530),
.B2(n_2539),
.C(n_1113),
.Y(n_2991)
);

AOI21xp5_ASAP7_75t_L g2992 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2992)
);

BUFx3_ASAP7_75t_L g2993 ( 
.A(n_2126),
.Y(n_2993)
);

AOI21xp5_ASAP7_75t_L g2994 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2994)
);

OAI22xp5_ASAP7_75t_SL g2995 ( 
.A1(n_2402),
.A2(n_2151),
.B1(n_2035),
.B2(n_2529),
.Y(n_2995)
);

NOR2xp33_ASAP7_75t_L g2996 ( 
.A(n_2491),
.B(n_529),
.Y(n_2996)
);

OAI21xp5_ASAP7_75t_L g2997 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_2997)
);

NOR2xp67_ASAP7_75t_L g2998 ( 
.A(n_2232),
.B(n_2474),
.Y(n_2998)
);

NOR2xp33_ASAP7_75t_L g2999 ( 
.A(n_2491),
.B(n_529),
.Y(n_2999)
);

AOI21xp33_ASAP7_75t_L g3000 ( 
.A1(n_2498),
.A2(n_1931),
.B(n_1113),
.Y(n_3000)
);

OAI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2035),
.A2(n_1800),
.B1(n_1868),
.B2(n_1863),
.Y(n_3001)
);

AOI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_SL g3003 ( 
.A(n_2235),
.B(n_2035),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2004),
.B(n_2487),
.Y(n_3004)
);

AOI21xp5_ASAP7_75t_L g3005 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_3005)
);

AOI21xp33_ASAP7_75t_L g3006 ( 
.A1(n_2498),
.A2(n_1931),
.B(n_1113),
.Y(n_3006)
);

AOI21xp5_ASAP7_75t_L g3007 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2180),
.B(n_2516),
.Y(n_3008)
);

A2O1A1Ixp33_ASAP7_75t_L g3009 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.C(n_2530),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2004),
.B(n_2487),
.Y(n_3010)
);

OAI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_2530),
.Y(n_3011)
);

INVx1_ASAP7_75t_SL g3012 ( 
.A(n_2287),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2035),
.A2(n_1800),
.B1(n_1868),
.B2(n_1863),
.Y(n_3013)
);

INVx2_ASAP7_75t_SL g3014 ( 
.A(n_2287),
.Y(n_3014)
);

OAI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.Y(n_3015)
);

OAI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2505),
.A2(n_1931),
.B(n_1113),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2004),
.B(n_2487),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_SL g3018 ( 
.A(n_2505),
.B(n_834),
.Y(n_3018)
);

OAI21x1_ASAP7_75t_SL g3019 ( 
.A1(n_2012),
.A2(n_2502),
.B(n_2488),
.Y(n_3019)
);

INVx1_ASAP7_75t_SL g3020 ( 
.A(n_2287),
.Y(n_3020)
);

INVxp67_ASAP7_75t_SL g3021 ( 
.A(n_2423),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2004),
.B(n_2487),
.Y(n_3022)
);

INVx4_ASAP7_75t_L g3023 ( 
.A(n_2603),
.Y(n_3023)
);

BUFx8_ASAP7_75t_L g3024 ( 
.A(n_2654),
.Y(n_3024)
);

INVx2_ASAP7_75t_SL g3025 ( 
.A(n_2624),
.Y(n_3025)
);

BUFx3_ASAP7_75t_L g3026 ( 
.A(n_2603),
.Y(n_3026)
);

AOI22xp33_ASAP7_75t_L g3027 ( 
.A1(n_2995),
.A2(n_3018),
.B1(n_2555),
.B2(n_2951),
.Y(n_3027)
);

NAND2x1p5_ASAP7_75t_L g3028 ( 
.A(n_2689),
.B(n_2818),
.Y(n_3028)
);

INVx5_ASAP7_75t_L g3029 ( 
.A(n_2581),
.Y(n_3029)
);

BUFx2_ASAP7_75t_SL g3030 ( 
.A(n_2717),
.Y(n_3030)
);

INVx2_ASAP7_75t_SL g3031 ( 
.A(n_2624),
.Y(n_3031)
);

CKINVDCx5p33_ASAP7_75t_R g3032 ( 
.A(n_2986),
.Y(n_3032)
);

BUFx6f_ASAP7_75t_L g3033 ( 
.A(n_2549),
.Y(n_3033)
);

INVx2_ASAP7_75t_SL g3034 ( 
.A(n_2930),
.Y(n_3034)
);

BUFx4f_ASAP7_75t_L g3035 ( 
.A(n_2899),
.Y(n_3035)
);

AO21x1_ASAP7_75t_L g3036 ( 
.A1(n_2966),
.A2(n_3018),
.B(n_2562),
.Y(n_3036)
);

INVx5_ASAP7_75t_L g3037 ( 
.A(n_2581),
.Y(n_3037)
);

INVx3_ASAP7_75t_L g3038 ( 
.A(n_2732),
.Y(n_3038)
);

INVx3_ASAP7_75t_L g3039 ( 
.A(n_2732),
.Y(n_3039)
);

BUFx2_ASAP7_75t_SL g3040 ( 
.A(n_2717),
.Y(n_3040)
);

BUFx2_ASAP7_75t_L g3041 ( 
.A(n_2742),
.Y(n_3041)
);

AOI22xp33_ASAP7_75t_L g3042 ( 
.A1(n_2995),
.A2(n_2555),
.B1(n_2951),
.B2(n_2552),
.Y(n_3042)
);

AND2x4_ASAP7_75t_L g3043 ( 
.A(n_2651),
.B(n_2708),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2545),
.B(n_2567),
.Y(n_3044)
);

INVx1_ASAP7_75t_SL g3045 ( 
.A(n_2930),
.Y(n_3045)
);

BUFx2_ASAP7_75t_SL g3046 ( 
.A(n_2654),
.Y(n_3046)
);

INVx6_ASAP7_75t_L g3047 ( 
.A(n_2689),
.Y(n_3047)
);

INVxp67_ASAP7_75t_SL g3048 ( 
.A(n_2598),
.Y(n_3048)
);

BUFx3_ASAP7_75t_L g3049 ( 
.A(n_2603),
.Y(n_3049)
);

BUFx12f_ASAP7_75t_L g3050 ( 
.A(n_2576),
.Y(n_3050)
);

INVx1_ASAP7_75t_SL g3051 ( 
.A(n_2640),
.Y(n_3051)
);

BUFx4_ASAP7_75t_SL g3052 ( 
.A(n_2583),
.Y(n_3052)
);

INVx2_ASAP7_75t_SL g3053 ( 
.A(n_2697),
.Y(n_3053)
);

BUFx3_ASAP7_75t_L g3054 ( 
.A(n_2742),
.Y(n_3054)
);

INVx4_ASAP7_75t_L g3055 ( 
.A(n_2689),
.Y(n_3055)
);

BUFx4_ASAP7_75t_SL g3056 ( 
.A(n_2569),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2782),
.Y(n_3057)
);

BUFx2_ASAP7_75t_L g3058 ( 
.A(n_2739),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2630),
.Y(n_3059)
);

NAND2x1p5_ASAP7_75t_L g3060 ( 
.A(n_2689),
.B(n_2818),
.Y(n_3060)
);

INVx3_ASAP7_75t_L g3061 ( 
.A(n_2618),
.Y(n_3061)
);

INVx5_ASAP7_75t_L g3062 ( 
.A(n_2581),
.Y(n_3062)
);

INVx3_ASAP7_75t_SL g3063 ( 
.A(n_2646),
.Y(n_3063)
);

BUFx4f_ASAP7_75t_L g3064 ( 
.A(n_2899),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2630),
.Y(n_3065)
);

BUFx2_ASAP7_75t_L g3066 ( 
.A(n_2739),
.Y(n_3066)
);

INVx3_ASAP7_75t_L g3067 ( 
.A(n_2618),
.Y(n_3067)
);

CKINVDCx20_ASAP7_75t_R g3068 ( 
.A(n_2570),
.Y(n_3068)
);

BUFx3_ASAP7_75t_L g3069 ( 
.A(n_2871),
.Y(n_3069)
);

CKINVDCx5p33_ASAP7_75t_R g3070 ( 
.A(n_2807),
.Y(n_3070)
);

BUFx3_ASAP7_75t_L g3071 ( 
.A(n_2871),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2631),
.Y(n_3072)
);

BUFx3_ASAP7_75t_L g3073 ( 
.A(n_2773),
.Y(n_3073)
);

BUFx2_ASAP7_75t_L g3074 ( 
.A(n_2787),
.Y(n_3074)
);

INVx3_ASAP7_75t_SL g3075 ( 
.A(n_2646),
.Y(n_3075)
);

INVx2_ASAP7_75t_L g3076 ( 
.A(n_2782),
.Y(n_3076)
);

INVx5_ASAP7_75t_L g3077 ( 
.A(n_2581),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2631),
.Y(n_3078)
);

INVx3_ASAP7_75t_L g3079 ( 
.A(n_2618),
.Y(n_3079)
);

BUFx8_ASAP7_75t_L g3080 ( 
.A(n_2654),
.Y(n_3080)
);

BUFx12f_ASAP7_75t_L g3081 ( 
.A(n_2576),
.Y(n_3081)
);

OAI22xp5_ASAP7_75t_L g3082 ( 
.A1(n_2969),
.A2(n_2563),
.B1(n_2966),
.B2(n_2922),
.Y(n_3082)
);

CKINVDCx20_ASAP7_75t_R g3083 ( 
.A(n_2570),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2545),
.B(n_2567),
.Y(n_3084)
);

INVx1_ASAP7_75t_SL g3085 ( 
.A(n_2640),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_2879),
.B(n_2880),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2684),
.B(n_2879),
.Y(n_3087)
);

BUFx8_ASAP7_75t_L g3088 ( 
.A(n_2777),
.Y(n_3088)
);

CKINVDCx6p67_ASAP7_75t_R g3089 ( 
.A(n_2784),
.Y(n_3089)
);

BUFx8_ASAP7_75t_L g3090 ( 
.A(n_2777),
.Y(n_3090)
);

BUFx4_ASAP7_75t_SL g3091 ( 
.A(n_2807),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2632),
.Y(n_3092)
);

INVxp67_ASAP7_75t_SL g3093 ( 
.A(n_2598),
.Y(n_3093)
);

INVx1_ASAP7_75t_SL g3094 ( 
.A(n_3012),
.Y(n_3094)
);

BUFx2_ASAP7_75t_SL g3095 ( 
.A(n_2837),
.Y(n_3095)
);

NAND2x1p5_ASAP7_75t_L g3096 ( 
.A(n_2689),
.B(n_2826),
.Y(n_3096)
);

CKINVDCx6p67_ASAP7_75t_R g3097 ( 
.A(n_2784),
.Y(n_3097)
);

BUFx12f_ASAP7_75t_L g3098 ( 
.A(n_2576),
.Y(n_3098)
);

INVx2_ASAP7_75t_SL g3099 ( 
.A(n_2697),
.Y(n_3099)
);

HB1xp67_ASAP7_75t_L g3100 ( 
.A(n_2904),
.Y(n_3100)
);

BUFx2_ASAP7_75t_R g3101 ( 
.A(n_2882),
.Y(n_3101)
);

BUFx4_ASAP7_75t_SL g3102 ( 
.A(n_2578),
.Y(n_3102)
);

HB1xp67_ASAP7_75t_L g3103 ( 
.A(n_3012),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2632),
.Y(n_3104)
);

INVxp67_ASAP7_75t_SL g3105 ( 
.A(n_2785),
.Y(n_3105)
);

INVx5_ASAP7_75t_SL g3106 ( 
.A(n_2651),
.Y(n_3106)
);

BUFx3_ASAP7_75t_L g3107 ( 
.A(n_2773),
.Y(n_3107)
);

BUFx3_ASAP7_75t_L g3108 ( 
.A(n_2639),
.Y(n_3108)
);

BUFx3_ASAP7_75t_L g3109 ( 
.A(n_2639),
.Y(n_3109)
);

INVx4_ASAP7_75t_L g3110 ( 
.A(n_2689),
.Y(n_3110)
);

BUFx2_ASAP7_75t_L g3111 ( 
.A(n_2787),
.Y(n_3111)
);

BUFx4_ASAP7_75t_SL g3112 ( 
.A(n_2578),
.Y(n_3112)
);

BUFx2_ASAP7_75t_SL g3113 ( 
.A(n_2837),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2668),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2880),
.B(n_2896),
.Y(n_3115)
);

NAND2x1p5_ASAP7_75t_L g3116 ( 
.A(n_2826),
.B(n_2836),
.Y(n_3116)
);

BUFx6f_ASAP7_75t_SL g3117 ( 
.A(n_2817),
.Y(n_3117)
);

BUFx6f_ASAP7_75t_SL g3118 ( 
.A(n_2817),
.Y(n_3118)
);

INVx2_ASAP7_75t_SL g3119 ( 
.A(n_2762),
.Y(n_3119)
);

INVx1_ASAP7_75t_SL g3120 ( 
.A(n_3020),
.Y(n_3120)
);

NAND2x1p5_ASAP7_75t_L g3121 ( 
.A(n_2836),
.B(n_2998),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2896),
.B(n_2949),
.Y(n_3122)
);

CKINVDCx20_ASAP7_75t_R g3123 ( 
.A(n_2947),
.Y(n_3123)
);

AOI22xp5_ASAP7_75t_L g3124 ( 
.A1(n_2552),
.A2(n_2877),
.B1(n_2941),
.B2(n_2873),
.Y(n_3124)
);

BUFx2_ASAP7_75t_L g3125 ( 
.A(n_2776),
.Y(n_3125)
);

BUFx3_ASAP7_75t_L g3126 ( 
.A(n_2639),
.Y(n_3126)
);

AND2x2_ASAP7_75t_L g3127 ( 
.A(n_2949),
.B(n_2964),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2668),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2782),
.Y(n_3129)
);

INVx3_ASAP7_75t_L g3130 ( 
.A(n_2636),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2696),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2828),
.Y(n_3132)
);

INVx3_ASAP7_75t_L g3133 ( 
.A(n_2636),
.Y(n_3133)
);

CKINVDCx20_ASAP7_75t_R g3134 ( 
.A(n_2947),
.Y(n_3134)
);

INVx3_ASAP7_75t_L g3135 ( 
.A(n_2636),
.Y(n_3135)
);

BUFx4f_ASAP7_75t_SL g3136 ( 
.A(n_2810),
.Y(n_3136)
);

INVx3_ASAP7_75t_L g3137 ( 
.A(n_2921),
.Y(n_3137)
);

INVx3_ASAP7_75t_L g3138 ( 
.A(n_2921),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_2943),
.B(n_2960),
.Y(n_3139)
);

INVx2_ASAP7_75t_SL g3140 ( 
.A(n_2762),
.Y(n_3140)
);

CKINVDCx8_ASAP7_75t_R g3141 ( 
.A(n_2557),
.Y(n_3141)
);

INVx3_ASAP7_75t_SL g3142 ( 
.A(n_2646),
.Y(n_3142)
);

INVx1_ASAP7_75t_SL g3143 ( 
.A(n_3020),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2828),
.Y(n_3144)
);

AND2x4_ASAP7_75t_L g3145 ( 
.A(n_2651),
.B(n_2708),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2964),
.B(n_2974),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_2921),
.Y(n_3147)
);

INVx3_ASAP7_75t_L g3148 ( 
.A(n_2925),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_2974),
.B(n_2979),
.Y(n_3149)
);

BUFx2_ASAP7_75t_L g3150 ( 
.A(n_2776),
.Y(n_3150)
);

BUFx12f_ASAP7_75t_L g3151 ( 
.A(n_2576),
.Y(n_3151)
);

BUFx3_ASAP7_75t_L g3152 ( 
.A(n_2604),
.Y(n_3152)
);

INVx8_ASAP7_75t_L g3153 ( 
.A(n_2777),
.Y(n_3153)
);

BUFx12f_ASAP7_75t_L g3154 ( 
.A(n_2811),
.Y(n_3154)
);

INVx8_ASAP7_75t_L g3155 ( 
.A(n_2738),
.Y(n_3155)
);

BUFx4f_ASAP7_75t_SL g3156 ( 
.A(n_2810),
.Y(n_3156)
);

BUFx16f_ASAP7_75t_R g3157 ( 
.A(n_2547),
.Y(n_3157)
);

BUFx3_ASAP7_75t_L g3158 ( 
.A(n_2604),
.Y(n_3158)
);

AOI22xp33_ASAP7_75t_L g3159 ( 
.A1(n_3001),
.A2(n_3013),
.B1(n_2590),
.B2(n_2591),
.Y(n_3159)
);

BUFx2_ASAP7_75t_L g3160 ( 
.A(n_2592),
.Y(n_3160)
);

BUFx4f_ASAP7_75t_L g3161 ( 
.A(n_2899),
.Y(n_3161)
);

BUFx2_ASAP7_75t_R g3162 ( 
.A(n_2946),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2696),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2715),
.Y(n_3164)
);

OR2x6_ASAP7_75t_L g3165 ( 
.A(n_2581),
.B(n_2672),
.Y(n_3165)
);

BUFx2_ASAP7_75t_L g3166 ( 
.A(n_2592),
.Y(n_3166)
);

INVx3_ASAP7_75t_L g3167 ( 
.A(n_2925),
.Y(n_3167)
);

BUFx2_ASAP7_75t_SL g3168 ( 
.A(n_2650),
.Y(n_3168)
);

BUFx2_ASAP7_75t_L g3169 ( 
.A(n_2601),
.Y(n_3169)
);

AND2x2_ASAP7_75t_L g3170 ( 
.A(n_2979),
.B(n_3008),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2715),
.Y(n_3171)
);

BUFx3_ASAP7_75t_L g3172 ( 
.A(n_2794),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2736),
.Y(n_3173)
);

BUFx3_ASAP7_75t_L g3174 ( 
.A(n_2794),
.Y(n_3174)
);

CKINVDCx5p33_ASAP7_75t_R g3175 ( 
.A(n_2811),
.Y(n_3175)
);

BUFx3_ASAP7_75t_L g3176 ( 
.A(n_2774),
.Y(n_3176)
);

NOR2x1_ASAP7_75t_L g3177 ( 
.A(n_2628),
.B(n_2550),
.Y(n_3177)
);

AND2x4_ASAP7_75t_L g3178 ( 
.A(n_2651),
.B(n_2708),
.Y(n_3178)
);

CKINVDCx20_ASAP7_75t_R g3179 ( 
.A(n_2612),
.Y(n_3179)
);

AND2x4_ASAP7_75t_L g3180 ( 
.A(n_2708),
.B(n_2738),
.Y(n_3180)
);

INVx3_ASAP7_75t_SL g3181 ( 
.A(n_2698),
.Y(n_3181)
);

INVx1_ASAP7_75t_SL g3182 ( 
.A(n_2723),
.Y(n_3182)
);

INVx2_ASAP7_75t_SL g3183 ( 
.A(n_2601),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2736),
.Y(n_3184)
);

BUFx3_ASAP7_75t_L g3185 ( 
.A(n_2774),
.Y(n_3185)
);

BUFx3_ASAP7_75t_L g3186 ( 
.A(n_2704),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2737),
.Y(n_3187)
);

AND2x2_ASAP7_75t_L g3188 ( 
.A(n_3008),
.B(n_2608),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2608),
.B(n_2617),
.Y(n_3189)
);

INVx5_ASAP7_75t_L g3190 ( 
.A(n_2672),
.Y(n_3190)
);

INVx6_ASAP7_75t_L g3191 ( 
.A(n_2738),
.Y(n_3191)
);

BUFx2_ASAP7_75t_L g3192 ( 
.A(n_2885),
.Y(n_3192)
);

INVx1_ASAP7_75t_SL g3193 ( 
.A(n_2723),
.Y(n_3193)
);

NOR2xp33_ASAP7_75t_L g3194 ( 
.A(n_2963),
.B(n_2996),
.Y(n_3194)
);

NAND2x1p5_ASAP7_75t_L g3195 ( 
.A(n_2998),
.B(n_2565),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2737),
.Y(n_3196)
);

BUFx2_ASAP7_75t_R g3197 ( 
.A(n_3003),
.Y(n_3197)
);

BUFx2_ASAP7_75t_SL g3198 ( 
.A(n_2709),
.Y(n_3198)
);

INVxp67_ASAP7_75t_SL g3199 ( 
.A(n_2554),
.Y(n_3199)
);

INVx8_ASAP7_75t_L g3200 ( 
.A(n_2738),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2617),
.B(n_2621),
.Y(n_3201)
);

INVxp67_ASAP7_75t_SL g3202 ( 
.A(n_2709),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2621),
.B(n_2600),
.Y(n_3203)
);

INVx2_ASAP7_75t_SL g3204 ( 
.A(n_2885),
.Y(n_3204)
);

INVx2_ASAP7_75t_SL g3205 ( 
.A(n_2892),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2550),
.B(n_2551),
.Y(n_3206)
);

NOR2xp33_ASAP7_75t_L g3207 ( 
.A(n_2999),
.B(n_2579),
.Y(n_3207)
);

INVx3_ASAP7_75t_L g3208 ( 
.A(n_2925),
.Y(n_3208)
);

BUFx3_ASAP7_75t_L g3209 ( 
.A(n_2704),
.Y(n_3209)
);

BUFx3_ASAP7_75t_L g3210 ( 
.A(n_2870),
.Y(n_3210)
);

AND2x2_ASAP7_75t_L g3211 ( 
.A(n_2813),
.B(n_2686),
.Y(n_3211)
);

NOR2xp33_ASAP7_75t_L g3212 ( 
.A(n_2546),
.B(n_2556),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2828),
.Y(n_3213)
);

INVx3_ASAP7_75t_L g3214 ( 
.A(n_2912),
.Y(n_3214)
);

BUFx6f_ASAP7_75t_SL g3215 ( 
.A(n_2612),
.Y(n_3215)
);

BUFx2_ASAP7_75t_L g3216 ( 
.A(n_2892),
.Y(n_3216)
);

BUFx2_ASAP7_75t_L g3217 ( 
.A(n_2937),
.Y(n_3217)
);

BUFx2_ASAP7_75t_L g3218 ( 
.A(n_2937),
.Y(n_3218)
);

CKINVDCx6p67_ASAP7_75t_R g3219 ( 
.A(n_2683),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2828),
.Y(n_3220)
);

CKINVDCx16_ASAP7_75t_R g3221 ( 
.A(n_2683),
.Y(n_3221)
);

OAI22xp5_ASAP7_75t_L g3222 ( 
.A1(n_2969),
.A2(n_2891),
.B1(n_2981),
.B2(n_2950),
.Y(n_3222)
);

NAND2x1p5_ASAP7_75t_L g3223 ( 
.A(n_2596),
.B(n_2738),
.Y(n_3223)
);

INVx1_ASAP7_75t_SL g3224 ( 
.A(n_2765),
.Y(n_3224)
);

NAND2x1p5_ASAP7_75t_L g3225 ( 
.A(n_2740),
.B(n_2657),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2745),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2745),
.Y(n_3227)
);

INVx1_ASAP7_75t_SL g3228 ( 
.A(n_2765),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2764),
.Y(n_3229)
);

NAND2x1p5_ASAP7_75t_L g3230 ( 
.A(n_2740),
.B(n_2649),
.Y(n_3230)
);

INVx8_ASAP7_75t_L g3231 ( 
.A(n_2672),
.Y(n_3231)
);

BUFx3_ASAP7_75t_L g3232 ( 
.A(n_2870),
.Y(n_3232)
);

BUFx3_ASAP7_75t_L g3233 ( 
.A(n_2659),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2764),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2792),
.Y(n_3235)
);

BUFx4f_ASAP7_75t_SL g3236 ( 
.A(n_2886),
.Y(n_3236)
);

BUFx12f_ASAP7_75t_L g3237 ( 
.A(n_2741),
.Y(n_3237)
);

INVx3_ASAP7_75t_L g3238 ( 
.A(n_2912),
.Y(n_3238)
);

INVx1_ASAP7_75t_SL g3239 ( 
.A(n_2687),
.Y(n_3239)
);

BUFx2_ASAP7_75t_L g3240 ( 
.A(n_3014),
.Y(n_3240)
);

BUFx2_ASAP7_75t_SL g3241 ( 
.A(n_2741),
.Y(n_3241)
);

BUFx12f_ASAP7_75t_L g3242 ( 
.A(n_2741),
.Y(n_3242)
);

BUFx3_ASAP7_75t_L g3243 ( 
.A(n_2659),
.Y(n_3243)
);

CKINVDCx16_ASAP7_75t_R g3244 ( 
.A(n_2886),
.Y(n_3244)
);

INVx4_ASAP7_75t_L g3245 ( 
.A(n_2670),
.Y(n_3245)
);

INVx2_ASAP7_75t_SL g3246 ( 
.A(n_3014),
.Y(n_3246)
);

CKINVDCx8_ASAP7_75t_R g3247 ( 
.A(n_2557),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_2813),
.B(n_2686),
.Y(n_3248)
);

INVx1_ASAP7_75t_SL g3249 ( 
.A(n_2687),
.Y(n_3249)
);

INVx1_ASAP7_75t_SL g3250 ( 
.A(n_2935),
.Y(n_3250)
);

CKINVDCx20_ASAP7_75t_R g3251 ( 
.A(n_2890),
.Y(n_3251)
);

BUFx3_ASAP7_75t_L g3252 ( 
.A(n_2754),
.Y(n_3252)
);

BUFx2_ASAP7_75t_L g3253 ( 
.A(n_2662),
.Y(n_3253)
);

BUFx3_ASAP7_75t_L g3254 ( 
.A(n_2754),
.Y(n_3254)
);

AOI22xp33_ASAP7_75t_L g3255 ( 
.A1(n_2591),
.A2(n_2568),
.B1(n_2562),
.B2(n_2571),
.Y(n_3255)
);

INVx1_ASAP7_75t_SL g3256 ( 
.A(n_2935),
.Y(n_3256)
);

CKINVDCx20_ASAP7_75t_R g3257 ( 
.A(n_2890),
.Y(n_3257)
);

BUFx2_ASAP7_75t_L g3258 ( 
.A(n_2662),
.Y(n_3258)
);

BUFx3_ASAP7_75t_L g3259 ( 
.A(n_2656),
.Y(n_3259)
);

INVx4_ASAP7_75t_L g3260 ( 
.A(n_2670),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2792),
.Y(n_3261)
);

BUFx3_ASAP7_75t_L g3262 ( 
.A(n_2656),
.Y(n_3262)
);

INVx3_ASAP7_75t_L g3263 ( 
.A(n_2938),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2801),
.Y(n_3264)
);

CKINVDCx20_ASAP7_75t_R g3265 ( 
.A(n_2895),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_2799),
.Y(n_3266)
);

BUFx2_ASAP7_75t_L g3267 ( 
.A(n_2662),
.Y(n_3267)
);

AND2x4_ASAP7_75t_L g3268 ( 
.A(n_2825),
.B(n_2838),
.Y(n_3268)
);

INVx5_ASAP7_75t_L g3269 ( 
.A(n_2694),
.Y(n_3269)
);

BUFx10_ASAP7_75t_L g3270 ( 
.A(n_2713),
.Y(n_3270)
);

INVx1_ASAP7_75t_SL g3271 ( 
.A(n_2820),
.Y(n_3271)
);

OR2x6_ASAP7_75t_L g3272 ( 
.A(n_2694),
.B(n_2755),
.Y(n_3272)
);

BUFx3_ASAP7_75t_L g3273 ( 
.A(n_2702),
.Y(n_3273)
);

AOI22xp33_ASAP7_75t_SL g3274 ( 
.A1(n_2903),
.A2(n_2916),
.B1(n_3019),
.B2(n_2910),
.Y(n_3274)
);

INVx5_ASAP7_75t_L g3275 ( 
.A(n_2694),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_2801),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2812),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2799),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2666),
.Y(n_3279)
);

BUFx3_ASAP7_75t_L g3280 ( 
.A(n_2702),
.Y(n_3280)
);

INVx1_ASAP7_75t_SL g3281 ( 
.A(n_2820),
.Y(n_3281)
);

BUFx2_ASAP7_75t_R g3282 ( 
.A(n_2895),
.Y(n_3282)
);

INVx2_ASAP7_75t_SL g3283 ( 
.A(n_2728),
.Y(n_3283)
);

INVx8_ASAP7_75t_L g3284 ( 
.A(n_2694),
.Y(n_3284)
);

BUFx3_ASAP7_75t_L g3285 ( 
.A(n_2629),
.Y(n_3285)
);

AND2x2_ASAP7_75t_SL g3286 ( 
.A(n_2718),
.B(n_2924),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_2551),
.B(n_2752),
.Y(n_3287)
);

BUFx4_ASAP7_75t_SL g3288 ( 
.A(n_2936),
.Y(n_3288)
);

INVx5_ASAP7_75t_L g3289 ( 
.A(n_2694),
.Y(n_3289)
);

OR2x2_ASAP7_75t_L g3290 ( 
.A(n_2808),
.B(n_2855),
.Y(n_3290)
);

CKINVDCx5p33_ASAP7_75t_R g3291 ( 
.A(n_2869),
.Y(n_3291)
);

BUFx3_ASAP7_75t_L g3292 ( 
.A(n_2629),
.Y(n_3292)
);

INVx1_ASAP7_75t_SL g3293 ( 
.A(n_2728),
.Y(n_3293)
);

BUFx3_ASAP7_75t_L g3294 ( 
.A(n_2748),
.Y(n_3294)
);

CKINVDCx8_ASAP7_75t_R g3295 ( 
.A(n_2781),
.Y(n_3295)
);

BUFx2_ASAP7_75t_SL g3296 ( 
.A(n_2909),
.Y(n_3296)
);

BUFx8_ASAP7_75t_SL g3297 ( 
.A(n_2905),
.Y(n_3297)
);

CKINVDCx16_ASAP7_75t_R g3298 ( 
.A(n_2936),
.Y(n_3298)
);

INVx3_ASAP7_75t_SL g3299 ( 
.A(n_2731),
.Y(n_3299)
);

INVx5_ASAP7_75t_L g3300 ( 
.A(n_2755),
.Y(n_3300)
);

INVx8_ASAP7_75t_L g3301 ( 
.A(n_2755),
.Y(n_3301)
);

NAND2x1p5_ASAP7_75t_L g3302 ( 
.A(n_2887),
.B(n_2984),
.Y(n_3302)
);

AOI22xp33_ASAP7_75t_L g3303 ( 
.A1(n_2591),
.A2(n_2568),
.B1(n_2586),
.B2(n_2641),
.Y(n_3303)
);

BUFx3_ASAP7_75t_L g3304 ( 
.A(n_2748),
.Y(n_3304)
);

INVx3_ASAP7_75t_SL g3305 ( 
.A(n_2781),
.Y(n_3305)
);

INVx3_ASAP7_75t_L g3306 ( 
.A(n_2938),
.Y(n_3306)
);

INVx5_ASAP7_75t_L g3307 ( 
.A(n_2755),
.Y(n_3307)
);

INVx5_ASAP7_75t_L g3308 ( 
.A(n_2755),
.Y(n_3308)
);

BUFx2_ASAP7_75t_L g3309 ( 
.A(n_2664),
.Y(n_3309)
);

AND2x4_ASAP7_75t_L g3310 ( 
.A(n_2825),
.B(n_2838),
.Y(n_3310)
);

BUFx4f_ASAP7_75t_L g3311 ( 
.A(n_2944),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_2638),
.B(n_2727),
.Y(n_3312)
);

BUFx3_ASAP7_75t_L g3313 ( 
.A(n_2643),
.Y(n_3313)
);

NAND2x1p5_ASAP7_75t_L g3314 ( 
.A(n_2984),
.B(n_2643),
.Y(n_3314)
);

INVx1_ASAP7_75t_SL g3315 ( 
.A(n_2744),
.Y(n_3315)
);

BUFx3_ASAP7_75t_L g3316 ( 
.A(n_2644),
.Y(n_3316)
);

CKINVDCx11_ASAP7_75t_R g3317 ( 
.A(n_2993),
.Y(n_3317)
);

OR2x2_ASAP7_75t_L g3318 ( 
.A(n_2808),
.B(n_2830),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2823),
.Y(n_3319)
);

INVx5_ASAP7_75t_L g3320 ( 
.A(n_2989),
.Y(n_3320)
);

BUFx3_ASAP7_75t_L g3321 ( 
.A(n_2644),
.Y(n_3321)
);

CKINVDCx5p33_ASAP7_75t_R g3322 ( 
.A(n_2993),
.Y(n_3322)
);

BUFx2_ASAP7_75t_L g3323 ( 
.A(n_2664),
.Y(n_3323)
);

INVx3_ASAP7_75t_L g3324 ( 
.A(n_2582),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_2638),
.B(n_2727),
.Y(n_3325)
);

BUFx3_ASAP7_75t_L g3326 ( 
.A(n_2700),
.Y(n_3326)
);

INVxp67_ASAP7_75t_SL g3327 ( 
.A(n_2673),
.Y(n_3327)
);

INVxp67_ASAP7_75t_SL g3328 ( 
.A(n_2733),
.Y(n_3328)
);

INVx1_ASAP7_75t_SL g3329 ( 
.A(n_2693),
.Y(n_3329)
);

INVx8_ASAP7_75t_L g3330 ( 
.A(n_2989),
.Y(n_3330)
);

AOI22xp33_ASAP7_75t_L g3331 ( 
.A1(n_2641),
.A2(n_2589),
.B1(n_2910),
.B2(n_2903),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2584),
.B(n_2753),
.Y(n_3332)
);

INVx1_ASAP7_75t_SL g3333 ( 
.A(n_2859),
.Y(n_3333)
);

BUFx2_ASAP7_75t_L g3334 ( 
.A(n_2788),
.Y(n_3334)
);

BUFx2_ASAP7_75t_SL g3335 ( 
.A(n_3021),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_2711),
.B(n_2830),
.Y(n_3336)
);

INVx2_ASAP7_75t_SL g3337 ( 
.A(n_2750),
.Y(n_3337)
);

INVx3_ASAP7_75t_L g3338 ( 
.A(n_2582),
.Y(n_3338)
);

BUFx3_ASAP7_75t_L g3339 ( 
.A(n_2700),
.Y(n_3339)
);

BUFx3_ASAP7_75t_L g3340 ( 
.A(n_2606),
.Y(n_3340)
);

NOR2xp33_ASAP7_75t_L g3341 ( 
.A(n_2558),
.B(n_2560),
.Y(n_3341)
);

INVx5_ASAP7_75t_L g3342 ( 
.A(n_2989),
.Y(n_3342)
);

BUFx3_ASAP7_75t_L g3343 ( 
.A(n_2606),
.Y(n_3343)
);

INVx5_ASAP7_75t_L g3344 ( 
.A(n_2989),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_2711),
.B(n_2816),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_2725),
.Y(n_3346)
);

BUFx3_ASAP7_75t_L g3347 ( 
.A(n_2594),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_2823),
.Y(n_3348)
);

NOR2xp33_ASAP7_75t_SL g3349 ( 
.A(n_2889),
.B(n_2561),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_2816),
.B(n_2842),
.Y(n_3350)
);

BUFx3_ASAP7_75t_L g3351 ( 
.A(n_2594),
.Y(n_3351)
);

BUFx2_ASAP7_75t_SL g3352 ( 
.A(n_2714),
.Y(n_3352)
);

INVx2_ASAP7_75t_SL g3353 ( 
.A(n_2757),
.Y(n_3353)
);

BUFx3_ASAP7_75t_L g3354 ( 
.A(n_2645),
.Y(n_3354)
);

AND2x4_ASAP7_75t_L g3355 ( 
.A(n_2825),
.B(n_2838),
.Y(n_3355)
);

BUFx3_ASAP7_75t_L g3356 ( 
.A(n_2645),
.Y(n_3356)
);

INVxp67_ASAP7_75t_SL g3357 ( 
.A(n_2733),
.Y(n_3357)
);

OR2x6_ASAP7_75t_L g3358 ( 
.A(n_2724),
.B(n_2800),
.Y(n_3358)
);

AND2x2_ASAP7_75t_L g3359 ( 
.A(n_2842),
.B(n_2844),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_2853),
.Y(n_3360)
);

AOI22xp5_ASAP7_75t_L g3361 ( 
.A1(n_2610),
.A2(n_2889),
.B1(n_2924),
.B2(n_2605),
.Y(n_3361)
);

BUFx12f_ASAP7_75t_L g3362 ( 
.A(n_2846),
.Y(n_3362)
);

OR2x6_ASAP7_75t_L g3363 ( 
.A(n_2724),
.B(n_2800),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_2584),
.B(n_2548),
.Y(n_3364)
);

AND2x4_ASAP7_75t_L g3365 ( 
.A(n_2814),
.B(n_2588),
.Y(n_3365)
);

HB1xp67_ASAP7_75t_L g3366 ( 
.A(n_2758),
.Y(n_3366)
);

CKINVDCx20_ASAP7_75t_R g3367 ( 
.A(n_2905),
.Y(n_3367)
);

NAND2x1p5_ASAP7_75t_L g3368 ( 
.A(n_2815),
.B(n_2674),
.Y(n_3368)
);

CKINVDCx5p33_ASAP7_75t_R g3369 ( 
.A(n_2821),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_2729),
.Y(n_3370)
);

BUFx3_ASAP7_75t_L g3371 ( 
.A(n_2735),
.Y(n_3371)
);

AND2x4_ASAP7_75t_L g3372 ( 
.A(n_2814),
.B(n_2661),
.Y(n_3372)
);

BUFx12f_ASAP7_75t_L g3373 ( 
.A(n_2846),
.Y(n_3373)
);

INVx5_ASAP7_75t_L g3374 ( 
.A(n_2814),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_2584),
.B(n_2705),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_2844),
.B(n_2854),
.Y(n_3376)
);

INVxp67_ASAP7_75t_SL g3377 ( 
.A(n_2554),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_R g3378 ( 
.A(n_2671),
.B(n_2905),
.Y(n_3378)
);

INVx5_ASAP7_75t_L g3379 ( 
.A(n_2975),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_L g3380 ( 
.A(n_2566),
.B(n_2874),
.Y(n_3380)
);

BUFx2_ASAP7_75t_SL g3381 ( 
.A(n_2730),
.Y(n_3381)
);

INVxp67_ASAP7_75t_SL g3382 ( 
.A(n_2691),
.Y(n_3382)
);

BUFx3_ASAP7_75t_L g3383 ( 
.A(n_2695),
.Y(n_3383)
);

CKINVDCx20_ASAP7_75t_R g3384 ( 
.A(n_2953),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_2768),
.Y(n_3385)
);

HB1xp67_ASAP7_75t_L g3386 ( 
.A(n_2761),
.Y(n_3386)
);

BUFx2_ASAP7_75t_L g3387 ( 
.A(n_2851),
.Y(n_3387)
);

INVx1_ASAP7_75t_SL g3388 ( 
.A(n_2872),
.Y(n_3388)
);

BUFx3_ASAP7_75t_L g3389 ( 
.A(n_2695),
.Y(n_3389)
);

BUFx4_ASAP7_75t_SL g3390 ( 
.A(n_2953),
.Y(n_3390)
);

AND2x4_ASAP7_75t_L g3391 ( 
.A(n_2854),
.B(n_2572),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_2665),
.B(n_2660),
.Y(n_3392)
);

INVx6_ASAP7_75t_L g3393 ( 
.A(n_2824),
.Y(n_3393)
);

INVx6_ASAP7_75t_SL g3394 ( 
.A(n_2642),
.Y(n_3394)
);

INVx5_ASAP7_75t_SL g3395 ( 
.A(n_2848),
.Y(n_3395)
);

BUFx3_ASAP7_75t_L g3396 ( 
.A(n_2866),
.Y(n_3396)
);

BUFx3_ASAP7_75t_L g3397 ( 
.A(n_2635),
.Y(n_3397)
);

BUFx10_ASAP7_75t_L g3398 ( 
.A(n_2658),
.Y(n_3398)
);

CKINVDCx5p33_ASAP7_75t_R g3399 ( 
.A(n_2953),
.Y(n_3399)
);

CKINVDCx20_ASAP7_75t_R g3400 ( 
.A(n_2793),
.Y(n_3400)
);

INVx1_ASAP7_75t_SL g3401 ( 
.A(n_2747),
.Y(n_3401)
);

AOI22xp33_ASAP7_75t_L g3402 ( 
.A1(n_2641),
.A2(n_2589),
.B1(n_3019),
.B2(n_2916),
.Y(n_3402)
);

INVx6_ASAP7_75t_SL g3403 ( 
.A(n_2642),
.Y(n_3403)
);

BUFx3_ASAP7_75t_L g3404 ( 
.A(n_2635),
.Y(n_3404)
);

BUFx8_ASAP7_75t_L g3405 ( 
.A(n_2809),
.Y(n_3405)
);

INVx1_ASAP7_75t_SL g3406 ( 
.A(n_2867),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_2809),
.Y(n_3407)
);

AND2x2_ASAP7_75t_L g3408 ( 
.A(n_2778),
.B(n_2780),
.Y(n_3408)
);

CKINVDCx5p33_ASAP7_75t_R g3409 ( 
.A(n_2888),
.Y(n_3409)
);

BUFx6f_ASAP7_75t_L g3410 ( 
.A(n_2720),
.Y(n_3410)
);

BUFx4f_ASAP7_75t_L g3411 ( 
.A(n_2724),
.Y(n_3411)
);

BUFx3_ASAP7_75t_L g3412 ( 
.A(n_2691),
.Y(n_3412)
);

BUFx2_ASAP7_75t_L g3413 ( 
.A(n_2851),
.Y(n_3413)
);

INVx5_ASAP7_75t_SL g3414 ( 
.A(n_2848),
.Y(n_3414)
);

NAND2x1p5_ASAP7_75t_L g3415 ( 
.A(n_2815),
.B(n_2674),
.Y(n_3415)
);

BUFx3_ASAP7_75t_L g3416 ( 
.A(n_2720),
.Y(n_3416)
);

NOR2xp33_ASAP7_75t_L g3417 ( 
.A(n_2893),
.B(n_2900),
.Y(n_3417)
);

OAI22xp5_ASAP7_75t_L g3418 ( 
.A1(n_2987),
.A2(n_3009),
.B1(n_2542),
.B2(n_2898),
.Y(n_3418)
);

INVx1_ASAP7_75t_SL g3419 ( 
.A(n_2751),
.Y(n_3419)
);

INVx1_ASAP7_75t_SL g3420 ( 
.A(n_2746),
.Y(n_3420)
);

BUFx12f_ASAP7_75t_L g3421 ( 
.A(n_2597),
.Y(n_3421)
);

INVx1_ASAP7_75t_SL g3422 ( 
.A(n_2749),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_2802),
.Y(n_3423)
);

INVx4_ASAP7_75t_L g3424 ( 
.A(n_2597),
.Y(n_3424)
);

INVx4_ASAP7_75t_L g3425 ( 
.A(n_2669),
.Y(n_3425)
);

HB1xp67_ASAP7_75t_L g3426 ( 
.A(n_2791),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_2802),
.Y(n_3427)
);

BUFx4f_ASAP7_75t_L g3428 ( 
.A(n_2800),
.Y(n_3428)
);

INVx3_ASAP7_75t_SL g3429 ( 
.A(n_2718),
.Y(n_3429)
);

CKINVDCx5p33_ASAP7_75t_R g3430 ( 
.A(n_2919),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_2853),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_2577),
.Y(n_3432)
);

INVx6_ASAP7_75t_L g3433 ( 
.A(n_2824),
.Y(n_3433)
);

AND2x4_ASAP7_75t_L g3434 ( 
.A(n_2634),
.B(n_2827),
.Y(n_3434)
);

INVx1_ASAP7_75t_SL g3435 ( 
.A(n_2756),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_2789),
.B(n_2790),
.Y(n_3436)
);

BUFx4_ASAP7_75t_SL g3437 ( 
.A(n_2681),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_2857),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_2857),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_2577),
.Y(n_3440)
);

INVx1_ASAP7_75t_SL g3441 ( 
.A(n_2718),
.Y(n_3441)
);

BUFx6f_ASAP7_75t_SL g3442 ( 
.A(n_2609),
.Y(n_3442)
);

BUFx4f_ASAP7_75t_L g3443 ( 
.A(n_2688),
.Y(n_3443)
);

CKINVDCx5p33_ASAP7_75t_R g3444 ( 
.A(n_2920),
.Y(n_3444)
);

BUFx12f_ASAP7_75t_L g3445 ( 
.A(n_2688),
.Y(n_3445)
);

CKINVDCx11_ASAP7_75t_R g3446 ( 
.A(n_2625),
.Y(n_3446)
);

INVx1_ASAP7_75t_SL g3447 ( 
.A(n_2718),
.Y(n_3447)
);

INVx2_ASAP7_75t_SL g3448 ( 
.A(n_2806),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_2860),
.Y(n_3449)
);

INVxp67_ASAP7_75t_SL g3450 ( 
.A(n_2609),
.Y(n_3450)
);

INVx1_ASAP7_75t_SL g3451 ( 
.A(n_2806),
.Y(n_3451)
);

BUFx6f_ASAP7_75t_L g3452 ( 
.A(n_2580),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_2797),
.B(n_2803),
.Y(n_3453)
);

BUFx6f_ASAP7_75t_L g3454 ( 
.A(n_2580),
.Y(n_3454)
);

AND2x2_ASAP7_75t_L g3455 ( 
.A(n_2804),
.B(n_2611),
.Y(n_3455)
);

INVx3_ASAP7_75t_SL g3456 ( 
.A(n_2627),
.Y(n_3456)
);

BUFx8_ASAP7_75t_L g3457 ( 
.A(n_2681),
.Y(n_3457)
);

INVxp67_ASAP7_75t_SL g3458 ( 
.A(n_2881),
.Y(n_3458)
);

INVx6_ASAP7_75t_L g3459 ( 
.A(n_2868),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_2881),
.Y(n_3460)
);

INVx1_ASAP7_75t_SL g3461 ( 
.A(n_2627),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2894),
.Y(n_3462)
);

BUFx8_ASAP7_75t_L g3463 ( 
.A(n_2927),
.Y(n_3463)
);

CKINVDCx14_ASAP7_75t_R g3464 ( 
.A(n_2679),
.Y(n_3464)
);

BUFx3_ASAP7_75t_L g3465 ( 
.A(n_2770),
.Y(n_3465)
);

INVx3_ASAP7_75t_SL g3466 ( 
.A(n_2627),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_2860),
.Y(n_3467)
);

BUFx2_ASAP7_75t_SL g3468 ( 
.A(n_2726),
.Y(n_3468)
);

INVx3_ASAP7_75t_L g3469 ( 
.A(n_2876),
.Y(n_3469)
);

BUFx10_ASAP7_75t_L g3470 ( 
.A(n_2894),
.Y(n_3470)
);

BUFx3_ASAP7_75t_L g3471 ( 
.A(n_2845),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_2907),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_2861),
.Y(n_3473)
);

INVx5_ASAP7_75t_SL g3474 ( 
.A(n_2848),
.Y(n_3474)
);

INVx3_ASAP7_75t_L g3475 ( 
.A(n_2876),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_2861),
.Y(n_3476)
);

BUFx12f_ASAP7_75t_L g3477 ( 
.A(n_2841),
.Y(n_3477)
);

BUFx3_ASAP7_75t_L g3478 ( 
.A(n_2845),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_2907),
.Y(n_3479)
);

NAND2x1p5_ASAP7_75t_L g3480 ( 
.A(n_2682),
.B(n_2767),
.Y(n_3480)
);

CKINVDCx5p33_ASAP7_75t_R g3481 ( 
.A(n_2923),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_2908),
.Y(n_3482)
);

BUFx3_ASAP7_75t_L g3483 ( 
.A(n_2626),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_2908),
.Y(n_3484)
);

BUFx4f_ASAP7_75t_SL g3485 ( 
.A(n_2918),
.Y(n_3485)
);

BUFx3_ASAP7_75t_L g3486 ( 
.A(n_2626),
.Y(n_3486)
);

OAI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_3418),
.A2(n_2958),
.B(n_2884),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_3036),
.A2(n_2875),
.B1(n_2948),
.B2(n_2898),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3287),
.B(n_2573),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3059),
.Y(n_3490)
);

AOI22xp33_ASAP7_75t_L g3491 ( 
.A1(n_3036),
.A2(n_2875),
.B1(n_2956),
.B2(n_2948),
.Y(n_3491)
);

AO21x2_ASAP7_75t_L g3492 ( 
.A1(n_3364),
.A2(n_2593),
.B(n_2675),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_3202),
.A2(n_2897),
.B(n_2883),
.Y(n_3493)
);

OA21x2_ASAP7_75t_L g3494 ( 
.A1(n_3048),
.A2(n_2831),
.B(n_2685),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3059),
.Y(n_3495)
);

OA21x2_ASAP7_75t_L g3496 ( 
.A1(n_3093),
.A2(n_2831),
.B(n_2712),
.Y(n_3496)
);

INVx2_ASAP7_75t_L g3497 ( 
.A(n_3057),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3065),
.Y(n_3498)
);

OAI21x1_ASAP7_75t_L g3499 ( 
.A1(n_3480),
.A2(n_2988),
.B(n_2959),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3044),
.B(n_2611),
.Y(n_3500)
);

CKINVDCx11_ASAP7_75t_R g3501 ( 
.A(n_3068),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3287),
.B(n_2573),
.Y(n_3502)
);

BUFx6f_ASAP7_75t_L g3503 ( 
.A(n_3033),
.Y(n_3503)
);

OAI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_3418),
.A2(n_2906),
.B(n_2901),
.Y(n_3504)
);

AOI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_3082),
.A2(n_2913),
.B(n_2911),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3065),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3057),
.Y(n_3507)
);

OAI221xp5_ASAP7_75t_L g3508 ( 
.A1(n_3361),
.A2(n_2679),
.B1(n_2633),
.B2(n_2595),
.C(n_2602),
.Y(n_3508)
);

NAND2x1p5_ASAP7_75t_L g3509 ( 
.A(n_3055),
.B(n_2622),
.Y(n_3509)
);

AND2x4_ASAP7_75t_L g3510 ( 
.A(n_3152),
.B(n_2648),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3072),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3072),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3078),
.Y(n_3513)
);

BUFx10_ASAP7_75t_L g3514 ( 
.A(n_3215),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3078),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3092),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3057),
.Y(n_3517)
);

AOI22xp33_ASAP7_75t_L g3518 ( 
.A1(n_3303),
.A2(n_2956),
.B1(n_2980),
.B2(n_2976),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_3207),
.B(n_3139),
.Y(n_3519)
);

OR2x2_ASAP7_75t_L g3520 ( 
.A(n_3239),
.B(n_2678),
.Y(n_3520)
);

CKINVDCx20_ASAP7_75t_R g3521 ( 
.A(n_3123),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3044),
.B(n_2703),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3092),
.Y(n_3523)
);

OR2x6_ASAP7_75t_L g3524 ( 
.A(n_3074),
.B(n_2835),
.Y(n_3524)
);

INVx2_ASAP7_75t_L g3525 ( 
.A(n_3076),
.Y(n_3525)
);

AOI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_3027),
.A2(n_2976),
.B1(n_2997),
.B2(n_2980),
.Y(n_3526)
);

OR2x2_ASAP7_75t_L g3527 ( 
.A(n_3239),
.B(n_2692),
.Y(n_3527)
);

HB1xp67_ASAP7_75t_L g3528 ( 
.A(n_3041),
.Y(n_3528)
);

AOI222xp33_ASAP7_75t_L g3529 ( 
.A1(n_3082),
.A2(n_3222),
.B1(n_3255),
.B2(n_3042),
.C1(n_2574),
.C2(n_2553),
.Y(n_3529)
);

AOI221xp5_ASAP7_75t_L g3530 ( 
.A1(n_3328),
.A2(n_2543),
.B1(n_2595),
.B2(n_2707),
.C(n_3006),
.Y(n_3530)
);

AND2x4_ASAP7_75t_L g3531 ( 
.A(n_3152),
.B(n_2647),
.Y(n_3531)
);

HB1xp67_ASAP7_75t_L g3532 ( 
.A(n_3041),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3104),
.Y(n_3533)
);

NOR2x1_ASAP7_75t_R g3534 ( 
.A(n_3050),
.B(n_2933),
.Y(n_3534)
);

NOR2xp33_ASAP7_75t_L g3535 ( 
.A(n_3194),
.B(n_2934),
.Y(n_3535)
);

O2A1O1Ixp33_ASAP7_75t_L g3536 ( 
.A1(n_3222),
.A2(n_2902),
.B(n_2971),
.C(n_3016),
.Y(n_3536)
);

OAI22xp5_ASAP7_75t_L g3537 ( 
.A1(n_3361),
.A2(n_3124),
.B1(n_2553),
.B2(n_3198),
.Y(n_3537)
);

CKINVDCx20_ASAP7_75t_R g3538 ( 
.A(n_3134),
.Y(n_3538)
);

NAND2x1p5_ASAP7_75t_L g3539 ( 
.A(n_3110),
.B(n_2743),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3104),
.Y(n_3540)
);

CKINVDCx6p67_ASAP7_75t_R g3541 ( 
.A(n_3050),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3114),
.Y(n_3542)
);

AOI21x1_ASAP7_75t_L g3543 ( 
.A1(n_3177),
.A2(n_2955),
.B(n_2954),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3114),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3128),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_SL g3546 ( 
.A(n_3108),
.B(n_2783),
.Y(n_3546)
);

AND2x4_ASAP7_75t_L g3547 ( 
.A(n_3152),
.B(n_3158),
.Y(n_3547)
);

OAI21xp5_ASAP7_75t_L g3548 ( 
.A1(n_3177),
.A2(n_2917),
.B(n_2915),
.Y(n_3548)
);

AND2x6_ASAP7_75t_SL g3549 ( 
.A(n_3157),
.B(n_2939),
.Y(n_3549)
);

INVx4_ASAP7_75t_L g3550 ( 
.A(n_3050),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3128),
.Y(n_3551)
);

BUFx12f_ASAP7_75t_L g3552 ( 
.A(n_3317),
.Y(n_3552)
);

INVxp67_ASAP7_75t_L g3553 ( 
.A(n_3103),
.Y(n_3553)
);

INVx3_ASAP7_75t_SL g3554 ( 
.A(n_3322),
.Y(n_3554)
);

OAI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3357),
.A2(n_2931),
.B(n_2926),
.Y(n_3555)
);

AND2x4_ASAP7_75t_L g3556 ( 
.A(n_3158),
.B(n_2663),
.Y(n_3556)
);

BUFx3_ASAP7_75t_L g3557 ( 
.A(n_3081),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3332),
.B(n_2775),
.Y(n_3558)
);

OAI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_3349),
.A2(n_2965),
.B(n_2932),
.Y(n_3559)
);

A2O1A1Ixp33_ASAP7_75t_L g3560 ( 
.A1(n_3074),
.A2(n_2707),
.B(n_2928),
.C(n_3007),
.Y(n_3560)
);

BUFx2_ASAP7_75t_L g3561 ( 
.A(n_3023),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_3349),
.A2(n_2985),
.B(n_2978),
.Y(n_3562)
);

OR2x6_ASAP7_75t_L g3563 ( 
.A(n_3111),
.B(n_2835),
.Y(n_3563)
);

BUFx2_ASAP7_75t_L g3564 ( 
.A(n_3023),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3131),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3131),
.Y(n_3566)
);

CKINVDCx5p33_ASAP7_75t_R g3567 ( 
.A(n_3052),
.Y(n_3567)
);

O2A1O1Ixp33_ASAP7_75t_SL g3568 ( 
.A1(n_3083),
.A2(n_3015),
.B(n_2952),
.C(n_2929),
.Y(n_3568)
);

OAI22xp5_ASAP7_75t_L g3569 ( 
.A1(n_3124),
.A2(n_2994),
.B1(n_3002),
.B2(n_2992),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3163),
.Y(n_3570)
);

AOI22xp33_ASAP7_75t_SL g3571 ( 
.A1(n_3111),
.A2(n_2613),
.B1(n_2616),
.B2(n_2997),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3163),
.Y(n_3572)
);

BUFx2_ASAP7_75t_L g3573 ( 
.A(n_3023),
.Y(n_3573)
);

INVx2_ASAP7_75t_SL g3574 ( 
.A(n_3054),
.Y(n_3574)
);

AO21x2_ASAP7_75t_L g3575 ( 
.A1(n_3423),
.A2(n_2977),
.B(n_2970),
.Y(n_3575)
);

AOI22xp33_ASAP7_75t_SL g3576 ( 
.A1(n_3198),
.A2(n_3011),
.B1(n_3005),
.B2(n_2763),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3164),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3164),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3171),
.Y(n_3579)
);

OAI22xp5_ASAP7_75t_L g3580 ( 
.A1(n_3159),
.A2(n_3011),
.B1(n_2680),
.B2(n_3000),
.Y(n_3580)
);

OA21x2_ASAP7_75t_L g3581 ( 
.A1(n_3382),
.A2(n_3132),
.B(n_3129),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3171),
.Y(n_3582)
);

BUFx2_ASAP7_75t_L g3583 ( 
.A(n_3023),
.Y(n_3583)
);

OAI21x1_ASAP7_75t_L g3584 ( 
.A1(n_3469),
.A2(n_2585),
.B(n_2559),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3332),
.B(n_2775),
.Y(n_3585)
);

AOI22xp33_ASAP7_75t_L g3586 ( 
.A1(n_3464),
.A2(n_2878),
.B1(n_2667),
.B2(n_2699),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3173),
.Y(n_3587)
);

OAI22xp5_ASAP7_75t_L g3588 ( 
.A1(n_3302),
.A2(n_2676),
.B1(n_2544),
.B2(n_2722),
.Y(n_3588)
);

CKINVDCx12_ASAP7_75t_R g3589 ( 
.A(n_3056),
.Y(n_3589)
);

HB1xp67_ASAP7_75t_L g3590 ( 
.A(n_3045),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3173),
.Y(n_3591)
);

AOI22xp33_ASAP7_75t_L g3592 ( 
.A1(n_3108),
.A2(n_2763),
.B1(n_2652),
.B2(n_2796),
.Y(n_3592)
);

HB1xp67_ASAP7_75t_L g3593 ( 
.A(n_3045),
.Y(n_3593)
);

AND2x4_ASAP7_75t_L g3594 ( 
.A(n_3043),
.B(n_2858),
.Y(n_3594)
);

AOI22xp33_ASAP7_75t_SL g3595 ( 
.A1(n_3108),
.A2(n_2914),
.B1(n_2587),
.B2(n_2564),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3184),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3184),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3187),
.Y(n_3598)
);

AOI22xp33_ASAP7_75t_L g3599 ( 
.A1(n_3109),
.A2(n_2849),
.B1(n_2690),
.B2(n_2864),
.Y(n_3599)
);

INVx1_ASAP7_75t_SL g3600 ( 
.A(n_3451),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3187),
.Y(n_3601)
);

OAI21x1_ASAP7_75t_L g3602 ( 
.A1(n_3475),
.A2(n_2599),
.B(n_2710),
.Y(n_3602)
);

BUFx3_ASAP7_75t_L g3603 ( 
.A(n_3081),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_3206),
.A2(n_2991),
.B(n_2721),
.Y(n_3604)
);

BUFx3_ASAP7_75t_L g3605 ( 
.A(n_3081),
.Y(n_3605)
);

AND2x4_ASAP7_75t_L g3606 ( 
.A(n_3043),
.B(n_2834),
.Y(n_3606)
);

OAI21x1_ASAP7_75t_SL g3607 ( 
.A1(n_3206),
.A2(n_2840),
.B(n_2795),
.Y(n_3607)
);

OA21x2_ASAP7_75t_L g3608 ( 
.A1(n_3144),
.A2(n_2587),
.B(n_2863),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_3213),
.Y(n_3609)
);

OAI21x1_ASAP7_75t_L g3610 ( 
.A1(n_3475),
.A2(n_2701),
.B(n_2843),
.Y(n_3610)
);

AOI22xp33_ASAP7_75t_SL g3611 ( 
.A1(n_3109),
.A2(n_2564),
.B1(n_2627),
.B2(n_2962),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_3286),
.A2(n_2833),
.B(n_2856),
.Y(n_3612)
);

OAI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3302),
.A2(n_2982),
.B(n_2957),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_SL g3614 ( 
.A1(n_3302),
.A2(n_2833),
.B(n_2862),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3375),
.B(n_2564),
.Y(n_3615)
);

BUFx2_ASAP7_75t_L g3616 ( 
.A(n_3405),
.Y(n_3616)
);

CKINVDCx9p33_ASAP7_75t_R g3617 ( 
.A(n_3390),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3084),
.B(n_2940),
.Y(n_3618)
);

AND2x4_ASAP7_75t_L g3619 ( 
.A(n_3043),
.B(n_2564),
.Y(n_3619)
);

AOI22xp33_ASAP7_75t_L g3620 ( 
.A1(n_3109),
.A2(n_2849),
.B1(n_2865),
.B2(n_2771),
.Y(n_3620)
);

OAI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_3435),
.A2(n_3022),
.B1(n_3017),
.B2(n_2967),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3196),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3196),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_3220),
.Y(n_3624)
);

INVx6_ASAP7_75t_L g3625 ( 
.A(n_3457),
.Y(n_3625)
);

NOR2xp33_ASAP7_75t_L g3626 ( 
.A(n_3221),
.B(n_2942),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3220),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3226),
.Y(n_3628)
);

AND2x2_ASAP7_75t_L g3629 ( 
.A(n_3084),
.B(n_2940),
.Y(n_3629)
);

CKINVDCx8_ASAP7_75t_R g3630 ( 
.A(n_3030),
.Y(n_3630)
);

BUFx3_ASAP7_75t_L g3631 ( 
.A(n_3098),
.Y(n_3631)
);

INVx8_ASAP7_75t_L g3632 ( 
.A(n_3098),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3226),
.Y(n_3633)
);

INVx3_ASAP7_75t_L g3634 ( 
.A(n_3371),
.Y(n_3634)
);

NOR2xp33_ASAP7_75t_L g3635 ( 
.A(n_3221),
.B(n_3010),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3227),
.Y(n_3636)
);

AND2x4_ASAP7_75t_L g3637 ( 
.A(n_3043),
.B(n_2564),
.Y(n_3637)
);

NOR2x1_ASAP7_75t_SL g3638 ( 
.A(n_3026),
.B(n_2760),
.Y(n_3638)
);

BUFx2_ASAP7_75t_SL g3639 ( 
.A(n_3141),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3375),
.B(n_2822),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3227),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3229),
.Y(n_3642)
);

OAI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3435),
.A2(n_2972),
.B(n_2945),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3229),
.Y(n_3644)
);

AND2x2_ASAP7_75t_L g3645 ( 
.A(n_3086),
.B(n_2962),
.Y(n_3645)
);

AND2x4_ASAP7_75t_L g3646 ( 
.A(n_3145),
.B(n_2779),
.Y(n_3646)
);

AOI22xp5_ASAP7_75t_L g3647 ( 
.A1(n_3400),
.A2(n_3004),
.B1(n_2968),
.B2(n_2973),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3234),
.Y(n_3648)
);

OR2x2_ASAP7_75t_L g3649 ( 
.A(n_3249),
.B(n_2772),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3234),
.Y(n_3650)
);

CKINVDCx11_ASAP7_75t_R g3651 ( 
.A(n_3179),
.Y(n_3651)
);

BUFx3_ASAP7_75t_L g3652 ( 
.A(n_3098),
.Y(n_3652)
);

BUFx12f_ASAP7_75t_L g3653 ( 
.A(n_3151),
.Y(n_3653)
);

AND2x2_ASAP7_75t_L g3654 ( 
.A(n_3086),
.B(n_2962),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3235),
.Y(n_3655)
);

OR2x6_ASAP7_75t_L g3656 ( 
.A(n_3165),
.B(n_2819),
.Y(n_3656)
);

OAI22xp5_ASAP7_75t_L g3657 ( 
.A1(n_3331),
.A2(n_2990),
.B1(n_2961),
.B2(n_2983),
.Y(n_3657)
);

AND2x2_ASAP7_75t_L g3658 ( 
.A(n_3127),
.B(n_2962),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3235),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3401),
.B(n_3420),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3127),
.B(n_2962),
.Y(n_3661)
);

A2O1A1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_3126),
.A2(n_2653),
.B(n_2607),
.C(n_2614),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3261),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3261),
.Y(n_3664)
);

BUFx3_ASAP7_75t_L g3665 ( 
.A(n_3151),
.Y(n_3665)
);

AOI22xp33_ASAP7_75t_L g3666 ( 
.A1(n_3126),
.A2(n_2849),
.B1(n_2766),
.B2(n_2734),
.Y(n_3666)
);

O2A1O1Ixp33_ASAP7_75t_SL g3667 ( 
.A1(n_3367),
.A2(n_2677),
.B(n_2615),
.C(n_2619),
.Y(n_3667)
);

INVx4_ASAP7_75t_SL g3668 ( 
.A(n_3191),
.Y(n_3668)
);

NAND2x1p5_ASAP7_75t_L g3669 ( 
.A(n_3035),
.B(n_2849),
.Y(n_3669)
);

OAI22x1_ASAP7_75t_L g3670 ( 
.A1(n_3429),
.A2(n_2623),
.B1(n_2575),
.B2(n_2655),
.Y(n_3670)
);

AOI22xp33_ASAP7_75t_L g3671 ( 
.A1(n_3126),
.A2(n_3419),
.B1(n_3299),
.B2(n_3286),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3401),
.B(n_2940),
.Y(n_3672)
);

OAI22xp33_ASAP7_75t_L g3673 ( 
.A1(n_3299),
.A2(n_2786),
.B1(n_2798),
.B2(n_2805),
.Y(n_3673)
);

NOR2xp33_ASAP7_75t_L g3674 ( 
.A(n_3244),
.B(n_2832),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3264),
.Y(n_3675)
);

OAI21x1_ASAP7_75t_L g3676 ( 
.A1(n_3324),
.A2(n_3338),
.B(n_3314),
.Y(n_3676)
);

OAI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_3274),
.A2(n_2940),
.B(n_2716),
.Y(n_3677)
);

BUFx3_ASAP7_75t_L g3678 ( 
.A(n_3151),
.Y(n_3678)
);

AOI21xp5_ASAP7_75t_L g3679 ( 
.A1(n_3286),
.A2(n_2719),
.B(n_2940),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3420),
.B(n_2637),
.Y(n_3680)
);

AOI22xp33_ASAP7_75t_L g3681 ( 
.A1(n_3419),
.A2(n_2868),
.B1(n_2829),
.B2(n_2839),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3264),
.Y(n_3682)
);

AND2x4_ASAP7_75t_L g3683 ( 
.A(n_3145),
.B(n_2620),
.Y(n_3683)
);

AOI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_3035),
.A2(n_2850),
.B(n_2706),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3244),
.B(n_2847),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3276),
.Y(n_3686)
);

BUFx4f_ASAP7_75t_L g3687 ( 
.A(n_3028),
.Y(n_3687)
);

INVx2_ASAP7_75t_SL g3688 ( 
.A(n_3054),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3276),
.Y(n_3689)
);

AOI22xp33_ASAP7_75t_L g3690 ( 
.A1(n_3299),
.A2(n_2852),
.B1(n_2706),
.B2(n_2637),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3277),
.Y(n_3691)
);

AND2x4_ASAP7_75t_L g3692 ( 
.A(n_3145),
.B(n_2620),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3277),
.Y(n_3693)
);

OAI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3274),
.A2(n_2637),
.B(n_2620),
.Y(n_3694)
);

NAND2xp33_ASAP7_75t_R g3695 ( 
.A(n_3032),
.B(n_2637),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_3422),
.B(n_2620),
.Y(n_3696)
);

OAI21x1_ASAP7_75t_L g3697 ( 
.A1(n_3314),
.A2(n_2706),
.B(n_2759),
.Y(n_3697)
);

NOR2xp33_ASAP7_75t_L g3698 ( 
.A(n_3298),
.B(n_2769),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3279),
.Y(n_3699)
);

AOI21xp5_ASAP7_75t_L g3700 ( 
.A1(n_3035),
.A2(n_2759),
.B(n_2769),
.Y(n_3700)
);

OAI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3402),
.A2(n_3426),
.B(n_3157),
.Y(n_3701)
);

AOI22xp33_ASAP7_75t_L g3702 ( 
.A1(n_3455),
.A2(n_2759),
.B1(n_2769),
.B2(n_3446),
.Y(n_3702)
);

OAI21x1_ASAP7_75t_L g3703 ( 
.A1(n_3038),
.A2(n_3039),
.B(n_3368),
.Y(n_3703)
);

OAI21x1_ASAP7_75t_L g3704 ( 
.A1(n_3038),
.A2(n_3039),
.B(n_3368),
.Y(n_3704)
);

OAI21x1_ASAP7_75t_L g3705 ( 
.A1(n_3038),
.A2(n_3039),
.B(n_3368),
.Y(n_3705)
);

OAI21x1_ASAP7_75t_L g3706 ( 
.A1(n_3038),
.A2(n_3039),
.B(n_3415),
.Y(n_3706)
);

AND2x4_ASAP7_75t_L g3707 ( 
.A(n_3178),
.B(n_3180),
.Y(n_3707)
);

OAI21x1_ASAP7_75t_L g3708 ( 
.A1(n_3415),
.A2(n_3223),
.B(n_3214),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3279),
.Y(n_3709)
);

CKINVDCx5p33_ASAP7_75t_R g3710 ( 
.A(n_3091),
.Y(n_3710)
);

CKINVDCx11_ASAP7_75t_R g3711 ( 
.A(n_3251),
.Y(n_3711)
);

OAI21x1_ASAP7_75t_L g3712 ( 
.A1(n_3415),
.A2(n_3223),
.B(n_3214),
.Y(n_3712)
);

OAI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_3334),
.A2(n_3066),
.B(n_3058),
.Y(n_3713)
);

OAI21x1_ASAP7_75t_L g3714 ( 
.A1(n_3223),
.A2(n_3238),
.B(n_3214),
.Y(n_3714)
);

OAI21x1_ASAP7_75t_L g3715 ( 
.A1(n_3214),
.A2(n_3263),
.B(n_3238),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3422),
.B(n_3203),
.Y(n_3716)
);

AO31x2_ASAP7_75t_L g3717 ( 
.A1(n_3427),
.A2(n_3440),
.A3(n_3460),
.B(n_3432),
.Y(n_3717)
);

AOI22xp33_ASAP7_75t_SL g3718 ( 
.A1(n_3026),
.A2(n_3049),
.B1(n_3381),
.B2(n_3352),
.Y(n_3718)
);

A2O1A1Ixp33_ASAP7_75t_L g3719 ( 
.A1(n_3026),
.A2(n_3049),
.B(n_3381),
.C(n_3209),
.Y(n_3719)
);

OAI21x1_ASAP7_75t_L g3720 ( 
.A1(n_3238),
.A2(n_3306),
.B(n_3263),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3058),
.B(n_3066),
.Y(n_3721)
);

OAI221xp5_ASAP7_75t_L g3722 ( 
.A1(n_3429),
.A2(n_3168),
.B1(n_3352),
.B2(n_3334),
.C(n_3456),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3149),
.B(n_3170),
.Y(n_3723)
);

INVx2_ASAP7_75t_SL g3724 ( 
.A(n_3054),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3224),
.B(n_3228),
.Y(n_3725)
);

OAI21x1_ASAP7_75t_L g3726 ( 
.A1(n_3238),
.A2(n_3306),
.B(n_3263),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3224),
.B(n_3228),
.Y(n_3727)
);

AOI22xp33_ASAP7_75t_L g3728 ( 
.A1(n_3455),
.A2(n_3429),
.B1(n_3049),
.B2(n_3209),
.Y(n_3728)
);

HB1xp67_ASAP7_75t_L g3729 ( 
.A(n_3100),
.Y(n_3729)
);

OA21x2_ASAP7_75t_L g3730 ( 
.A1(n_3105),
.A2(n_3431),
.B(n_3360),
.Y(n_3730)
);

AND2x4_ASAP7_75t_L g3731 ( 
.A(n_3178),
.B(n_3180),
.Y(n_3731)
);

NOR2xp67_ASAP7_75t_SL g3732 ( 
.A(n_3141),
.B(n_3247),
.Y(n_3732)
);

A2O1A1Ixp33_ASAP7_75t_L g3733 ( 
.A1(n_3186),
.A2(n_3209),
.B(n_3447),
.C(n_3441),
.Y(n_3733)
);

OAI21x1_ASAP7_75t_L g3734 ( 
.A1(n_3263),
.A2(n_3306),
.B(n_3195),
.Y(n_3734)
);

OAI21x1_ASAP7_75t_L g3735 ( 
.A1(n_3306),
.A2(n_3195),
.B(n_3230),
.Y(n_3735)
);

BUFx2_ASAP7_75t_R g3736 ( 
.A(n_3297),
.Y(n_3736)
);

OAI211xp5_ASAP7_75t_SL g3737 ( 
.A1(n_3327),
.A2(n_3293),
.B(n_3315),
.C(n_3283),
.Y(n_3737)
);

AO21x2_ASAP7_75t_L g3738 ( 
.A1(n_3360),
.A2(n_3438),
.B(n_3431),
.Y(n_3738)
);

CKINVDCx11_ASAP7_75t_R g3739 ( 
.A(n_3257),
.Y(n_3739)
);

OAI21x1_ASAP7_75t_L g3740 ( 
.A1(n_3195),
.A2(n_3230),
.B(n_3225),
.Y(n_3740)
);

INVx4_ASAP7_75t_L g3741 ( 
.A(n_3237),
.Y(n_3741)
);

INVx2_ASAP7_75t_SL g3742 ( 
.A(n_3025),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3087),
.B(n_3250),
.Y(n_3743)
);

INVx1_ASAP7_75t_SL g3744 ( 
.A(n_3451),
.Y(n_3744)
);

OAI21x1_ASAP7_75t_L g3745 ( 
.A1(n_3230),
.A2(n_3225),
.B(n_3360),
.Y(n_3745)
);

NOR2xp33_ASAP7_75t_L g3746 ( 
.A(n_3298),
.B(n_3154),
.Y(n_3746)
);

AOI22xp33_ASAP7_75t_L g3747 ( 
.A1(n_3186),
.A2(n_3107),
.B1(n_3073),
.B2(n_3463),
.Y(n_3747)
);

CKINVDCx5p33_ASAP7_75t_R g3748 ( 
.A(n_3102),
.Y(n_3748)
);

CKINVDCx20_ASAP7_75t_R g3749 ( 
.A(n_3265),
.Y(n_3749)
);

OAI21x1_ASAP7_75t_L g3750 ( 
.A1(n_3438),
.A2(n_3449),
.B(n_3439),
.Y(n_3750)
);

OR2x2_ASAP7_75t_L g3751 ( 
.A(n_3256),
.B(n_3318),
.Y(n_3751)
);

AO31x2_ASAP7_75t_L g3752 ( 
.A1(n_3432),
.A2(n_3440),
.A3(n_3462),
.B(n_3460),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3149),
.B(n_3170),
.Y(n_3753)
);

CKINVDCx5p33_ASAP7_75t_R g3754 ( 
.A(n_3112),
.Y(n_3754)
);

OAI21x1_ASAP7_75t_L g3755 ( 
.A1(n_3439),
.A2(n_3467),
.B(n_3449),
.Y(n_3755)
);

OAI21x1_ASAP7_75t_L g3756 ( 
.A1(n_3439),
.A2(n_3467),
.B(n_3449),
.Y(n_3756)
);

OAI21x1_ASAP7_75t_L g3757 ( 
.A1(n_3467),
.A2(n_3476),
.B(n_3473),
.Y(n_3757)
);

OR2x2_ASAP7_75t_L g3758 ( 
.A(n_3256),
.B(n_3318),
.Y(n_3758)
);

BUFx12f_ASAP7_75t_L g3759 ( 
.A(n_3070),
.Y(n_3759)
);

INVx4_ASAP7_75t_L g3760 ( 
.A(n_3237),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3087),
.B(n_3051),
.Y(n_3761)
);

AOI22xp33_ASAP7_75t_SL g3762 ( 
.A1(n_3168),
.A2(n_3441),
.B1(n_3447),
.B2(n_3186),
.Y(n_3762)
);

BUFx8_ASAP7_75t_L g3763 ( 
.A(n_3215),
.Y(n_3763)
);

BUFx3_ASAP7_75t_L g3764 ( 
.A(n_3024),
.Y(n_3764)
);

AO21x2_ASAP7_75t_L g3765 ( 
.A1(n_3473),
.A2(n_3476),
.B(n_3472),
.Y(n_3765)
);

AND2x4_ASAP7_75t_L g3766 ( 
.A(n_3178),
.B(n_3180),
.Y(n_3766)
);

OAI21x1_ASAP7_75t_L g3767 ( 
.A1(n_3028),
.A2(n_3096),
.B(n_3060),
.Y(n_3767)
);

BUFx3_ASAP7_75t_L g3768 ( 
.A(n_3024),
.Y(n_3768)
);

OAI21x1_ASAP7_75t_L g3769 ( 
.A1(n_3028),
.A2(n_3096),
.B(n_3060),
.Y(n_3769)
);

BUFx3_ASAP7_75t_L g3770 ( 
.A(n_3024),
.Y(n_3770)
);

OA21x2_ASAP7_75t_L g3771 ( 
.A1(n_3461),
.A2(n_3377),
.B(n_3199),
.Y(n_3771)
);

HB1xp67_ASAP7_75t_L g3772 ( 
.A(n_3125),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3211),
.B(n_3248),
.Y(n_3773)
);

BUFx3_ASAP7_75t_L g3774 ( 
.A(n_3024),
.Y(n_3774)
);

AOI21xp5_ASAP7_75t_L g3775 ( 
.A1(n_3064),
.A2(n_3311),
.B(n_3161),
.Y(n_3775)
);

OAI21x1_ASAP7_75t_L g3776 ( 
.A1(n_3096),
.A2(n_3116),
.B(n_3121),
.Y(n_3776)
);

CKINVDCx5p33_ASAP7_75t_R g3777 ( 
.A(n_3288),
.Y(n_3777)
);

AO21x2_ASAP7_75t_L g3778 ( 
.A1(n_3462),
.A2(n_3479),
.B(n_3472),
.Y(n_3778)
);

OAI21x1_ASAP7_75t_L g3779 ( 
.A1(n_3116),
.A2(n_3121),
.B(n_3199),
.Y(n_3779)
);

OAI21x1_ASAP7_75t_L g3780 ( 
.A1(n_3116),
.A2(n_3121),
.B(n_3377),
.Y(n_3780)
);

AO31x2_ASAP7_75t_L g3781 ( 
.A1(n_3479),
.A2(n_3484),
.A3(n_3482),
.B(n_3278),
.Y(n_3781)
);

OAI21x1_ASAP7_75t_L g3782 ( 
.A1(n_3482),
.A2(n_3484),
.B(n_3067),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3051),
.B(n_3085),
.Y(n_3783)
);

AOI22xp33_ASAP7_75t_SL g3784 ( 
.A1(n_3347),
.A2(n_3351),
.B1(n_3107),
.B2(n_3073),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3457),
.B(n_3448),
.Y(n_3785)
);

BUFx2_ASAP7_75t_SL g3786 ( 
.A(n_3141),
.Y(n_3786)
);

OAI22xp5_ASAP7_75t_L g3787 ( 
.A1(n_3347),
.A2(n_3351),
.B1(n_3430),
.B2(n_3409),
.Y(n_3787)
);

NOR2xp33_ASAP7_75t_L g3788 ( 
.A(n_3154),
.B(n_3369),
.Y(n_3788)
);

OR2x4_ASAP7_75t_L g3789 ( 
.A(n_3290),
.B(n_3437),
.Y(n_3789)
);

OAI21x1_ASAP7_75t_L g3790 ( 
.A1(n_3061),
.A2(n_3079),
.B(n_3067),
.Y(n_3790)
);

OR2x2_ASAP7_75t_L g3791 ( 
.A(n_3115),
.B(n_3122),
.Y(n_3791)
);

AO21x2_ASAP7_75t_L g3792 ( 
.A1(n_3450),
.A2(n_3458),
.B(n_3278),
.Y(n_3792)
);

OAI21x1_ASAP7_75t_L g3793 ( 
.A1(n_3061),
.A2(n_3079),
.B(n_3067),
.Y(n_3793)
);

OAI21x1_ASAP7_75t_L g3794 ( 
.A1(n_3061),
.A2(n_3079),
.B(n_3067),
.Y(n_3794)
);

AO21x2_ASAP7_75t_L g3795 ( 
.A1(n_3266),
.A2(n_3319),
.B(n_3278),
.Y(n_3795)
);

OAI22xp5_ASAP7_75t_L g3796 ( 
.A1(n_3347),
.A2(n_3351),
.B1(n_3481),
.B2(n_3444),
.Y(n_3796)
);

OAI21x1_ASAP7_75t_L g3797 ( 
.A1(n_3061),
.A2(n_3130),
.B(n_3079),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_SL g3798 ( 
.A(n_3457),
.B(n_3448),
.Y(n_3798)
);

NOR2xp33_ASAP7_75t_L g3799 ( 
.A(n_3154),
.B(n_3236),
.Y(n_3799)
);

OAI21x1_ASAP7_75t_L g3800 ( 
.A1(n_3130),
.A2(n_3135),
.B(n_3133),
.Y(n_3800)
);

OAI21xp5_ASAP7_75t_L g3801 ( 
.A1(n_3387),
.A2(n_3413),
.B(n_3461),
.Y(n_3801)
);

AND2x2_ASAP7_75t_L g3802 ( 
.A(n_3211),
.B(n_3248),
.Y(n_3802)
);

NOR2xp33_ASAP7_75t_L g3803 ( 
.A(n_3282),
.B(n_3291),
.Y(n_3803)
);

HB1xp67_ASAP7_75t_L g3804 ( 
.A(n_3125),
.Y(n_3804)
);

AOI22xp33_ASAP7_75t_L g3805 ( 
.A1(n_3073),
.A2(n_3107),
.B1(n_3463),
.B2(n_3284),
.Y(n_3805)
);

AOI22xp33_ASAP7_75t_SL g3806 ( 
.A1(n_3465),
.A2(n_3185),
.B1(n_3176),
.B2(n_3457),
.Y(n_3806)
);

OAI21x1_ASAP7_75t_L g3807 ( 
.A1(n_3130),
.A2(n_3135),
.B(n_3133),
.Y(n_3807)
);

NOR2x1_ASAP7_75t_SL g3808 ( 
.A(n_3421),
.B(n_3445),
.Y(n_3808)
);

OA21x2_ASAP7_75t_L g3809 ( 
.A1(n_3434),
.A2(n_3413),
.B(n_3387),
.Y(n_3809)
);

NOR2xp33_ASAP7_75t_SL g3810 ( 
.A(n_3101),
.B(n_3162),
.Y(n_3810)
);

AND2x4_ASAP7_75t_L g3811 ( 
.A(n_3178),
.B(n_3180),
.Y(n_3811)
);

OA21x2_ASAP7_75t_L g3812 ( 
.A1(n_3434),
.A2(n_3391),
.B(n_3372),
.Y(n_3812)
);

OAI22xp5_ASAP7_75t_L g3813 ( 
.A1(n_3101),
.A2(n_3197),
.B1(n_3162),
.B2(n_3122),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3085),
.B(n_3094),
.Y(n_3814)
);

INVxp67_ASAP7_75t_L g3815 ( 
.A(n_3283),
.Y(n_3815)
);

OAI21x1_ASAP7_75t_L g3816 ( 
.A1(n_3130),
.A2(n_3135),
.B(n_3133),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3094),
.B(n_3120),
.Y(n_3817)
);

INVxp67_ASAP7_75t_L g3818 ( 
.A(n_3160),
.Y(n_3818)
);

HB1xp67_ASAP7_75t_L g3819 ( 
.A(n_3150),
.Y(n_3819)
);

OAI22xp33_ASAP7_75t_L g3820 ( 
.A1(n_3456),
.A2(n_3466),
.B1(n_3394),
.B2(n_3403),
.Y(n_3820)
);

OA21x2_ASAP7_75t_L g3821 ( 
.A1(n_3434),
.A2(n_3391),
.B(n_3372),
.Y(n_3821)
);

OAI222xp33_ASAP7_75t_L g3822 ( 
.A1(n_3115),
.A2(n_3146),
.B1(n_3201),
.B2(n_3189),
.C1(n_3165),
.C2(n_3272),
.Y(n_3822)
);

OAI21x1_ASAP7_75t_L g3823 ( 
.A1(n_3133),
.A2(n_3137),
.B(n_3135),
.Y(n_3823)
);

OAI21x1_ASAP7_75t_L g3824 ( 
.A1(n_3137),
.A2(n_3147),
.B(n_3138),
.Y(n_3824)
);

AND2x4_ASAP7_75t_L g3825 ( 
.A(n_3233),
.B(n_3243),
.Y(n_3825)
);

AND2x4_ASAP7_75t_L g3826 ( 
.A(n_3233),
.B(n_3243),
.Y(n_3826)
);

AOI221xp5_ASAP7_75t_L g3827 ( 
.A1(n_3329),
.A2(n_3315),
.B1(n_3212),
.B2(n_3380),
.C(n_3341),
.Y(n_3827)
);

OAI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3417),
.A2(n_3143),
.B(n_3120),
.Y(n_3828)
);

OA21x2_ASAP7_75t_L g3829 ( 
.A1(n_3434),
.A2(n_3391),
.B(n_3372),
.Y(n_3829)
);

AOI21x1_ASAP7_75t_L g3830 ( 
.A1(n_3253),
.A2(n_3267),
.B(n_3258),
.Y(n_3830)
);

AO21x2_ASAP7_75t_L g3831 ( 
.A1(n_3319),
.A2(n_3348),
.B(n_3346),
.Y(n_3831)
);

O2A1O1Ixp33_ASAP7_75t_SL g3832 ( 
.A1(n_3384),
.A2(n_3293),
.B(n_3031),
.C(n_3034),
.Y(n_3832)
);

OAI22xp5_ASAP7_75t_L g3833 ( 
.A1(n_3197),
.A2(n_3146),
.B1(n_3201),
.B2(n_3189),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3064),
.A2(n_3311),
.B(n_3161),
.Y(n_3834)
);

AND2x2_ASAP7_75t_L g3835 ( 
.A(n_3188),
.B(n_3336),
.Y(n_3835)
);

AND2x4_ASAP7_75t_L g3836 ( 
.A(n_3233),
.B(n_3243),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3188),
.B(n_3336),
.Y(n_3837)
);

INVx3_ASAP7_75t_L g3838 ( 
.A(n_3483),
.Y(n_3838)
);

O2A1O1Ixp33_ASAP7_75t_L g3839 ( 
.A1(n_3456),
.A2(n_3466),
.B(n_3182),
.C(n_3193),
.Y(n_3839)
);

OA21x2_ASAP7_75t_L g3840 ( 
.A1(n_3391),
.A2(n_3372),
.B(n_3258),
.Y(n_3840)
);

OAI21x1_ASAP7_75t_L g3841 ( 
.A1(n_3137),
.A2(n_3147),
.B(n_3138),
.Y(n_3841)
);

OAI21x1_ASAP7_75t_L g3842 ( 
.A1(n_3137),
.A2(n_3147),
.B(n_3138),
.Y(n_3842)
);

AOI21xp5_ASAP7_75t_L g3843 ( 
.A1(n_3161),
.A2(n_3311),
.B(n_3443),
.Y(n_3843)
);

OAI21xp5_ASAP7_75t_L g3844 ( 
.A1(n_3143),
.A2(n_3193),
.B(n_3182),
.Y(n_3844)
);

OAI22xp33_ASAP7_75t_L g3845 ( 
.A1(n_3466),
.A2(n_3394),
.B1(n_3403),
.B2(n_3393),
.Y(n_3845)
);

OR2x2_ASAP7_75t_L g3846 ( 
.A(n_3290),
.B(n_3337),
.Y(n_3846)
);

OAI221xp5_ASAP7_75t_L g3847 ( 
.A1(n_3465),
.A2(n_3071),
.B1(n_3069),
.B2(n_3329),
.C(n_3185),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3271),
.B(n_3281),
.Y(n_3848)
);

OAI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3271),
.A2(n_3281),
.B(n_3031),
.Y(n_3849)
);

AOI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_3443),
.A2(n_3428),
.B(n_3411),
.Y(n_3850)
);

OAI21x1_ASAP7_75t_L g3851 ( 
.A1(n_3138),
.A2(n_3148),
.B(n_3147),
.Y(n_3851)
);

INVx1_ASAP7_75t_SL g3852 ( 
.A(n_3160),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_3025),
.B(n_3034),
.Y(n_3853)
);

INVx1_ASAP7_75t_SL g3854 ( 
.A(n_3166),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3370),
.Y(n_3855)
);

INVx5_ASAP7_75t_L g3856 ( 
.A(n_3191),
.Y(n_3856)
);

INVx6_ASAP7_75t_L g3857 ( 
.A(n_3088),
.Y(n_3857)
);

OAI222xp33_ASAP7_75t_L g3858 ( 
.A1(n_3165),
.A2(n_3272),
.B1(n_3388),
.B2(n_3406),
.C1(n_3392),
.C2(n_3308),
.Y(n_3858)
);

OAI21x1_ASAP7_75t_L g3859 ( 
.A1(n_3167),
.A2(n_3208),
.B(n_3385),
.Y(n_3859)
);

OAI21x1_ASAP7_75t_L g3860 ( 
.A1(n_3395),
.A2(n_3474),
.B(n_3414),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3366),
.B(n_3386),
.Y(n_3861)
);

AOI21xp5_ASAP7_75t_L g3862 ( 
.A1(n_3443),
.A2(n_3428),
.B(n_3411),
.Y(n_3862)
);

INVxp67_ASAP7_75t_SL g3863 ( 
.A(n_3150),
.Y(n_3863)
);

A2O1A1Ixp33_ASAP7_75t_L g3864 ( 
.A1(n_3465),
.A2(n_3185),
.B(n_3176),
.C(n_3071),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_SL g3865 ( 
.A(n_3247),
.B(n_3270),
.Y(n_3865)
);

OAI21x1_ASAP7_75t_L g3866 ( 
.A1(n_3395),
.A2(n_3474),
.B(n_3414),
.Y(n_3866)
);

HB1xp67_ASAP7_75t_L g3867 ( 
.A(n_3166),
.Y(n_3867)
);

OAI22xp33_ASAP7_75t_L g3868 ( 
.A1(n_3394),
.A2(n_3403),
.B1(n_3433),
.B2(n_3393),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3408),
.B(n_3436),
.Y(n_3869)
);

OAI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3428),
.A2(n_3443),
.B(n_3204),
.Y(n_3870)
);

OAI21x1_ASAP7_75t_L g3871 ( 
.A1(n_3395),
.A2(n_3474),
.B(n_3414),
.Y(n_3871)
);

CKINVDCx20_ASAP7_75t_R g3872 ( 
.A(n_3136),
.Y(n_3872)
);

AOI22xp33_ASAP7_75t_L g3873 ( 
.A1(n_3463),
.A2(n_3231),
.B1(n_3301),
.B2(n_3284),
.Y(n_3873)
);

CKINVDCx5p33_ASAP7_75t_R g3874 ( 
.A(n_3175),
.Y(n_3874)
);

NAND3xp33_ASAP7_75t_L g3875 ( 
.A(n_3463),
.B(n_3080),
.C(n_3169),
.Y(n_3875)
);

AND2x4_ASAP7_75t_L g3876 ( 
.A(n_3365),
.B(n_3374),
.Y(n_3876)
);

OAI21x1_ASAP7_75t_L g3877 ( 
.A1(n_3395),
.A2(n_3474),
.B(n_3414),
.Y(n_3877)
);

AOI21xp5_ASAP7_75t_SL g3878 ( 
.A1(n_3285),
.A2(n_3292),
.B(n_3215),
.Y(n_3878)
);

OAI22xp5_ASAP7_75t_L g3879 ( 
.A1(n_3247),
.A2(n_3433),
.B1(n_3393),
.B2(n_3353),
.Y(n_3879)
);

AO21x2_ASAP7_75t_L g3880 ( 
.A1(n_3392),
.A2(n_3378),
.B(n_3365),
.Y(n_3880)
);

BUFx2_ASAP7_75t_SL g3881 ( 
.A(n_3215),
.Y(n_3881)
);

AOI22xp33_ASAP7_75t_L g3882 ( 
.A1(n_3231),
.A2(n_3284),
.B1(n_3330),
.B2(n_3301),
.Y(n_3882)
);

OAI21x1_ASAP7_75t_L g3883 ( 
.A1(n_3407),
.A2(n_3359),
.B(n_3350),
.Y(n_3883)
);

OAI21x1_ASAP7_75t_L g3884 ( 
.A1(n_3350),
.A2(n_3376),
.B(n_3359),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3408),
.B(n_3436),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3312),
.B(n_3325),
.Y(n_3886)
);

AND2x2_ASAP7_75t_L g3887 ( 
.A(n_3312),
.B(n_3325),
.Y(n_3887)
);

O2A1O1Ixp33_ASAP7_75t_L g3888 ( 
.A1(n_3183),
.A2(n_3205),
.B(n_3246),
.C(n_3204),
.Y(n_3888)
);

INVx8_ASAP7_75t_L g3889 ( 
.A(n_3237),
.Y(n_3889)
);

BUFx4f_ASAP7_75t_SL g3890 ( 
.A(n_3219),
.Y(n_3890)
);

OAI22xp33_ASAP7_75t_L g3891 ( 
.A1(n_3394),
.A2(n_3403),
.B1(n_3433),
.B2(n_3393),
.Y(n_3891)
);

CKINVDCx20_ASAP7_75t_R g3892 ( 
.A(n_3156),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3453),
.B(n_3388),
.Y(n_3893)
);

OAI22xp5_ASAP7_75t_L g3894 ( 
.A1(n_3433),
.A2(n_3040),
.B1(n_3030),
.B2(n_3089),
.Y(n_3894)
);

INVx3_ASAP7_75t_L g3895 ( 
.A(n_3483),
.Y(n_3895)
);

AND2x4_ASAP7_75t_L g3896 ( 
.A(n_3365),
.B(n_3374),
.Y(n_3896)
);

NOR2x1_ASAP7_75t_L g3897 ( 
.A(n_3471),
.B(n_3478),
.Y(n_3897)
);

AOI22xp33_ASAP7_75t_SL g3898 ( 
.A1(n_3176),
.A2(n_3468),
.B1(n_3485),
.B2(n_3254),
.Y(n_3898)
);

BUFx2_ASAP7_75t_L g3899 ( 
.A(n_3789),
.Y(n_3899)
);

NAND2x1p5_ASAP7_75t_L g3900 ( 
.A(n_3687),
.B(n_3379),
.Y(n_3900)
);

AOI22xp33_ASAP7_75t_L g3901 ( 
.A1(n_3508),
.A2(n_3071),
.B1(n_3069),
.B2(n_3272),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3795),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3752),
.Y(n_3903)
);

AOI21x1_ASAP7_75t_L g3904 ( 
.A1(n_3543),
.A2(n_3323),
.B(n_3309),
.Y(n_3904)
);

AND2x4_ASAP7_75t_L g3905 ( 
.A(n_3668),
.B(n_3365),
.Y(n_3905)
);

INVxp33_ASAP7_75t_L g3906 ( 
.A(n_3651),
.Y(n_3906)
);

INVx5_ASAP7_75t_L g3907 ( 
.A(n_3524),
.Y(n_3907)
);

AOI22xp5_ASAP7_75t_L g3908 ( 
.A1(n_3529),
.A2(n_3468),
.B1(n_3477),
.B2(n_3333),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3752),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3752),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3752),
.Y(n_3911)
);

OAI21x1_ASAP7_75t_L g3912 ( 
.A1(n_3735),
.A2(n_3442),
.B(n_3483),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3752),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3795),
.Y(n_3914)
);

OAI22xp33_ASAP7_75t_L g3915 ( 
.A1(n_3537),
.A2(n_3810),
.B1(n_3559),
.B2(n_3562),
.Y(n_3915)
);

AOI22xp33_ASAP7_75t_L g3916 ( 
.A1(n_3488),
.A2(n_3069),
.B1(n_3284),
.B2(n_3231),
.Y(n_3916)
);

OAI22xp5_ASAP7_75t_L g3917 ( 
.A1(n_3491),
.A2(n_3040),
.B1(n_3295),
.B2(n_3296),
.Y(n_3917)
);

BUFx10_ASAP7_75t_L g3918 ( 
.A(n_3857),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3771),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3723),
.B(n_3345),
.Y(n_3920)
);

INVx2_ASAP7_75t_L g3921 ( 
.A(n_3795),
.Y(n_3921)
);

AOI22xp33_ASAP7_75t_L g3922 ( 
.A1(n_3571),
.A2(n_3284),
.B1(n_3301),
.B2(n_3231),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3795),
.Y(n_3923)
);

INVx3_ASAP7_75t_L g3924 ( 
.A(n_3812),
.Y(n_3924)
);

OAI22xp5_ASAP7_75t_L g3925 ( 
.A1(n_3576),
.A2(n_3295),
.B1(n_3335),
.B2(n_3296),
.Y(n_3925)
);

OR2x6_ASAP7_75t_L g3926 ( 
.A(n_3524),
.B(n_3231),
.Y(n_3926)
);

OA21x2_ASAP7_75t_L g3927 ( 
.A1(n_3694),
.A2(n_3192),
.B(n_3169),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3752),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3781),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_3778),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3781),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3723),
.B(n_3192),
.Y(n_3932)
);

BUFx12f_ASAP7_75t_L g3933 ( 
.A(n_3552),
.Y(n_3933)
);

OAI21x1_ASAP7_75t_L g3934 ( 
.A1(n_3735),
.A2(n_3442),
.B(n_3486),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3781),
.Y(n_3935)
);

AOI22xp33_ASAP7_75t_L g3936 ( 
.A1(n_3529),
.A2(n_3301),
.B1(n_3330),
.B2(n_3442),
.Y(n_3936)
);

HB1xp67_ASAP7_75t_L g3937 ( 
.A(n_3528),
.Y(n_3937)
);

INVxp67_ASAP7_75t_L g3938 ( 
.A(n_3729),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3778),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3778),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3771),
.Y(n_3941)
);

BUFx8_ASAP7_75t_SL g3942 ( 
.A(n_3552),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3778),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3581),
.Y(n_3944)
);

OAI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3537),
.A2(n_3029),
.B1(n_3190),
.B2(n_3037),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3781),
.Y(n_3946)
);

NAND2x1p5_ASAP7_75t_L g3947 ( 
.A(n_3687),
.B(n_3379),
.Y(n_3947)
);

AOI22xp33_ASAP7_75t_SL g3948 ( 
.A1(n_3810),
.A2(n_3252),
.B1(n_3254),
.B2(n_3259),
.Y(n_3948)
);

HB1xp67_ASAP7_75t_L g3949 ( 
.A(n_3532),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3581),
.Y(n_3950)
);

CKINVDCx5p33_ASAP7_75t_R g3951 ( 
.A(n_3711),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3489),
.B(n_3453),
.Y(n_3952)
);

INVx6_ASAP7_75t_L g3953 ( 
.A(n_3552),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_3489),
.B(n_3216),
.Y(n_3954)
);

INVx3_ASAP7_75t_SL g3955 ( 
.A(n_3777),
.Y(n_3955)
);

AOI22xp33_ASAP7_75t_L g3956 ( 
.A1(n_3580),
.A2(n_3330),
.B1(n_3301),
.B2(n_3442),
.Y(n_3956)
);

BUFx6f_ASAP7_75t_L g3957 ( 
.A(n_3764),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3781),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3781),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3717),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3581),
.Y(n_3961)
);

OAI21x1_ASAP7_75t_L g3962 ( 
.A1(n_3740),
.A2(n_3486),
.B(n_3404),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3717),
.Y(n_3963)
);

HB1xp67_ASAP7_75t_L g3964 ( 
.A(n_3772),
.Y(n_3964)
);

AOI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_3505),
.A2(n_3292),
.B(n_3285),
.Y(n_3965)
);

AND2x4_ASAP7_75t_L g3966 ( 
.A(n_3668),
.B(n_3876),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3717),
.Y(n_3967)
);

NAND2x1p5_ASAP7_75t_L g3968 ( 
.A(n_3687),
.B(n_3379),
.Y(n_3968)
);

INVx3_ASAP7_75t_L g3969 ( 
.A(n_3812),
.Y(n_3969)
);

HB1xp67_ASAP7_75t_L g3970 ( 
.A(n_3804),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3581),
.Y(n_3971)
);

INVx2_ASAP7_75t_SL g3972 ( 
.A(n_3789),
.Y(n_3972)
);

OR2x2_ASAP7_75t_L g3973 ( 
.A(n_3751),
.B(n_3216),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3771),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3771),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3717),
.Y(n_3976)
);

OAI21x1_ASAP7_75t_L g3977 ( 
.A1(n_3740),
.A2(n_3486),
.B(n_3404),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3765),
.Y(n_3978)
);

CKINVDCx5p33_ASAP7_75t_R g3979 ( 
.A(n_3739),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3753),
.B(n_3217),
.Y(n_3980)
);

BUFx2_ASAP7_75t_L g3981 ( 
.A(n_3789),
.Y(n_3981)
);

INVx4_ASAP7_75t_L g3982 ( 
.A(n_3653),
.Y(n_3982)
);

OA21x2_ASAP7_75t_L g3983 ( 
.A1(n_3694),
.A2(n_3218),
.B(n_3217),
.Y(n_3983)
);

AOI21x1_ASAP7_75t_L g3984 ( 
.A1(n_3543),
.A2(n_3240),
.B(n_3218),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3717),
.Y(n_3985)
);

INVx1_ASAP7_75t_SL g3986 ( 
.A(n_3501),
.Y(n_3986)
);

BUFx2_ASAP7_75t_L g3987 ( 
.A(n_3707),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3502),
.B(n_3621),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_3717),
.Y(n_3989)
);

OAI22xp5_ASAP7_75t_L g3990 ( 
.A1(n_3560),
.A2(n_3526),
.B1(n_3518),
.B2(n_3504),
.Y(n_3990)
);

NAND2x1p5_ASAP7_75t_L g3991 ( 
.A(n_3687),
.B(n_3732),
.Y(n_3991)
);

AO21x2_ASAP7_75t_L g3992 ( 
.A1(n_3672),
.A2(n_3310),
.B(n_3268),
.Y(n_3992)
);

INVx2_ASAP7_75t_L g3993 ( 
.A(n_3765),
.Y(n_3993)
);

INVx3_ASAP7_75t_L g3994 ( 
.A(n_3812),
.Y(n_3994)
);

INVx2_ASAP7_75t_L g3995 ( 
.A(n_3765),
.Y(n_3995)
);

AND2x2_ASAP7_75t_L g3996 ( 
.A(n_3753),
.B(n_3240),
.Y(n_3996)
);

OAI21x1_ASAP7_75t_L g3997 ( 
.A1(n_3734),
.A2(n_3720),
.B(n_3715),
.Y(n_3997)
);

NAND2x1p5_ASAP7_75t_L g3998 ( 
.A(n_3732),
.B(n_3379),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3765),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3738),
.Y(n_4000)
);

INVx4_ASAP7_75t_L g4001 ( 
.A(n_3653),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3855),
.Y(n_4002)
);

BUFx3_ASAP7_75t_L g4003 ( 
.A(n_3653),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3855),
.Y(n_4004)
);

INVx2_ASAP7_75t_L g4005 ( 
.A(n_3738),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3855),
.Y(n_4006)
);

INVx6_ASAP7_75t_L g4007 ( 
.A(n_3763),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_L g4008 ( 
.A(n_3502),
.B(n_3183),
.Y(n_4008)
);

BUFx12f_ASAP7_75t_L g4009 ( 
.A(n_3567),
.Y(n_4009)
);

AOI21x1_ASAP7_75t_L g4010 ( 
.A1(n_3672),
.A2(n_3246),
.B(n_3205),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3490),
.Y(n_4011)
);

AOI22xp5_ASAP7_75t_L g4012 ( 
.A1(n_3580),
.A2(n_3477),
.B1(n_3333),
.B2(n_3363),
.Y(n_4012)
);

NAND2x1p5_ASAP7_75t_L g4013 ( 
.A(n_3767),
.B(n_3379),
.Y(n_4013)
);

INVx8_ASAP7_75t_L g4014 ( 
.A(n_3632),
.Y(n_4014)
);

BUFx6f_ASAP7_75t_L g4015 ( 
.A(n_3764),
.Y(n_4015)
);

INVx1_ASAP7_75t_SL g4016 ( 
.A(n_3749),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3490),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3495),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3738),
.Y(n_4019)
);

INVxp67_ASAP7_75t_SL g4020 ( 
.A(n_3638),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3495),
.Y(n_4021)
);

NOR2xp33_ASAP7_75t_R g4022 ( 
.A(n_3589),
.B(n_3399),
.Y(n_4022)
);

AND2x2_ASAP7_75t_L g4023 ( 
.A(n_3835),
.B(n_3396),
.Y(n_4023)
);

INVx3_ASAP7_75t_L g4024 ( 
.A(n_3812),
.Y(n_4024)
);

BUFx2_ASAP7_75t_L g4025 ( 
.A(n_3707),
.Y(n_4025)
);

INVx2_ASAP7_75t_L g4026 ( 
.A(n_3738),
.Y(n_4026)
);

AOI21x1_ASAP7_75t_L g4027 ( 
.A1(n_3546),
.A2(n_3830),
.B(n_3680),
.Y(n_4027)
);

AND2x2_ASAP7_75t_L g4028 ( 
.A(n_3835),
.B(n_3396),
.Y(n_4028)
);

BUFx2_ASAP7_75t_L g4029 ( 
.A(n_3707),
.Y(n_4029)
);

CKINVDCx20_ASAP7_75t_R g4030 ( 
.A(n_3521),
.Y(n_4030)
);

OR2x2_ASAP7_75t_L g4031 ( 
.A(n_3751),
.B(n_3053),
.Y(n_4031)
);

INVx3_ASAP7_75t_L g4032 ( 
.A(n_3821),
.Y(n_4032)
);

HB1xp67_ASAP7_75t_L g4033 ( 
.A(n_3819),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3792),
.Y(n_4034)
);

INVx2_ASAP7_75t_L g4035 ( 
.A(n_3792),
.Y(n_4035)
);

AOI22xp33_ASAP7_75t_L g4036 ( 
.A1(n_3530),
.A2(n_3620),
.B1(n_3559),
.B2(n_3586),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3498),
.Y(n_4037)
);

CKINVDCx20_ASAP7_75t_R g4038 ( 
.A(n_3538),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3498),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3506),
.Y(n_4040)
);

INVx4_ASAP7_75t_L g4041 ( 
.A(n_3632),
.Y(n_4041)
);

BUFx3_ASAP7_75t_L g4042 ( 
.A(n_3759),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3506),
.Y(n_4043)
);

BUFx6f_ASAP7_75t_L g4044 ( 
.A(n_3764),
.Y(n_4044)
);

BUFx6f_ASAP7_75t_L g4045 ( 
.A(n_3768),
.Y(n_4045)
);

BUFx2_ASAP7_75t_L g4046 ( 
.A(n_3707),
.Y(n_4046)
);

INVx2_ASAP7_75t_L g4047 ( 
.A(n_3792),
.Y(n_4047)
);

AOI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3701),
.A2(n_3330),
.B1(n_3300),
.B2(n_3037),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3792),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3511),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_3730),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3511),
.Y(n_4052)
);

OAI21xp5_ASAP7_75t_L g4053 ( 
.A1(n_3504),
.A2(n_3099),
.B(n_3053),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3512),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3512),
.Y(n_4055)
);

OAI21xp5_ASAP7_75t_SL g4056 ( 
.A1(n_3548),
.A2(n_3140),
.B(n_3119),
.Y(n_4056)
);

OAI21xp5_ASAP7_75t_L g4057 ( 
.A1(n_3493),
.A2(n_3099),
.B(n_3119),
.Y(n_4057)
);

OAI21x1_ASAP7_75t_L g4058 ( 
.A1(n_3734),
.A2(n_3404),
.B(n_3397),
.Y(n_4058)
);

OAI22xp33_ASAP7_75t_L g4059 ( 
.A1(n_3588),
.A2(n_3029),
.B1(n_3190),
.B2(n_3037),
.Y(n_4059)
);

AOI22xp33_ASAP7_75t_SL g4060 ( 
.A1(n_3813),
.A2(n_3252),
.B1(n_3254),
.B2(n_3259),
.Y(n_4060)
);

AOI22xp33_ASAP7_75t_L g4061 ( 
.A1(n_3701),
.A2(n_3666),
.B1(n_3569),
.B2(n_3813),
.Y(n_4061)
);

INVx2_ASAP7_75t_SL g4062 ( 
.A(n_3731),
.Y(n_4062)
);

AND2x2_ASAP7_75t_L g4063 ( 
.A(n_3837),
.B(n_3396),
.Y(n_4063)
);

INVxp33_ASAP7_75t_L g4064 ( 
.A(n_3803),
.Y(n_4064)
);

INVx3_ASAP7_75t_L g4065 ( 
.A(n_3821),
.Y(n_4065)
);

INVx3_ASAP7_75t_L g4066 ( 
.A(n_3821),
.Y(n_4066)
);

AND2x2_ASAP7_75t_L g4067 ( 
.A(n_3837),
.B(n_3106),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3513),
.Y(n_4068)
);

AND2x2_ASAP7_75t_L g4069 ( 
.A(n_3773),
.B(n_3106),
.Y(n_4069)
);

OAI21x1_ASAP7_75t_L g4070 ( 
.A1(n_3715),
.A2(n_3397),
.B(n_3470),
.Y(n_4070)
);

HB1xp67_ASAP7_75t_L g4071 ( 
.A(n_3590),
.Y(n_4071)
);

HB1xp67_ASAP7_75t_L g4072 ( 
.A(n_3593),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3513),
.Y(n_4073)
);

AND2x4_ASAP7_75t_L g4074 ( 
.A(n_3668),
.B(n_3259),
.Y(n_4074)
);

AOI21x1_ASAP7_75t_L g4075 ( 
.A1(n_3830),
.A2(n_3310),
.B(n_3268),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3831),
.Y(n_4076)
);

INVx2_ASAP7_75t_L g4077 ( 
.A(n_3831),
.Y(n_4077)
);

NAND2xp33_ASAP7_75t_SL g4078 ( 
.A(n_3554),
.B(n_3117),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_3569),
.A2(n_3330),
.B1(n_3342),
.B2(n_3037),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3831),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3831),
.Y(n_4081)
);

HB1xp67_ASAP7_75t_L g4082 ( 
.A(n_3867),
.Y(n_4082)
);

OAI22xp33_ASAP7_75t_L g4083 ( 
.A1(n_3588),
.A2(n_3029),
.B1(n_3190),
.B2(n_3037),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3515),
.Y(n_4084)
);

INVx2_ASAP7_75t_SL g4085 ( 
.A(n_3731),
.Y(n_4085)
);

INVx3_ASAP7_75t_L g4086 ( 
.A(n_3821),
.Y(n_4086)
);

OAI22xp5_ASAP7_75t_L g4087 ( 
.A1(n_3548),
.A2(n_3295),
.B1(n_3335),
.B2(n_3089),
.Y(n_4087)
);

INVx6_ASAP7_75t_L g4088 ( 
.A(n_3763),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_3621),
.B(n_3140),
.Y(n_4089)
);

BUFx2_ASAP7_75t_L g4090 ( 
.A(n_3731),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3515),
.Y(n_4091)
);

OAI21x1_ASAP7_75t_L g4092 ( 
.A1(n_3720),
.A2(n_3397),
.B(n_3470),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_3516),
.Y(n_4093)
);

INVx2_ASAP7_75t_L g4094 ( 
.A(n_3497),
.Y(n_4094)
);

OAI21xp5_ASAP7_75t_L g4095 ( 
.A1(n_3604),
.A2(n_3292),
.B(n_3285),
.Y(n_4095)
);

BUFx6f_ASAP7_75t_SL g4096 ( 
.A(n_3557),
.Y(n_4096)
);

HB1xp67_ASAP7_75t_L g4097 ( 
.A(n_3725),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3497),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3516),
.Y(n_4099)
);

BUFx4f_ASAP7_75t_SL g4100 ( 
.A(n_3872),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3523),
.Y(n_4101)
);

INVx3_ASAP7_75t_L g4102 ( 
.A(n_3829),
.Y(n_4102)
);

BUFx8_ASAP7_75t_L g4103 ( 
.A(n_3759),
.Y(n_4103)
);

HB1xp67_ASAP7_75t_L g4104 ( 
.A(n_3725),
.Y(n_4104)
);

BUFx8_ASAP7_75t_L g4105 ( 
.A(n_3759),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_3497),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3643),
.B(n_3406),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_SL g4108 ( 
.A1(n_3607),
.A2(n_3252),
.B1(n_3262),
.B2(n_3412),
.Y(n_4108)
);

OAI22xp33_ASAP7_75t_L g4109 ( 
.A1(n_3695),
.A2(n_3029),
.B1(n_3190),
.B2(n_3037),
.Y(n_4109)
);

HB1xp67_ASAP7_75t_L g4110 ( 
.A(n_3727),
.Y(n_4110)
);

AND2x2_ASAP7_75t_L g4111 ( 
.A(n_3773),
.B(n_3106),
.Y(n_4111)
);

AO21x2_ASAP7_75t_L g4112 ( 
.A1(n_3555),
.A2(n_3310),
.B(n_3268),
.Y(n_4112)
);

AOI22xp33_ASAP7_75t_L g4113 ( 
.A1(n_3555),
.A2(n_3029),
.B1(n_3190),
.B2(n_3037),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3523),
.Y(n_4114)
);

INVx2_ASAP7_75t_L g4115 ( 
.A(n_3730),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3533),
.Y(n_4116)
);

AOI22xp33_ASAP7_75t_L g4117 ( 
.A1(n_3599),
.A2(n_3029),
.B1(n_3344),
.B2(n_3342),
.Y(n_4117)
);

BUFx2_ASAP7_75t_L g4118 ( 
.A(n_3731),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_3730),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3533),
.Y(n_4120)
);

AO21x1_ASAP7_75t_L g4121 ( 
.A1(n_3833),
.A2(n_3425),
.B(n_3424),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3540),
.Y(n_4122)
);

BUFx3_ASAP7_75t_L g4123 ( 
.A(n_3632),
.Y(n_4123)
);

INVx2_ASAP7_75t_L g4124 ( 
.A(n_3507),
.Y(n_4124)
);

BUFx2_ASAP7_75t_SL g4125 ( 
.A(n_3630),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3540),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3802),
.B(n_3106),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3542),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3542),
.Y(n_4129)
);

AOI22xp33_ASAP7_75t_SL g4130 ( 
.A1(n_3607),
.A2(n_3262),
.B1(n_3412),
.B2(n_3313),
.Y(n_4130)
);

INVx2_ASAP7_75t_L g4131 ( 
.A(n_3507),
.Y(n_4131)
);

AOI222xp33_ASAP7_75t_L g4132 ( 
.A1(n_3487),
.A2(n_3262),
.B1(n_3412),
.B2(n_3383),
.C1(n_3389),
.C2(n_3326),
.Y(n_4132)
);

OAI21x1_ASAP7_75t_SL g4133 ( 
.A1(n_3808),
.A2(n_3425),
.B(n_3424),
.Y(n_4133)
);

CKINVDCx20_ASAP7_75t_R g4134 ( 
.A(n_3589),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_3802),
.B(n_3106),
.Y(n_4135)
);

HB1xp67_ASAP7_75t_L g4136 ( 
.A(n_3727),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3544),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_3507),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_3544),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_3545),
.Y(n_4140)
);

AOI22xp33_ASAP7_75t_SL g4141 ( 
.A1(n_3657),
.A2(n_3321),
.B1(n_3313),
.B2(n_3316),
.Y(n_4141)
);

BUFx6f_ASAP7_75t_L g4142 ( 
.A(n_3768),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3545),
.Y(n_4143)
);

AOI22xp33_ASAP7_75t_L g4144 ( 
.A1(n_3702),
.A2(n_3029),
.B1(n_3344),
.B2(n_3342),
.Y(n_4144)
);

INVxp67_ASAP7_75t_L g4145 ( 
.A(n_3519),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_3517),
.Y(n_4146)
);

HB1xp67_ASAP7_75t_L g4147 ( 
.A(n_3783),
.Y(n_4147)
);

HB1xp67_ASAP7_75t_L g4148 ( 
.A(n_3783),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3551),
.Y(n_4149)
);

OAI21x1_ASAP7_75t_L g4150 ( 
.A1(n_3726),
.A2(n_3470),
.B(n_3416),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_3551),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_3565),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3565),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3566),
.Y(n_4154)
);

HB1xp67_ASAP7_75t_L g4155 ( 
.A(n_3814),
.Y(n_4155)
);

OR2x2_ASAP7_75t_L g4156 ( 
.A(n_3758),
.B(n_3210),
.Y(n_4156)
);

INVx4_ASAP7_75t_L g4157 ( 
.A(n_3632),
.Y(n_4157)
);

BUFx12f_ASAP7_75t_L g4158 ( 
.A(n_3710),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_3643),
.B(n_3210),
.Y(n_4159)
);

BUFx3_ASAP7_75t_L g4160 ( 
.A(n_3632),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3566),
.Y(n_4161)
);

AOI21x1_ASAP7_75t_L g4162 ( 
.A1(n_3680),
.A2(n_3310),
.B(n_3268),
.Y(n_4162)
);

HB1xp67_ASAP7_75t_L g4163 ( 
.A(n_3814),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3517),
.Y(n_4164)
);

AOI22xp33_ASAP7_75t_L g4165 ( 
.A1(n_3487),
.A2(n_3190),
.B1(n_3308),
.B2(n_3307),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_3517),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3570),
.Y(n_4167)
);

BUFx12f_ASAP7_75t_L g4168 ( 
.A(n_3748),
.Y(n_4168)
);

BUFx3_ASAP7_75t_L g4169 ( 
.A(n_3630),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_3525),
.Y(n_4170)
);

BUFx2_ASAP7_75t_L g4171 ( 
.A(n_3766),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_3525),
.Y(n_4172)
);

BUFx6f_ASAP7_75t_L g4173 ( 
.A(n_3768),
.Y(n_4173)
);

BUFx3_ASAP7_75t_L g4174 ( 
.A(n_3763),
.Y(n_4174)
);

CKINVDCx6p67_ASAP7_75t_R g4175 ( 
.A(n_3617),
.Y(n_4175)
);

INVx3_ASAP7_75t_L g4176 ( 
.A(n_3829),
.Y(n_4176)
);

OA21x2_ASAP7_75t_L g4177 ( 
.A1(n_3703),
.A2(n_3355),
.B(n_3416),
.Y(n_4177)
);

AOI22xp33_ASAP7_75t_L g4178 ( 
.A1(n_3592),
.A2(n_3190),
.B1(n_3308),
.B2(n_3307),
.Y(n_4178)
);

INVx3_ASAP7_75t_L g4179 ( 
.A(n_3829),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_3570),
.Y(n_4180)
);

BUFx3_ASAP7_75t_L g4181 ( 
.A(n_3763),
.Y(n_4181)
);

AND2x4_ASAP7_75t_L g4182 ( 
.A(n_3668),
.B(n_3172),
.Y(n_4182)
);

AOI22xp5_ASAP7_75t_L g4183 ( 
.A1(n_3647),
.A2(n_3477),
.B1(n_3358),
.B2(n_3363),
.Y(n_4183)
);

HB1xp67_ASAP7_75t_L g4184 ( 
.A(n_3817),
.Y(n_4184)
);

NAND2x1p5_ASAP7_75t_L g4185 ( 
.A(n_3767),
.B(n_3379),
.Y(n_4185)
);

INVx3_ASAP7_75t_L g4186 ( 
.A(n_3829),
.Y(n_4186)
);

CKINVDCx11_ASAP7_75t_R g4187 ( 
.A(n_3892),
.Y(n_4187)
);

AND2x2_ASAP7_75t_L g4188 ( 
.A(n_3618),
.B(n_3172),
.Y(n_4188)
);

OAI22xp5_ASAP7_75t_L g4189 ( 
.A1(n_3536),
.A2(n_3089),
.B1(n_3097),
.B2(n_3219),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_3572),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_3572),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_3577),
.Y(n_4192)
);

CKINVDCx5p33_ASAP7_75t_R g4193 ( 
.A(n_3874),
.Y(n_4193)
);

INVxp33_ASAP7_75t_L g4194 ( 
.A(n_3788),
.Y(n_4194)
);

BUFx2_ASAP7_75t_L g4195 ( 
.A(n_3766),
.Y(n_4195)
);

HB1xp67_ASAP7_75t_L g4196 ( 
.A(n_3817),
.Y(n_4196)
);

AOI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_3657),
.A2(n_3611),
.B1(n_3833),
.B2(n_3595),
.Y(n_4197)
);

INVx3_ASAP7_75t_L g4198 ( 
.A(n_3876),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_3577),
.Y(n_4199)
);

AOI22xp33_ASAP7_75t_L g4200 ( 
.A1(n_3496),
.A2(n_3289),
.B1(n_3320),
.B2(n_3308),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_3578),
.Y(n_4201)
);

BUFx8_ASAP7_75t_L g4202 ( 
.A(n_3557),
.Y(n_4202)
);

AOI22xp5_ASAP7_75t_L g4203 ( 
.A1(n_3647),
.A2(n_3363),
.B1(n_3358),
.B2(n_3047),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3578),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3579),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_3579),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_3618),
.B(n_3210),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_3582),
.Y(n_4208)
);

BUFx3_ASAP7_75t_L g4209 ( 
.A(n_3770),
.Y(n_4209)
);

AOI22xp33_ASAP7_75t_L g4210 ( 
.A1(n_3496),
.A2(n_3308),
.B1(n_3269),
.B2(n_3275),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3582),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_3629),
.B(n_3232),
.Y(n_4212)
);

AND2x4_ASAP7_75t_L g4213 ( 
.A(n_3668),
.B(n_3172),
.Y(n_4213)
);

INVx3_ASAP7_75t_L g4214 ( 
.A(n_3876),
.Y(n_4214)
);

INVx3_ASAP7_75t_L g4215 ( 
.A(n_3876),
.Y(n_4215)
);

AND2x2_ASAP7_75t_L g4216 ( 
.A(n_3629),
.B(n_3645),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_3730),
.Y(n_4217)
);

BUFx3_ASAP7_75t_L g4218 ( 
.A(n_3770),
.Y(n_4218)
);

AOI22xp33_ASAP7_75t_L g4219 ( 
.A1(n_3496),
.A2(n_3308),
.B1(n_3269),
.B2(n_3275),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_3587),
.Y(n_4220)
);

INVx4_ASAP7_75t_L g4221 ( 
.A(n_3541),
.Y(n_4221)
);

BUFx3_ASAP7_75t_L g4222 ( 
.A(n_3770),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3587),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_3591),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3591),
.Y(n_4225)
);

OAI21xp33_ASAP7_75t_L g4226 ( 
.A1(n_3558),
.A2(n_3585),
.B(n_3713),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_3645),
.B(n_3174),
.Y(n_4227)
);

AOI22xp33_ASAP7_75t_L g4228 ( 
.A1(n_3496),
.A2(n_3308),
.B1(n_3269),
.B2(n_3275),
.Y(n_4228)
);

HB1xp67_ASAP7_75t_L g4229 ( 
.A(n_3848),
.Y(n_4229)
);

AOI22xp33_ASAP7_75t_L g4230 ( 
.A1(n_3698),
.A2(n_3062),
.B1(n_3320),
.B2(n_3307),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_3596),
.Y(n_4231)
);

HB1xp67_ASAP7_75t_L g4232 ( 
.A(n_3848),
.Y(n_4232)
);

AOI22xp33_ASAP7_75t_SL g4233 ( 
.A1(n_3524),
.A2(n_3313),
.B1(n_3321),
.B2(n_3316),
.Y(n_4233)
);

CKINVDCx11_ASAP7_75t_R g4234 ( 
.A(n_3554),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_3654),
.B(n_3658),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_3596),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_3654),
.B(n_3174),
.Y(n_4237)
);

NAND2x1p5_ASAP7_75t_L g4238 ( 
.A(n_3769),
.B(n_3379),
.Y(n_4238)
);

CKINVDCx6p67_ASAP7_75t_R g4239 ( 
.A(n_3554),
.Y(n_4239)
);

BUFx8_ASAP7_75t_L g4240 ( 
.A(n_3557),
.Y(n_4240)
);

BUFx6f_ASAP7_75t_L g4241 ( 
.A(n_3774),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_3492),
.A2(n_3062),
.B1(n_3320),
.B2(n_3307),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_3597),
.Y(n_4243)
);

OAI22xp5_ASAP7_75t_L g4244 ( 
.A1(n_3662),
.A2(n_3097),
.B1(n_3219),
.B2(n_3095),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3597),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_3598),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_3598),
.Y(n_4247)
);

BUFx12f_ASAP7_75t_L g4248 ( 
.A(n_3754),
.Y(n_4248)
);

OAI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_3677),
.A2(n_3097),
.B1(n_3095),
.B2(n_3113),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_3601),
.Y(n_4250)
);

INVx2_ASAP7_75t_SL g4251 ( 
.A(n_3766),
.Y(n_4251)
);

INVx2_ASAP7_75t_SL g4252 ( 
.A(n_3766),
.Y(n_4252)
);

OAI22xp5_ASAP7_75t_L g4253 ( 
.A1(n_3677),
.A2(n_3113),
.B1(n_3174),
.B2(n_3232),
.Y(n_4253)
);

OAI21x1_ASAP7_75t_L g4254 ( 
.A1(n_3726),
.A2(n_3470),
.B(n_3416),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_3658),
.B(n_3232),
.Y(n_4255)
);

AOI22xp33_ASAP7_75t_L g4256 ( 
.A1(n_3492),
.A2(n_3344),
.B1(n_3269),
.B2(n_3275),
.Y(n_4256)
);

BUFx2_ASAP7_75t_L g4257 ( 
.A(n_3811),
.Y(n_4257)
);

OA21x2_ASAP7_75t_L g4258 ( 
.A1(n_3703),
.A2(n_3355),
.B(n_3383),
.Y(n_4258)
);

CKINVDCx5p33_ASAP7_75t_R g4259 ( 
.A(n_3736),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3601),
.Y(n_4260)
);

INVx6_ASAP7_75t_L g4261 ( 
.A(n_3514),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_3622),
.Y(n_4262)
);

NAND2x1p5_ASAP7_75t_L g4263 ( 
.A(n_3769),
.B(n_3062),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3622),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_3623),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_3661),
.B(n_3340),
.Y(n_4266)
);

HB1xp67_ASAP7_75t_L g4267 ( 
.A(n_3553),
.Y(n_4267)
);

BUFx6f_ASAP7_75t_L g4268 ( 
.A(n_3774),
.Y(n_4268)
);

AOI22xp33_ASAP7_75t_L g4269 ( 
.A1(n_3492),
.A2(n_3344),
.B1(n_3269),
.B2(n_3275),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_3623),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_3628),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_3628),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_3633),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_3633),
.Y(n_4274)
);

BUFx2_ASAP7_75t_R g4275 ( 
.A(n_3603),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3636),
.Y(n_4276)
);

BUFx2_ASAP7_75t_L g4277 ( 
.A(n_3811),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_3636),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_3661),
.B(n_3340),
.Y(n_4279)
);

BUFx6f_ASAP7_75t_L g4280 ( 
.A(n_3774),
.Y(n_4280)
);

BUFx10_ASAP7_75t_L g4281 ( 
.A(n_3857),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_3660),
.B(n_3340),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_3641),
.Y(n_4283)
);

HB1xp67_ASAP7_75t_L g4284 ( 
.A(n_3758),
.Y(n_4284)
);

AOI22xp5_ASAP7_75t_L g4285 ( 
.A1(n_3568),
.A2(n_3358),
.B1(n_3363),
.B2(n_3047),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_3641),
.Y(n_4286)
);

BUFx3_ASAP7_75t_L g4287 ( 
.A(n_3603),
.Y(n_4287)
);

OR2x2_ASAP7_75t_L g4288 ( 
.A(n_3721),
.B(n_3383),
.Y(n_4288)
);

AOI22xp33_ASAP7_75t_SL g4289 ( 
.A1(n_3524),
.A2(n_3563),
.B1(n_3494),
.B2(n_3500),
.Y(n_4289)
);

BUFx12f_ASAP7_75t_L g4290 ( 
.A(n_3550),
.Y(n_4290)
);

OAI22xp5_ASAP7_75t_L g4291 ( 
.A1(n_3728),
.A2(n_3241),
.B1(n_3282),
.B2(n_3343),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_3642),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_3642),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_3644),
.Y(n_4294)
);

OAI22xp5_ASAP7_75t_L g4295 ( 
.A1(n_3535),
.A2(n_3241),
.B1(n_3343),
.B2(n_3046),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_3660),
.B(n_3343),
.Y(n_4296)
);

HB1xp67_ASAP7_75t_L g4297 ( 
.A(n_3852),
.Y(n_4297)
);

INVx2_ASAP7_75t_SL g4298 ( 
.A(n_3811),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_3644),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_3648),
.Y(n_4300)
);

INVx4_ASAP7_75t_L g4301 ( 
.A(n_3541),
.Y(n_4301)
);

OR2x2_ASAP7_75t_L g4302 ( 
.A(n_3721),
.B(n_3389),
.Y(n_4302)
);

OAI21x1_ASAP7_75t_L g4303 ( 
.A1(n_3860),
.A2(n_3280),
.B(n_3273),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_3648),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_3650),
.Y(n_4305)
);

BUFx3_ASAP7_75t_L g4306 ( 
.A(n_3603),
.Y(n_4306)
);

AND2x4_ASAP7_75t_L g4307 ( 
.A(n_3896),
.B(n_3354),
.Y(n_4307)
);

INVx6_ASAP7_75t_L g4308 ( 
.A(n_3514),
.Y(n_4308)
);

AOI21xp5_ASAP7_75t_L g4309 ( 
.A1(n_3614),
.A2(n_3478),
.B(n_3471),
.Y(n_4309)
);

AND2x2_ASAP7_75t_L g4310 ( 
.A(n_3886),
.B(n_3398),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_3650),
.Y(n_4311)
);

OAI22xp5_ASAP7_75t_L g4312 ( 
.A1(n_3787),
.A2(n_3046),
.B1(n_3142),
.B2(n_3075),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_3655),
.Y(n_4313)
);

OAI22xp5_ASAP7_75t_SL g4314 ( 
.A1(n_3787),
.A2(n_3796),
.B1(n_3746),
.B2(n_3875),
.Y(n_4314)
);

INVxp67_ASAP7_75t_L g4315 ( 
.A(n_3716),
.Y(n_4315)
);

OR2x6_ASAP7_75t_L g4316 ( 
.A(n_3524),
.B(n_3358),
.Y(n_4316)
);

AOI22xp33_ASAP7_75t_L g4317 ( 
.A1(n_3492),
.A2(n_3494),
.B1(n_3500),
.B2(n_3690),
.Y(n_4317)
);

BUFx8_ASAP7_75t_L g4318 ( 
.A(n_3605),
.Y(n_4318)
);

OAI21x1_ASAP7_75t_L g4319 ( 
.A1(n_3860),
.A2(n_3280),
.B(n_3273),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_3655),
.Y(n_4320)
);

CKINVDCx20_ASAP7_75t_R g4321 ( 
.A(n_3890),
.Y(n_4321)
);

BUFx10_ASAP7_75t_L g4322 ( 
.A(n_3857),
.Y(n_4322)
);

OAI21xp5_ASAP7_75t_SL g4323 ( 
.A1(n_3713),
.A2(n_3454),
.B(n_3452),
.Y(n_4323)
);

BUFx3_ASAP7_75t_L g4324 ( 
.A(n_3605),
.Y(n_4324)
);

INVxp33_ASAP7_75t_L g4325 ( 
.A(n_3534),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_3659),
.Y(n_4326)
);

AOI22xp33_ASAP7_75t_L g4327 ( 
.A1(n_3494),
.A2(n_3342),
.B1(n_3269),
.B2(n_3275),
.Y(n_4327)
);

AO21x1_ASAP7_75t_SL g4328 ( 
.A1(n_3558),
.A2(n_3585),
.B(n_3870),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_3659),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_3663),
.Y(n_4330)
);

INVx6_ASAP7_75t_L g4331 ( 
.A(n_3514),
.Y(n_4331)
);

OA21x2_ASAP7_75t_L g4332 ( 
.A1(n_3704),
.A2(n_3355),
.B(n_3389),
.Y(n_4332)
);

BUFx6f_ASAP7_75t_L g4333 ( 
.A(n_3605),
.Y(n_4333)
);

OAI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_3801),
.A2(n_3356),
.B(n_3354),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_3716),
.B(n_3459),
.Y(n_4335)
);

BUFx3_ASAP7_75t_L g4336 ( 
.A(n_3631),
.Y(n_4336)
);

HB1xp67_ASAP7_75t_L g4337 ( 
.A(n_3852),
.Y(n_4337)
);

HB1xp67_ASAP7_75t_L g4338 ( 
.A(n_3854),
.Y(n_4338)
);

OAI21x1_ASAP7_75t_L g4339 ( 
.A1(n_3866),
.A2(n_3280),
.B(n_3273),
.Y(n_4339)
);

BUFx10_ASAP7_75t_L g4340 ( 
.A(n_3857),
.Y(n_4340)
);

INVx1_ASAP7_75t_SL g4341 ( 
.A(n_3736),
.Y(n_4341)
);

CKINVDCx20_ASAP7_75t_R g4342 ( 
.A(n_3631),
.Y(n_4342)
);

BUFx8_ASAP7_75t_L g4343 ( 
.A(n_3631),
.Y(n_4343)
);

AOI21x1_ASAP7_75t_L g4344 ( 
.A1(n_3696),
.A2(n_3355),
.B(n_3358),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_3663),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_3886),
.B(n_3398),
.Y(n_4346)
);

AOI22xp33_ASAP7_75t_SL g4347 ( 
.A1(n_3563),
.A2(n_3316),
.B1(n_3321),
.B2(n_3356),
.Y(n_4347)
);

OAI21x1_ASAP7_75t_L g4348 ( 
.A1(n_3866),
.A2(n_3354),
.B(n_3356),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_3664),
.Y(n_4349)
);

OAI21x1_ASAP7_75t_L g4350 ( 
.A1(n_3871),
.A2(n_3294),
.B(n_3304),
.Y(n_4350)
);

INVx2_ASAP7_75t_SL g4351 ( 
.A(n_3811),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_3664),
.Y(n_4352)
);

AOI22xp33_ASAP7_75t_L g4353 ( 
.A1(n_3494),
.A2(n_3307),
.B1(n_3269),
.B2(n_3275),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_3675),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_3675),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_3682),
.Y(n_4356)
);

OA21x2_ASAP7_75t_L g4357 ( 
.A1(n_3704),
.A2(n_3452),
.B(n_3454),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_3682),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_3887),
.B(n_3522),
.Y(n_4359)
);

AOI22xp33_ASAP7_75t_SL g4360 ( 
.A1(n_3563),
.A2(n_3326),
.B1(n_3339),
.B2(n_3459),
.Y(n_4360)
);

AOI22xp33_ASAP7_75t_L g4361 ( 
.A1(n_3563),
.A2(n_3289),
.B1(n_3344),
.B2(n_3077),
.Y(n_4361)
);

BUFx12f_ASAP7_75t_L g4362 ( 
.A(n_3550),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_3887),
.B(n_3398),
.Y(n_4363)
);

OAI21x1_ASAP7_75t_L g4364 ( 
.A1(n_3871),
.A2(n_3304),
.B(n_3294),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_3686),
.Y(n_4365)
);

OAI22xp33_ASAP7_75t_L g4366 ( 
.A1(n_3563),
.A2(n_3289),
.B1(n_3300),
.B2(n_3307),
.Y(n_4366)
);

AND2x2_ASAP7_75t_L g4367 ( 
.A(n_3522),
.B(n_3398),
.Y(n_4367)
);

OA21x2_ASAP7_75t_L g4368 ( 
.A1(n_3705),
.A2(n_3452),
.B(n_3454),
.Y(n_4368)
);

AND2x4_ASAP7_75t_L g4369 ( 
.A(n_3896),
.B(n_3326),
.Y(n_4369)
);

NOR2xp33_ASAP7_75t_L g4370 ( 
.A(n_3799),
.B(n_3270),
.Y(n_4370)
);

AOI22xp33_ASAP7_75t_L g4371 ( 
.A1(n_3670),
.A2(n_3307),
.B1(n_3289),
.B2(n_3300),
.Y(n_4371)
);

AOI21x1_ASAP7_75t_L g4372 ( 
.A1(n_3696),
.A2(n_3363),
.B(n_3270),
.Y(n_4372)
);

BUFx8_ASAP7_75t_SL g4373 ( 
.A(n_3652),
.Y(n_4373)
);

BUFx2_ASAP7_75t_L g4374 ( 
.A(n_3897),
.Y(n_4374)
);

HB1xp67_ASAP7_75t_L g4375 ( 
.A(n_3854),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_3686),
.Y(n_4376)
);

OR2x6_ASAP7_75t_L g4377 ( 
.A(n_3878),
.B(n_3155),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_3689),
.Y(n_4378)
);

BUFx6f_ASAP7_75t_L g4379 ( 
.A(n_3652),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_3689),
.Y(n_4380)
);

CKINVDCx11_ASAP7_75t_R g4381 ( 
.A(n_3549),
.Y(n_4381)
);

AOI22xp33_ASAP7_75t_L g4382 ( 
.A1(n_3670),
.A2(n_3289),
.B1(n_3344),
.B2(n_3342),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_L g4383 ( 
.A(n_3640),
.B(n_3459),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_3691),
.Y(n_4384)
);

AOI21x1_ASAP7_75t_L g4385 ( 
.A1(n_3615),
.A2(n_3270),
.B(n_3080),
.Y(n_4385)
);

OAI21x1_ASAP7_75t_L g4386 ( 
.A1(n_3877),
.A2(n_3304),
.B(n_3294),
.Y(n_4386)
);

OA21x2_ASAP7_75t_L g4387 ( 
.A1(n_3705),
.A2(n_3452),
.B(n_3454),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_3691),
.Y(n_4388)
);

NAND2x1p5_ASAP7_75t_L g4389 ( 
.A(n_3776),
.B(n_3062),
.Y(n_4389)
);

OAI22xp33_ASAP7_75t_L g4390 ( 
.A1(n_3669),
.A2(n_3679),
.B1(n_3722),
.B2(n_3673),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_3693),
.Y(n_4391)
);

BUFx4f_ASAP7_75t_SL g4392 ( 
.A(n_3652),
.Y(n_4392)
);

AOI21x1_ASAP7_75t_L g4393 ( 
.A1(n_3615),
.A2(n_3080),
.B(n_3118),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_3693),
.Y(n_4394)
);

OAI21x1_ASAP7_75t_L g4395 ( 
.A1(n_3877),
.A2(n_3410),
.B(n_3339),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_SL g4396 ( 
.A(n_3613),
.B(n_3471),
.Y(n_4396)
);

AOI22xp33_ASAP7_75t_L g4397 ( 
.A1(n_3683),
.A2(n_3289),
.B1(n_3344),
.B2(n_3342),
.Y(n_4397)
);

AOI22xp33_ASAP7_75t_L g4398 ( 
.A1(n_3683),
.A2(n_3320),
.B1(n_3289),
.B2(n_3300),
.Y(n_4398)
);

NAND2x1p5_ASAP7_75t_L g4399 ( 
.A(n_3776),
.B(n_3062),
.Y(n_4399)
);

OAI22x1_ASAP7_75t_L g4400 ( 
.A1(n_3531),
.A2(n_3300),
.B1(n_3077),
.B2(n_3320),
.Y(n_4400)
);

AOI22xp33_ASAP7_75t_SL g4401 ( 
.A1(n_3638),
.A2(n_3339),
.B1(n_3405),
.B2(n_3320),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_3884),
.B(n_3305),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_3699),
.Y(n_4403)
);

AOI22xp33_ASAP7_75t_L g4404 ( 
.A1(n_3683),
.A2(n_3300),
.B1(n_3077),
.B2(n_3320),
.Y(n_4404)
);

NAND2x1p5_ASAP7_75t_L g4405 ( 
.A(n_3897),
.B(n_3062),
.Y(n_4405)
);

BUFx6f_ASAP7_75t_L g4406 ( 
.A(n_3665),
.Y(n_4406)
);

INVx3_ASAP7_75t_L g4407 ( 
.A(n_3896),
.Y(n_4407)
);

BUFx2_ASAP7_75t_L g4408 ( 
.A(n_3840),
.Y(n_4408)
);

CKINVDCx11_ASAP7_75t_R g4409 ( 
.A(n_3549),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_3699),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_3709),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_3709),
.Y(n_4412)
);

BUFx3_ASAP7_75t_L g4413 ( 
.A(n_3665),
.Y(n_4413)
);

BUFx2_ASAP7_75t_SL g4414 ( 
.A(n_3550),
.Y(n_4414)
);

OA21x2_ASAP7_75t_L g4415 ( 
.A1(n_3997),
.A2(n_3706),
.B(n_3676),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4011),
.Y(n_4416)
);

INVx3_ASAP7_75t_L g4417 ( 
.A(n_3927),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4011),
.Y(n_4418)
);

AND2x2_ASAP7_75t_L g4419 ( 
.A(n_3987),
.B(n_3884),
.Y(n_4419)
);

INVx2_ASAP7_75t_L g4420 ( 
.A(n_3944),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4017),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4017),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4018),
.Y(n_4423)
);

BUFx3_ASAP7_75t_L g4424 ( 
.A(n_3942),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4018),
.Y(n_4425)
);

INVx2_ASAP7_75t_L g4426 ( 
.A(n_3944),
.Y(n_4426)
);

INVx2_ASAP7_75t_L g4427 ( 
.A(n_3944),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4021),
.Y(n_4428)
);

INVx2_ASAP7_75t_L g4429 ( 
.A(n_3950),
.Y(n_4429)
);

OAI21x1_ASAP7_75t_L g4430 ( 
.A1(n_4075),
.A2(n_3859),
.B(n_3706),
.Y(n_4430)
);

INVx2_ASAP7_75t_SL g4431 ( 
.A(n_3953),
.Y(n_4431)
);

AO21x1_ASAP7_75t_SL g4432 ( 
.A1(n_4095),
.A2(n_4057),
.B(n_4089),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_3950),
.Y(n_4433)
);

AO21x1_ASAP7_75t_SL g4434 ( 
.A1(n_4053),
.A2(n_3870),
.B(n_3747),
.Y(n_4434)
);

INVx2_ASAP7_75t_L g4435 ( 
.A(n_3950),
.Y(n_4435)
);

NOR2xp33_ASAP7_75t_L g4436 ( 
.A(n_4175),
.B(n_3796),
.Y(n_4436)
);

INVx3_ASAP7_75t_L g4437 ( 
.A(n_3927),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_4021),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4037),
.Y(n_4439)
);

INVx3_ASAP7_75t_L g4440 ( 
.A(n_3927),
.Y(n_4440)
);

AOI22xp33_ASAP7_75t_L g4441 ( 
.A1(n_4036),
.A2(n_3683),
.B1(n_3692),
.B2(n_3531),
.Y(n_4441)
);

OAI21xp33_ASAP7_75t_SL g4442 ( 
.A1(n_4020),
.A2(n_3883),
.B(n_3780),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_3961),
.Y(n_4443)
);

OA21x2_ASAP7_75t_L g4444 ( 
.A1(n_3997),
.A2(n_3676),
.B(n_3782),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4037),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_3988),
.B(n_3827),
.Y(n_4446)
);

HB1xp67_ASAP7_75t_L g4447 ( 
.A(n_3937),
.Y(n_4447)
);

INVx2_ASAP7_75t_SL g4448 ( 
.A(n_3953),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_3987),
.B(n_3809),
.Y(n_4449)
);

INVx3_ASAP7_75t_L g4450 ( 
.A(n_3927),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4039),
.Y(n_4451)
);

HB1xp67_ASAP7_75t_L g4452 ( 
.A(n_3949),
.Y(n_4452)
);

AO21x1_ASAP7_75t_SL g4453 ( 
.A1(n_4197),
.A2(n_3801),
.B(n_3805),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_4039),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_3971),
.Y(n_4455)
);

INVxp67_ASAP7_75t_L g4456 ( 
.A(n_4267),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_4025),
.B(n_3809),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_3961),
.Y(n_4458)
);

INVx2_ASAP7_75t_L g4459 ( 
.A(n_3961),
.Y(n_4459)
);

INVx2_ASAP7_75t_SL g4460 ( 
.A(n_3953),
.Y(n_4460)
);

INVx3_ASAP7_75t_L g4461 ( 
.A(n_3983),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4040),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4040),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4043),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_L g4465 ( 
.A(n_4226),
.B(n_3828),
.Y(n_4465)
);

INVx1_ASAP7_75t_SL g4466 ( 
.A(n_4187),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4043),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4025),
.B(n_3809),
.Y(n_4468)
);

AO21x2_ASAP7_75t_L g4469 ( 
.A1(n_3960),
.A2(n_3864),
.B(n_3847),
.Y(n_4469)
);

HB1xp67_ASAP7_75t_L g4470 ( 
.A(n_3964),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_4226),
.B(n_3828),
.Y(n_4471)
);

OR2x2_ASAP7_75t_L g4472 ( 
.A(n_3952),
.B(n_3861),
.Y(n_4472)
);

INVx2_ASAP7_75t_SL g4473 ( 
.A(n_3953),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_3971),
.Y(n_4474)
);

AND2x2_ASAP7_75t_L g4475 ( 
.A(n_4029),
.B(n_3809),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4050),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_3971),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4050),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4052),
.Y(n_4479)
);

INVx2_ASAP7_75t_SL g4480 ( 
.A(n_3966),
.Y(n_4480)
);

BUFx3_ASAP7_75t_L g4481 ( 
.A(n_3933),
.Y(n_4481)
);

INVx2_ASAP7_75t_L g4482 ( 
.A(n_4051),
.Y(n_4482)
);

BUFx3_ASAP7_75t_L g4483 ( 
.A(n_3933),
.Y(n_4483)
);

OAI21x1_ASAP7_75t_L g4484 ( 
.A1(n_4075),
.A2(n_3859),
.B(n_3782),
.Y(n_4484)
);

CKINVDCx20_ASAP7_75t_R g4485 ( 
.A(n_4030),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_4051),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_4115),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4052),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4054),
.Y(n_4489)
);

HB1xp67_ASAP7_75t_L g4490 ( 
.A(n_3970),
.Y(n_4490)
);

INVx3_ASAP7_75t_L g4491 ( 
.A(n_3983),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4054),
.Y(n_4492)
);

OA21x2_ASAP7_75t_L g4493 ( 
.A1(n_4150),
.A2(n_3745),
.B(n_3750),
.Y(n_4493)
);

HB1xp67_ASAP7_75t_L g4494 ( 
.A(n_4033),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4055),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_4055),
.Y(n_4496)
);

O2A1O1Ixp33_ASAP7_75t_SL g4497 ( 
.A1(n_4341),
.A2(n_3719),
.B(n_3737),
.C(n_3865),
.Y(n_4497)
);

HB1xp67_ASAP7_75t_L g4498 ( 
.A(n_4082),
.Y(n_4498)
);

INVx1_ASAP7_75t_SL g4499 ( 
.A(n_4134),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_4068),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4029),
.B(n_3840),
.Y(n_4501)
);

OAI21x1_ASAP7_75t_L g4502 ( 
.A1(n_3984),
.A2(n_3780),
.B(n_3779),
.Y(n_4502)
);

AND2x4_ASAP7_75t_L g4503 ( 
.A(n_3907),
.B(n_3692),
.Y(n_4503)
);

INVxp67_ASAP7_75t_L g4504 ( 
.A(n_4071),
.Y(n_4504)
);

INVx2_ASAP7_75t_L g4505 ( 
.A(n_4115),
.Y(n_4505)
);

OAI21x1_ASAP7_75t_L g4506 ( 
.A1(n_3984),
.A2(n_3779),
.B(n_3714),
.Y(n_4506)
);

HB1xp67_ASAP7_75t_L g4507 ( 
.A(n_4072),
.Y(n_4507)
);

INVx2_ASAP7_75t_L g4508 ( 
.A(n_4119),
.Y(n_4508)
);

AND2x4_ASAP7_75t_SL g4509 ( 
.A(n_3918),
.B(n_3531),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4068),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4073),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_4097),
.B(n_3869),
.Y(n_4512)
);

INVx2_ASAP7_75t_L g4513 ( 
.A(n_4119),
.Y(n_4513)
);

BUFx12f_ASAP7_75t_L g4514 ( 
.A(n_4234),
.Y(n_4514)
);

INVx2_ASAP7_75t_L g4515 ( 
.A(n_4217),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4073),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_4084),
.Y(n_4517)
);

INVx3_ASAP7_75t_L g4518 ( 
.A(n_3983),
.Y(n_4518)
);

BUFx6f_ASAP7_75t_L g4519 ( 
.A(n_4003),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4084),
.Y(n_4520)
);

AND2x2_ASAP7_75t_L g4521 ( 
.A(n_4046),
.B(n_3840),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_4104),
.B(n_3869),
.Y(n_4522)
);

BUFx12f_ASAP7_75t_L g4523 ( 
.A(n_4259),
.Y(n_4523)
);

OAI21x1_ASAP7_75t_L g4524 ( 
.A1(n_3904),
.A2(n_3714),
.B(n_3745),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_4091),
.Y(n_4525)
);

INVx2_ASAP7_75t_L g4526 ( 
.A(n_4217),
.Y(n_4526)
);

OAI21x1_ASAP7_75t_L g4527 ( 
.A1(n_3904),
.A2(n_3712),
.B(n_3708),
.Y(n_4527)
);

AND2x2_ASAP7_75t_L g4528 ( 
.A(n_4046),
.B(n_3840),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4091),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4093),
.Y(n_4530)
);

INVx3_ASAP7_75t_L g4531 ( 
.A(n_3983),
.Y(n_4531)
);

AOI21xp5_ASAP7_75t_L g4532 ( 
.A1(n_3915),
.A2(n_3614),
.B(n_3878),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_4093),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4099),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4099),
.Y(n_4535)
);

AO21x1_ASAP7_75t_SL g4536 ( 
.A1(n_4061),
.A2(n_3849),
.B(n_3671),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4101),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4101),
.Y(n_4538)
);

NOR2xp33_ASAP7_75t_L g4539 ( 
.A(n_4175),
.B(n_3550),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4114),
.Y(n_4540)
);

CKINVDCx20_ASAP7_75t_R g4541 ( 
.A(n_4038),
.Y(n_4541)
);

AO21x2_ASAP7_75t_L g4542 ( 
.A1(n_3960),
.A2(n_3733),
.B(n_3575),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4114),
.Y(n_4543)
);

BUFx2_ASAP7_75t_L g4544 ( 
.A(n_3899),
.Y(n_4544)
);

INVx2_ASAP7_75t_L g4545 ( 
.A(n_3919),
.Y(n_4545)
);

AOI22xp33_ASAP7_75t_L g4546 ( 
.A1(n_3990),
.A2(n_3692),
.B1(n_3531),
.B2(n_3637),
.Y(n_4546)
);

OAI21x1_ASAP7_75t_L g4547 ( 
.A1(n_4150),
.A2(n_4254),
.B(n_4092),
.Y(n_4547)
);

BUFx8_ASAP7_75t_L g4548 ( 
.A(n_4009),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4116),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_3919),
.Y(n_4550)
);

AOI22xp33_ASAP7_75t_L g4551 ( 
.A1(n_4317),
.A2(n_3692),
.B1(n_3637),
.B2(n_3619),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4116),
.Y(n_4552)
);

INVx2_ASAP7_75t_L g4553 ( 
.A(n_3941),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4090),
.B(n_3561),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4120),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_3974),
.Y(n_4556)
);

INVx2_ASAP7_75t_L g4557 ( 
.A(n_3974),
.Y(n_4557)
);

BUFx6f_ASAP7_75t_L g4558 ( 
.A(n_4003),
.Y(n_4558)
);

INVx2_ASAP7_75t_L g4559 ( 
.A(n_3974),
.Y(n_4559)
);

AND2x2_ASAP7_75t_L g4560 ( 
.A(n_4090),
.B(n_3561),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_4120),
.Y(n_4561)
);

OAI21x1_ASAP7_75t_L g4562 ( 
.A1(n_4254),
.A2(n_3712),
.B(n_3708),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4122),
.Y(n_4563)
);

INVx3_ASAP7_75t_L g4564 ( 
.A(n_3924),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4122),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_3975),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_3975),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_3975),
.Y(n_4568)
);

HB1xp67_ASAP7_75t_L g4569 ( 
.A(n_4284),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4126),
.Y(n_4570)
);

INVx2_ASAP7_75t_SL g4571 ( 
.A(n_3966),
.Y(n_4571)
);

HB1xp67_ASAP7_75t_L g4572 ( 
.A(n_4110),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_L g4573 ( 
.A(n_4136),
.B(n_3885),
.Y(n_4573)
);

OR2x6_ASAP7_75t_L g4574 ( 
.A(n_4389),
.B(n_3669),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4126),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_3941),
.Y(n_4576)
);

OAI21x1_ASAP7_75t_L g4577 ( 
.A1(n_4070),
.A2(n_3793),
.B(n_3790),
.Y(n_4577)
);

BUFx2_ASAP7_75t_L g4578 ( 
.A(n_3899),
.Y(n_4578)
);

BUFx3_ASAP7_75t_L g4579 ( 
.A(n_4103),
.Y(n_4579)
);

INVx1_ASAP7_75t_SL g4580 ( 
.A(n_4100),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4128),
.Y(n_4581)
);

INVx3_ASAP7_75t_L g4582 ( 
.A(n_3924),
.Y(n_4582)
);

INVx2_ASAP7_75t_L g4583 ( 
.A(n_3978),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4128),
.Y(n_4584)
);

OAI21x1_ASAP7_75t_L g4585 ( 
.A1(n_4070),
.A2(n_3793),
.B(n_3790),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4129),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4129),
.Y(n_4587)
);

BUFx2_ASAP7_75t_L g4588 ( 
.A(n_3981),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_3978),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4137),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4137),
.Y(n_4591)
);

OAI21xp5_ASAP7_75t_L g4592 ( 
.A1(n_4108),
.A2(n_3613),
.B(n_3844),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4147),
.B(n_3885),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4139),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4139),
.Y(n_4595)
);

AND2x2_ASAP7_75t_L g4596 ( 
.A(n_4118),
.B(n_3564),
.Y(n_4596)
);

INVx1_ASAP7_75t_SL g4597 ( 
.A(n_3986),
.Y(n_4597)
);

HB1xp67_ASAP7_75t_SL g4598 ( 
.A(n_4103),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_4148),
.B(n_3640),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_3978),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_3993),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4118),
.B(n_3564),
.Y(n_4602)
);

INVx3_ASAP7_75t_L g4603 ( 
.A(n_3924),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4171),
.B(n_3573),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_3993),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4140),
.Y(n_4606)
);

INVx2_ASAP7_75t_L g4607 ( 
.A(n_3993),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4140),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4143),
.Y(n_4609)
);

BUFx2_ASAP7_75t_L g4610 ( 
.A(n_3981),
.Y(n_4610)
);

AND2x4_ASAP7_75t_L g4611 ( 
.A(n_3907),
.B(n_3619),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4143),
.Y(n_4612)
);

BUFx6f_ASAP7_75t_L g4613 ( 
.A(n_4003),
.Y(n_4613)
);

BUFx2_ASAP7_75t_L g4614 ( 
.A(n_3966),
.Y(n_4614)
);

BUFx2_ASAP7_75t_L g4615 ( 
.A(n_3966),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_3995),
.Y(n_4616)
);

INVxp67_ASAP7_75t_L g4617 ( 
.A(n_4159),
.Y(n_4617)
);

BUFx2_ASAP7_75t_L g4618 ( 
.A(n_4112),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_3995),
.Y(n_4619)
);

OAI21x1_ASAP7_75t_L g4620 ( 
.A1(n_4092),
.A2(n_3797),
.B(n_3794),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4149),
.Y(n_4621)
);

CKINVDCx20_ASAP7_75t_R g4622 ( 
.A(n_3951),
.Y(n_4622)
);

HB1xp67_ASAP7_75t_SL g4623 ( 
.A(n_4103),
.Y(n_4623)
);

INVx3_ASAP7_75t_L g4624 ( 
.A(n_3924),
.Y(n_4624)
);

INVx2_ASAP7_75t_L g4625 ( 
.A(n_3995),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4149),
.Y(n_4626)
);

AND2x2_ASAP7_75t_L g4627 ( 
.A(n_4171),
.B(n_3573),
.Y(n_4627)
);

CKINVDCx5p33_ASAP7_75t_R g4628 ( 
.A(n_3979),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_4155),
.B(n_4163),
.Y(n_4629)
);

INVx2_ASAP7_75t_L g4630 ( 
.A(n_3902),
.Y(n_4630)
);

INVx3_ASAP7_75t_L g4631 ( 
.A(n_3969),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4151),
.Y(n_4632)
);

HB1xp67_ASAP7_75t_L g4633 ( 
.A(n_4184),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4151),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4152),
.Y(n_4635)
);

INVx3_ASAP7_75t_L g4636 ( 
.A(n_3969),
.Y(n_4636)
);

HB1xp67_ASAP7_75t_L g4637 ( 
.A(n_4196),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4152),
.Y(n_4638)
);

NAND2x1p5_ASAP7_75t_L g4639 ( 
.A(n_3907),
.B(n_3856),
.Y(n_4639)
);

INVxp67_ASAP7_75t_SL g4640 ( 
.A(n_4121),
.Y(n_4640)
);

BUFx2_ASAP7_75t_L g4641 ( 
.A(n_4112),
.Y(n_4641)
);

NOR2x1_ASAP7_75t_SL g4642 ( 
.A(n_4377),
.B(n_4125),
.Y(n_4642)
);

INVx2_ASAP7_75t_SL g4643 ( 
.A(n_4042),
.Y(n_4643)
);

BUFx3_ASAP7_75t_L g4644 ( 
.A(n_4103),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_3902),
.Y(n_4645)
);

BUFx6f_ASAP7_75t_L g4646 ( 
.A(n_4333),
.Y(n_4646)
);

INVx2_ASAP7_75t_L g4647 ( 
.A(n_3902),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4153),
.Y(n_4648)
);

BUFx3_ASAP7_75t_L g4649 ( 
.A(n_4105),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4153),
.Y(n_4650)
);

BUFx3_ASAP7_75t_L g4651 ( 
.A(n_4105),
.Y(n_4651)
);

INVx2_ASAP7_75t_L g4652 ( 
.A(n_3914),
.Y(n_4652)
);

INVx2_ASAP7_75t_L g4653 ( 
.A(n_3914),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_SL g4654 ( 
.A(n_4121),
.B(n_3718),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_3914),
.Y(n_4655)
);

INVx2_ASAP7_75t_L g4656 ( 
.A(n_3921),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4154),
.Y(n_4657)
);

INVx2_ASAP7_75t_L g4658 ( 
.A(n_3921),
.Y(n_4658)
);

INVx3_ASAP7_75t_L g4659 ( 
.A(n_3969),
.Y(n_4659)
);

NAND2xp5_ASAP7_75t_L g4660 ( 
.A(n_4229),
.B(n_3600),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4154),
.Y(n_4661)
);

INVx2_ASAP7_75t_L g4662 ( 
.A(n_3921),
.Y(n_4662)
);

INVx2_ASAP7_75t_L g4663 ( 
.A(n_3923),
.Y(n_4663)
);

BUFx2_ASAP7_75t_L g4664 ( 
.A(n_4112),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_4232),
.B(n_3600),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4161),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_3923),
.Y(n_4667)
);

AOI22xp33_ASAP7_75t_L g4668 ( 
.A1(n_4289),
.A2(n_3637),
.B1(n_3619),
.B2(n_3880),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_3923),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4161),
.Y(n_4670)
);

OAI21x1_ASAP7_75t_L g4671 ( 
.A1(n_4010),
.A2(n_3797),
.B(n_3794),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4076),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4167),
.Y(n_4673)
);

HB1xp67_ASAP7_75t_L g4674 ( 
.A(n_4297),
.Y(n_4674)
);

INVx3_ASAP7_75t_L g4675 ( 
.A(n_3969),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4167),
.Y(n_4676)
);

BUFx3_ASAP7_75t_L g4677 ( 
.A(n_4105),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4180),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4195),
.B(n_4257),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4180),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4190),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4190),
.Y(n_4682)
);

NOR2xp33_ASAP7_75t_L g4683 ( 
.A(n_3955),
.B(n_3665),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4191),
.Y(n_4684)
);

BUFx2_ASAP7_75t_L g4685 ( 
.A(n_4169),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4191),
.Y(n_4686)
);

BUFx2_ASAP7_75t_SL g4687 ( 
.A(n_4169),
.Y(n_4687)
);

HB1xp67_ASAP7_75t_L g4688 ( 
.A(n_4337),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4192),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4192),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4199),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_L g4692 ( 
.A(n_4315),
.B(n_3744),
.Y(n_4692)
);

INVx2_ASAP7_75t_L g4693 ( 
.A(n_3999),
.Y(n_4693)
);

NAND2x1p5_ASAP7_75t_L g4694 ( 
.A(n_3907),
.B(n_3856),
.Y(n_4694)
);

AND2x2_ASAP7_75t_L g4695 ( 
.A(n_4195),
.B(n_3583),
.Y(n_4695)
);

INVx3_ASAP7_75t_L g4696 ( 
.A(n_3994),
.Y(n_4696)
);

INVxp33_ASAP7_75t_L g4697 ( 
.A(n_4022),
.Y(n_4697)
);

NOR2xp33_ASAP7_75t_L g4698 ( 
.A(n_3955),
.B(n_3678),
.Y(n_4698)
);

INVx4_ASAP7_75t_L g4699 ( 
.A(n_3982),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4199),
.Y(n_4700)
);

AOI22xp5_ASAP7_75t_L g4701 ( 
.A1(n_4381),
.A2(n_3667),
.B1(n_3608),
.B2(n_3635),
.Y(n_4701)
);

INVx2_ASAP7_75t_L g4702 ( 
.A(n_3999),
.Y(n_4702)
);

OAI21xp5_ASAP7_75t_L g4703 ( 
.A1(n_4130),
.A2(n_3844),
.B(n_3839),
.Y(n_4703)
);

AND2x4_ASAP7_75t_L g4704 ( 
.A(n_3907),
.B(n_3619),
.Y(n_4704)
);

OAI21x1_ASAP7_75t_L g4705 ( 
.A1(n_4010),
.A2(n_3807),
.B(n_3800),
.Y(n_4705)
);

INVx3_ASAP7_75t_L g4706 ( 
.A(n_3994),
.Y(n_4706)
);

OAI21x1_ASAP7_75t_L g4707 ( 
.A1(n_4027),
.A2(n_4058),
.B(n_4350),
.Y(n_4707)
);

NOR2xp33_ASAP7_75t_SL g4708 ( 
.A(n_4275),
.B(n_3534),
.Y(n_4708)
);

CKINVDCx16_ASAP7_75t_R g4709 ( 
.A(n_4009),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4201),
.Y(n_4710)
);

OR2x2_ASAP7_75t_L g4711 ( 
.A(n_4235),
.B(n_3861),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4201),
.Y(n_4712)
);

BUFx3_ASAP7_75t_L g4713 ( 
.A(n_4105),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4257),
.B(n_3583),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4204),
.Y(n_4715)
);

AND2x2_ASAP7_75t_L g4716 ( 
.A(n_4277),
.B(n_3547),
.Y(n_4716)
);

OAI21x1_ASAP7_75t_L g4717 ( 
.A1(n_4027),
.A2(n_3807),
.B(n_3800),
.Y(n_4717)
);

OR2x2_ASAP7_75t_L g4718 ( 
.A(n_3954),
.B(n_3761),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4204),
.Y(n_4719)
);

AO21x2_ASAP7_75t_L g4720 ( 
.A1(n_3963),
.A2(n_3575),
.B(n_3722),
.Y(n_4720)
);

HB1xp67_ASAP7_75t_L g4721 ( 
.A(n_4338),
.Y(n_4721)
);

INVx2_ASAP7_75t_L g4722 ( 
.A(n_3999),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_4205),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4205),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4206),
.Y(n_4725)
);

CKINVDCx11_ASAP7_75t_R g4726 ( 
.A(n_3955),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4206),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4145),
.B(n_4107),
.Y(n_4728)
);

OR2x2_ASAP7_75t_L g4729 ( 
.A(n_4216),
.B(n_3761),
.Y(n_4729)
);

AND2x4_ASAP7_75t_L g4730 ( 
.A(n_3907),
.B(n_3637),
.Y(n_4730)
);

OA21x2_ASAP7_75t_L g4731 ( 
.A1(n_3963),
.A2(n_3976),
.B(n_3967),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4208),
.Y(n_4732)
);

INVx2_ASAP7_75t_L g4733 ( 
.A(n_4000),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4208),
.Y(n_4734)
);

AND2x4_ASAP7_75t_L g4735 ( 
.A(n_3905),
.B(n_3896),
.Y(n_4735)
);

OA21x2_ASAP7_75t_L g4736 ( 
.A1(n_3967),
.A2(n_3755),
.B(n_3750),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4000),
.Y(n_4737)
);

HB1xp67_ASAP7_75t_L g4738 ( 
.A(n_4375),
.Y(n_4738)
);

AND2x2_ASAP7_75t_L g4739 ( 
.A(n_4277),
.B(n_3547),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4211),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4211),
.Y(n_4741)
);

INVx2_ASAP7_75t_L g4742 ( 
.A(n_4000),
.Y(n_4742)
);

NAND2x1p5_ASAP7_75t_L g4743 ( 
.A(n_4174),
.B(n_3856),
.Y(n_4743)
);

HB1xp67_ASAP7_75t_L g4744 ( 
.A(n_3938),
.Y(n_4744)
);

BUFx3_ASAP7_75t_L g4745 ( 
.A(n_4158),
.Y(n_4745)
);

INVx2_ASAP7_75t_L g4746 ( 
.A(n_4005),
.Y(n_4746)
);

INVx2_ASAP7_75t_L g4747 ( 
.A(n_4005),
.Y(n_4747)
);

INVx2_ASAP7_75t_L g4748 ( 
.A(n_4005),
.Y(n_4748)
);

OA21x2_ASAP7_75t_L g4749 ( 
.A1(n_3976),
.A2(n_3756),
.B(n_3755),
.Y(n_4749)
);

OAI21x1_ASAP7_75t_L g4750 ( 
.A1(n_4058),
.A2(n_3823),
.B(n_3816),
.Y(n_4750)
);

AOI22xp5_ASAP7_75t_L g4751 ( 
.A1(n_4409),
.A2(n_3608),
.B1(n_3626),
.B2(n_3669),
.Y(n_4751)
);

INVx2_ASAP7_75t_L g4752 ( 
.A(n_4019),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4220),
.Y(n_4753)
);

BUFx3_ASAP7_75t_L g4754 ( 
.A(n_4158),
.Y(n_4754)
);

NAND2x1_ASAP7_75t_L g4755 ( 
.A(n_4374),
.B(n_4408),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4220),
.Y(n_4756)
);

BUFx2_ASAP7_75t_L g4757 ( 
.A(n_4169),
.Y(n_4757)
);

OAI21xp5_ASAP7_75t_L g4758 ( 
.A1(n_3908),
.A2(n_3888),
.B(n_3849),
.Y(n_4758)
);

INVx2_ASAP7_75t_L g4759 ( 
.A(n_4019),
.Y(n_4759)
);

OR2x2_ASAP7_75t_L g4760 ( 
.A(n_4216),
.B(n_3791),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4223),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4359),
.B(n_3744),
.Y(n_4762)
);

OR2x6_ASAP7_75t_L g4763 ( 
.A(n_4389),
.B(n_4399),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4223),
.Y(n_4764)
);

INVx4_ASAP7_75t_L g4765 ( 
.A(n_3982),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4224),
.Y(n_4766)
);

INVx2_ASAP7_75t_L g4767 ( 
.A(n_4019),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4026),
.Y(n_4768)
);

INVx2_ASAP7_75t_L g4769 ( 
.A(n_4026),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4224),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4225),
.Y(n_4771)
);

AND2x2_ASAP7_75t_L g4772 ( 
.A(n_4359),
.B(n_3547),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4225),
.Y(n_4773)
);

INVx2_ASAP7_75t_L g4774 ( 
.A(n_4026),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4231),
.Y(n_4775)
);

OAI22xp5_ASAP7_75t_L g4776 ( 
.A1(n_3908),
.A2(n_3762),
.B1(n_3875),
.B2(n_3539),
.Y(n_4776)
);

AO21x2_ASAP7_75t_L g4777 ( 
.A1(n_3985),
.A2(n_3575),
.B(n_3700),
.Y(n_4777)
);

INVx2_ASAP7_75t_L g4778 ( 
.A(n_4076),
.Y(n_4778)
);

OAI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4141),
.A2(n_3612),
.B(n_3685),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4076),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4231),
.Y(n_4781)
);

INVx2_ASAP7_75t_L g4782 ( 
.A(n_4077),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4236),
.Y(n_4783)
);

NOR2xp33_ASAP7_75t_L g4784 ( 
.A(n_3906),
.B(n_3678),
.Y(n_4784)
);

HB1xp67_ASAP7_75t_L g4785 ( 
.A(n_3973),
.Y(n_4785)
);

INVx2_ASAP7_75t_L g4786 ( 
.A(n_4077),
.Y(n_4786)
);

BUFx2_ASAP7_75t_L g4787 ( 
.A(n_4290),
.Y(n_4787)
);

AND2x2_ASAP7_75t_L g4788 ( 
.A(n_4062),
.B(n_3547),
.Y(n_4788)
);

INVx2_ASAP7_75t_L g4789 ( 
.A(n_4077),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4236),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4243),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4243),
.Y(n_4792)
);

INVx2_ASAP7_75t_SL g4793 ( 
.A(n_4042),
.Y(n_4793)
);

INVx2_ASAP7_75t_L g4794 ( 
.A(n_4080),
.Y(n_4794)
);

BUFx3_ASAP7_75t_L g4795 ( 
.A(n_4168),
.Y(n_4795)
);

AOI22xp33_ASAP7_75t_SL g4796 ( 
.A1(n_4408),
.A2(n_3880),
.B1(n_3826),
.B2(n_3836),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4245),
.Y(n_4797)
);

INVx2_ASAP7_75t_L g4798 ( 
.A(n_4080),
.Y(n_4798)
);

OAI21x1_ASAP7_75t_L g4799 ( 
.A1(n_4350),
.A2(n_4386),
.B(n_4364),
.Y(n_4799)
);

INVx2_ASAP7_75t_L g4800 ( 
.A(n_4080),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4245),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_3920),
.B(n_3893),
.Y(n_4802)
);

AND2x2_ASAP7_75t_SL g4803 ( 
.A(n_4182),
.B(n_3556),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4081),
.Y(n_4804)
);

AOI22xp33_ASAP7_75t_SL g4805 ( 
.A1(n_4334),
.A2(n_3880),
.B1(n_3826),
.B2(n_3836),
.Y(n_4805)
);

OAI21x1_ASAP7_75t_L g4806 ( 
.A1(n_4364),
.A2(n_3823),
.B(n_3816),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4062),
.B(n_3883),
.Y(n_4807)
);

INVx2_ASAP7_75t_L g4808 ( 
.A(n_4081),
.Y(n_4808)
);

NAND3xp33_ASAP7_75t_L g4809 ( 
.A(n_4132),
.B(n_3784),
.C(n_3684),
.Y(n_4809)
);

OR2x2_ASAP7_75t_L g4810 ( 
.A(n_3973),
.B(n_4008),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4246),
.Y(n_4811)
);

AND2x4_ASAP7_75t_L g4812 ( 
.A(n_3905),
.B(n_3646),
.Y(n_4812)
);

CKINVDCx5p33_ASAP7_75t_R g4813 ( 
.A(n_4193),
.Y(n_4813)
);

AND2x2_ASAP7_75t_L g4814 ( 
.A(n_4085),
.B(n_3880),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4246),
.Y(n_4815)
);

INVx2_ASAP7_75t_L g4816 ( 
.A(n_4081),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4034),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4247),
.Y(n_4818)
);

INVxp33_ASAP7_75t_L g4819 ( 
.A(n_4373),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4247),
.Y(n_4820)
);

INVx2_ASAP7_75t_L g4821 ( 
.A(n_4034),
.Y(n_4821)
);

OR2x2_ASAP7_75t_L g4822 ( 
.A(n_4031),
.B(n_3791),
.Y(n_4822)
);

INVx2_ASAP7_75t_L g4823 ( 
.A(n_4035),
.Y(n_4823)
);

INVx2_ASAP7_75t_L g4824 ( 
.A(n_4035),
.Y(n_4824)
);

INVx2_ASAP7_75t_L g4825 ( 
.A(n_4047),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4250),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4250),
.Y(n_4827)
);

BUFx2_ASAP7_75t_L g4828 ( 
.A(n_4290),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4260),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4260),
.Y(n_4830)
);

AOI21x1_ASAP7_75t_L g4831 ( 
.A1(n_3930),
.A2(n_3826),
.B(n_3825),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4262),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4262),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4264),
.Y(n_4834)
);

OA21x2_ASAP7_75t_L g4835 ( 
.A1(n_3985),
.A2(n_3757),
.B(n_3756),
.Y(n_4835)
);

INVx2_ASAP7_75t_L g4836 ( 
.A(n_4047),
.Y(n_4836)
);

INVx1_ASAP7_75t_L g4837 ( 
.A(n_4264),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4265),
.Y(n_4838)
);

HB1xp67_ASAP7_75t_L g4839 ( 
.A(n_4031),
.Y(n_4839)
);

INVx2_ASAP7_75t_SL g4840 ( 
.A(n_4042),
.Y(n_4840)
);

HB1xp67_ASAP7_75t_L g4841 ( 
.A(n_4265),
.Y(n_4841)
);

BUFx2_ASAP7_75t_L g4842 ( 
.A(n_4362),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4270),
.Y(n_4843)
);

INVx3_ASAP7_75t_L g4844 ( 
.A(n_3994),
.Y(n_4844)
);

AO31x2_ASAP7_75t_L g4845 ( 
.A1(n_3989),
.A2(n_3624),
.A3(n_3627),
.B(n_3609),
.Y(n_4845)
);

INVx2_ASAP7_75t_SL g4846 ( 
.A(n_4202),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4270),
.Y(n_4847)
);

NOR2xp33_ASAP7_75t_L g4848 ( 
.A(n_4239),
.B(n_3678),
.Y(n_4848)
);

INVx2_ASAP7_75t_L g4849 ( 
.A(n_4049),
.Y(n_4849)
);

HB1xp67_ASAP7_75t_L g4850 ( 
.A(n_4271),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4271),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4272),
.Y(n_4852)
);

OAI22xp5_ASAP7_75t_L g4853 ( 
.A1(n_4314),
.A2(n_3539),
.B1(n_3879),
.B2(n_3606),
.Y(n_4853)
);

INVx2_ASAP7_75t_L g4854 ( 
.A(n_4049),
.Y(n_4854)
);

BUFx6f_ASAP7_75t_L g4855 ( 
.A(n_4333),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4085),
.B(n_3606),
.Y(n_4856)
);

HB1xp67_ASAP7_75t_L g4857 ( 
.A(n_4272),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4273),
.Y(n_4858)
);

AND2x2_ASAP7_75t_L g4859 ( 
.A(n_4251),
.B(n_3606),
.Y(n_4859)
);

INVx2_ASAP7_75t_L g4860 ( 
.A(n_3994),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4251),
.B(n_3606),
.Y(n_4861)
);

AOI22xp33_ASAP7_75t_L g4862 ( 
.A1(n_4060),
.A2(n_3594),
.B1(n_3656),
.B2(n_3806),
.Y(n_4862)
);

INVx2_ASAP7_75t_L g4863 ( 
.A(n_4024),
.Y(n_4863)
);

OA21x2_ASAP7_75t_L g4864 ( 
.A1(n_3989),
.A2(n_3757),
.B(n_3584),
.Y(n_4864)
);

INVx2_ASAP7_75t_L g4865 ( 
.A(n_4024),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4273),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4274),
.Y(n_4867)
);

HB1xp67_ASAP7_75t_L g4868 ( 
.A(n_4274),
.Y(n_4868)
);

INVx2_ASAP7_75t_L g4869 ( 
.A(n_4094),
.Y(n_4869)
);

INVx3_ASAP7_75t_L g4870 ( 
.A(n_4024),
.Y(n_4870)
);

INVx2_ASAP7_75t_L g4871 ( 
.A(n_4094),
.Y(n_4871)
);

OAI21x1_ASAP7_75t_L g4872 ( 
.A1(n_4386),
.A2(n_3841),
.B(n_3824),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4276),
.Y(n_4873)
);

AND2x4_ASAP7_75t_L g4874 ( 
.A(n_3905),
.B(n_3646),
.Y(n_4874)
);

HB1xp67_ASAP7_75t_L g4875 ( 
.A(n_4276),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_L g4876 ( 
.A(n_3920),
.B(n_3893),
.Y(n_4876)
);

INVxp33_ASAP7_75t_L g4877 ( 
.A(n_4064),
.Y(n_4877)
);

OR2x2_ASAP7_75t_L g4878 ( 
.A(n_4156),
.B(n_3846),
.Y(n_4878)
);

INVx3_ASAP7_75t_L g4879 ( 
.A(n_4024),
.Y(n_4879)
);

INVx2_ASAP7_75t_L g4880 ( 
.A(n_4094),
.Y(n_4880)
);

HB1xp67_ASAP7_75t_L g4881 ( 
.A(n_4278),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4278),
.Y(n_4882)
);

INVx2_ASAP7_75t_L g4883 ( 
.A(n_4032),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4283),
.Y(n_4884)
);

AOI22xp33_ASAP7_75t_L g4885 ( 
.A1(n_3901),
.A2(n_3594),
.B1(n_3656),
.B2(n_3608),
.Y(n_4885)
);

HB1xp67_ASAP7_75t_L g4886 ( 
.A(n_4283),
.Y(n_4886)
);

AOI22xp33_ASAP7_75t_L g4887 ( 
.A1(n_3948),
.A2(n_3594),
.B1(n_3656),
.B2(n_3608),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4286),
.Y(n_4888)
);

INVx2_ASAP7_75t_L g4889 ( 
.A(n_4098),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4286),
.Y(n_4890)
);

INVxp67_ASAP7_75t_L g4891 ( 
.A(n_4125),
.Y(n_4891)
);

INVx2_ASAP7_75t_L g4892 ( 
.A(n_4098),
.Y(n_4892)
);

INVx2_ASAP7_75t_L g4893 ( 
.A(n_4098),
.Y(n_4893)
);

HB1xp67_ASAP7_75t_L g4894 ( 
.A(n_4292),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_4252),
.B(n_3646),
.Y(n_4895)
);

INVx2_ASAP7_75t_L g4896 ( 
.A(n_4106),
.Y(n_4896)
);

INVx2_ASAP7_75t_L g4897 ( 
.A(n_4106),
.Y(n_4897)
);

OAI21xp5_ASAP7_75t_L g4898 ( 
.A1(n_4390),
.A2(n_3539),
.B(n_3818),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4292),
.Y(n_4899)
);

OAI21x1_ASAP7_75t_L g4900 ( 
.A1(n_4348),
.A2(n_3841),
.B(n_3824),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4293),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4293),
.Y(n_4902)
);

OAI22xp33_ASAP7_75t_L g4903 ( 
.A1(n_4183),
.A2(n_3656),
.B1(n_3856),
.B2(n_3743),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4294),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4294),
.Y(n_4905)
);

INVx2_ASAP7_75t_L g4906 ( 
.A(n_4106),
.Y(n_4906)
);

OR2x2_ASAP7_75t_L g4907 ( 
.A(n_4156),
.B(n_3846),
.Y(n_4907)
);

NAND2x1p5_ASAP7_75t_L g4908 ( 
.A(n_4174),
.B(n_3856),
.Y(n_4908)
);

INVx1_ASAP7_75t_L g4909 ( 
.A(n_4299),
.Y(n_4909)
);

INVx3_ASAP7_75t_L g4910 ( 
.A(n_4032),
.Y(n_4910)
);

OAI21x1_ASAP7_75t_L g4911 ( 
.A1(n_4348),
.A2(n_3851),
.B(n_3842),
.Y(n_4911)
);

HB1xp67_ASAP7_75t_L g4912 ( 
.A(n_4299),
.Y(n_4912)
);

INVx2_ASAP7_75t_L g4913 ( 
.A(n_4032),
.Y(n_4913)
);

BUFx6f_ASAP7_75t_L g4914 ( 
.A(n_4333),
.Y(n_4914)
);

BUFx6f_ASAP7_75t_L g4915 ( 
.A(n_4333),
.Y(n_4915)
);

O2A1O1Ixp33_ASAP7_75t_L g4916 ( 
.A1(n_4323),
.A2(n_3832),
.B(n_3822),
.C(n_3509),
.Y(n_4916)
);

INVx1_ASAP7_75t_SL g4917 ( 
.A(n_4016),
.Y(n_4917)
);

AND2x2_ASAP7_75t_L g4918 ( 
.A(n_4252),
.B(n_3646),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4300),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4300),
.Y(n_4920)
);

INVxp33_ASAP7_75t_L g4921 ( 
.A(n_3957),
.Y(n_4921)
);

BUFx2_ASAP7_75t_L g4922 ( 
.A(n_4362),
.Y(n_4922)
);

INVx2_ASAP7_75t_L g4923 ( 
.A(n_4032),
.Y(n_4923)
);

AO21x2_ASAP7_75t_L g4924 ( 
.A1(n_3930),
.A2(n_3575),
.B(n_3697),
.Y(n_4924)
);

INVx2_ASAP7_75t_L g4925 ( 
.A(n_4065),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4304),
.Y(n_4926)
);

BUFx3_ASAP7_75t_L g4927 ( 
.A(n_4514),
.Y(n_4927)
);

INVx2_ASAP7_75t_L g4928 ( 
.A(n_4731),
.Y(n_4928)
);

INVx2_ASAP7_75t_L g4929 ( 
.A(n_4731),
.Y(n_4929)
);

AND2x2_ASAP7_75t_L g4930 ( 
.A(n_4432),
.B(n_4642),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4841),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_4850),
.Y(n_4932)
);

AND2x2_ASAP7_75t_L g4933 ( 
.A(n_4432),
.B(n_4642),
.Y(n_4933)
);

INVx2_ASAP7_75t_L g4934 ( 
.A(n_4731),
.Y(n_4934)
);

HB1xp67_ASAP7_75t_L g4935 ( 
.A(n_4674),
.Y(n_4935)
);

AND2x4_ASAP7_75t_L g4936 ( 
.A(n_4614),
.B(n_3905),
.Y(n_4936)
);

OA21x2_ASAP7_75t_L g4937 ( 
.A1(n_4484),
.A2(n_3939),
.B(n_3930),
.Y(n_4937)
);

AO21x2_ASAP7_75t_L g4938 ( 
.A1(n_4640),
.A2(n_4707),
.B(n_4779),
.Y(n_4938)
);

OA21x2_ASAP7_75t_L g4939 ( 
.A1(n_4484),
.A2(n_3940),
.B(n_3939),
.Y(n_4939)
);

OR2x2_ASAP7_75t_L g4940 ( 
.A(n_4760),
.B(n_4288),
.Y(n_4940)
);

AO21x2_ASAP7_75t_L g4941 ( 
.A1(n_4707),
.A2(n_3940),
.B(n_3939),
.Y(n_4941)
);

INVx4_ASAP7_75t_SL g4942 ( 
.A(n_4514),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_4857),
.Y(n_4943)
);

OAI21xp5_ASAP7_75t_L g4944 ( 
.A1(n_4446),
.A2(n_3965),
.B(n_4309),
.Y(n_4944)
);

OR2x2_ASAP7_75t_L g4945 ( 
.A(n_4760),
.B(n_4288),
.Y(n_4945)
);

OR2x2_ASAP7_75t_L g4946 ( 
.A(n_4472),
.B(n_4302),
.Y(n_4946)
);

INVx2_ASAP7_75t_L g4947 ( 
.A(n_4731),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4868),
.Y(n_4948)
);

INVx2_ASAP7_75t_L g4949 ( 
.A(n_4924),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4875),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4881),
.Y(n_4951)
);

INVx3_ASAP7_75t_L g4952 ( 
.A(n_4417),
.Y(n_4952)
);

INVx2_ASAP7_75t_L g4953 ( 
.A(n_4924),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_L g4954 ( 
.A(n_4465),
.B(n_4471),
.Y(n_4954)
);

AND2x2_ASAP7_75t_L g4955 ( 
.A(n_4614),
.B(n_4328),
.Y(n_4955)
);

CKINVDCx5p33_ASAP7_75t_R g4956 ( 
.A(n_4726),
.Y(n_4956)
);

INVx2_ASAP7_75t_L g4957 ( 
.A(n_4924),
.Y(n_4957)
);

INVx2_ASAP7_75t_L g4958 ( 
.A(n_4736),
.Y(n_4958)
);

AO21x2_ASAP7_75t_L g4959 ( 
.A1(n_4809),
.A2(n_3943),
.B(n_3940),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4886),
.Y(n_4960)
);

OR2x2_ASAP7_75t_L g4961 ( 
.A(n_4472),
.B(n_4302),
.Y(n_4961)
);

INVx2_ASAP7_75t_L g4962 ( 
.A(n_4736),
.Y(n_4962)
);

BUFx2_ASAP7_75t_L g4963 ( 
.A(n_4579),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4894),
.Y(n_4964)
);

BUFx6f_ASAP7_75t_L g4965 ( 
.A(n_4424),
.Y(n_4965)
);

AND2x2_ASAP7_75t_L g4966 ( 
.A(n_4615),
.B(n_4328),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4912),
.Y(n_4967)
);

INVx3_ASAP7_75t_L g4968 ( 
.A(n_4417),
.Y(n_4968)
);

AO21x2_ASAP7_75t_L g4969 ( 
.A1(n_4777),
.A2(n_3943),
.B(n_3909),
.Y(n_4969)
);

INVx3_ASAP7_75t_L g4970 ( 
.A(n_4417),
.Y(n_4970)
);

AND2x2_ASAP7_75t_L g4971 ( 
.A(n_4615),
.B(n_3972),
.Y(n_4971)
);

OR2x2_ASAP7_75t_L g4972 ( 
.A(n_4822),
.B(n_3903),
.Y(n_4972)
);

AND2x2_ASAP7_75t_L g4973 ( 
.A(n_4803),
.B(n_3972),
.Y(n_4973)
);

AND2x2_ASAP7_75t_L g4974 ( 
.A(n_4803),
.B(n_4298),
.Y(n_4974)
);

AND2x2_ASAP7_75t_L g4975 ( 
.A(n_4803),
.B(n_4298),
.Y(n_4975)
);

HB1xp67_ASAP7_75t_L g4976 ( 
.A(n_4688),
.Y(n_4976)
);

INVx2_ASAP7_75t_L g4977 ( 
.A(n_4736),
.Y(n_4977)
);

AND2x2_ASAP7_75t_L g4978 ( 
.A(n_4685),
.B(n_4351),
.Y(n_4978)
);

AND2x2_ASAP7_75t_L g4979 ( 
.A(n_4685),
.B(n_4351),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4416),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4416),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4418),
.Y(n_4982)
);

OR2x2_ASAP7_75t_L g4983 ( 
.A(n_4822),
.B(n_3903),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_4418),
.Y(n_4984)
);

AND2x2_ASAP7_75t_L g4985 ( 
.A(n_4757),
.B(n_4735),
.Y(n_4985)
);

INVx3_ASAP7_75t_L g4986 ( 
.A(n_4417),
.Y(n_4986)
);

INVx2_ASAP7_75t_SL g4987 ( 
.A(n_4579),
.Y(n_4987)
);

BUFx2_ASAP7_75t_L g4988 ( 
.A(n_4579),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_SL g4989 ( 
.A(n_4532),
.B(n_4314),
.Y(n_4989)
);

HB1xp67_ASAP7_75t_L g4990 ( 
.A(n_4721),
.Y(n_4990)
);

HB1xp67_ASAP7_75t_L g4991 ( 
.A(n_4738),
.Y(n_4991)
);

INVx2_ASAP7_75t_L g4992 ( 
.A(n_4736),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4421),
.Y(n_4993)
);

BUFx10_ASAP7_75t_L g4994 ( 
.A(n_4539),
.Y(n_4994)
);

OR2x6_ASAP7_75t_L g4995 ( 
.A(n_4639),
.B(n_4414),
.Y(n_4995)
);

AND2x2_ASAP7_75t_L g4996 ( 
.A(n_4757),
.B(n_4198),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4421),
.Y(n_4997)
);

INVx3_ASAP7_75t_L g4998 ( 
.A(n_4437),
.Y(n_4998)
);

INVx2_ASAP7_75t_SL g4999 ( 
.A(n_4644),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4422),
.Y(n_5000)
);

INVx2_ASAP7_75t_L g5001 ( 
.A(n_4749),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4422),
.Y(n_5002)
);

INVx3_ASAP7_75t_L g5003 ( 
.A(n_4437),
.Y(n_5003)
);

HB1xp67_ASAP7_75t_L g5004 ( 
.A(n_4507),
.Y(n_5004)
);

BUFx3_ASAP7_75t_L g5005 ( 
.A(n_4424),
.Y(n_5005)
);

HB1xp67_ASAP7_75t_L g5006 ( 
.A(n_4447),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_4735),
.B(n_4198),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4423),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4423),
.Y(n_5009)
);

INVx2_ASAP7_75t_L g5010 ( 
.A(n_4749),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4425),
.Y(n_5011)
);

OAI21x1_ASAP7_75t_L g5012 ( 
.A1(n_4437),
.A2(n_3934),
.B(n_3912),
.Y(n_5012)
);

INVx2_ASAP7_75t_L g5013 ( 
.A(n_4749),
.Y(n_5013)
);

AO21x2_ASAP7_75t_L g5014 ( 
.A1(n_4777),
.A2(n_3943),
.B(n_3910),
.Y(n_5014)
);

OR2x6_ASAP7_75t_L g5015 ( 
.A(n_4639),
.B(n_4414),
.Y(n_5015)
);

HB1xp67_ASAP7_75t_L g5016 ( 
.A(n_4452),
.Y(n_5016)
);

OA21x2_ASAP7_75t_L g5017 ( 
.A1(n_4430),
.A2(n_3910),
.B(n_3909),
.Y(n_5017)
);

AOI21x1_ASAP7_75t_L g5018 ( 
.A1(n_4787),
.A2(n_4374),
.B(n_3913),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4425),
.Y(n_5019)
);

OA21x2_ASAP7_75t_L g5020 ( 
.A1(n_4430),
.A2(n_3913),
.B(n_3911),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_4428),
.Y(n_5021)
);

INVx2_ASAP7_75t_L g5022 ( 
.A(n_4749),
.Y(n_5022)
);

AND2x2_ASAP7_75t_L g5023 ( 
.A(n_4735),
.B(n_4198),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4428),
.Y(n_5024)
);

INVx2_ASAP7_75t_L g5025 ( 
.A(n_4835),
.Y(n_5025)
);

NAND2xp5_ASAP7_75t_L g5026 ( 
.A(n_4504),
.B(n_4456),
.Y(n_5026)
);

OR2x2_ASAP7_75t_L g5027 ( 
.A(n_4718),
.B(n_3911),
.Y(n_5027)
);

INVx2_ASAP7_75t_L g5028 ( 
.A(n_4835),
.Y(n_5028)
);

INVx2_ASAP7_75t_L g5029 ( 
.A(n_4835),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4438),
.Y(n_5030)
);

INVx2_ASAP7_75t_L g5031 ( 
.A(n_4835),
.Y(n_5031)
);

INVx2_ASAP7_75t_L g5032 ( 
.A(n_4864),
.Y(n_5032)
);

OAI21xp5_ASAP7_75t_L g5033 ( 
.A1(n_4654),
.A2(n_4244),
.B(n_4056),
.Y(n_5033)
);

OR2x6_ASAP7_75t_L g5034 ( 
.A(n_4639),
.B(n_4389),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4438),
.Y(n_5035)
);

OR2x2_ASAP7_75t_L g5036 ( 
.A(n_4718),
.B(n_4599),
.Y(n_5036)
);

AND2x2_ASAP7_75t_L g5037 ( 
.A(n_4735),
.B(n_4198),
.Y(n_5037)
);

INVx2_ASAP7_75t_SL g5038 ( 
.A(n_4644),
.Y(n_5038)
);

AND2x2_ASAP7_75t_L g5039 ( 
.A(n_4772),
.B(n_4214),
.Y(n_5039)
);

INVx1_ASAP7_75t_L g5040 ( 
.A(n_4439),
.Y(n_5040)
);

INVx2_ASAP7_75t_L g5041 ( 
.A(n_4864),
.Y(n_5041)
);

AOI22xp33_ASAP7_75t_L g5042 ( 
.A1(n_4453),
.A2(n_4316),
.B1(n_4233),
.B2(n_4347),
.Y(n_5042)
);

INVxp33_ASAP7_75t_L g5043 ( 
.A(n_4708),
.Y(n_5043)
);

AND2x2_ASAP7_75t_L g5044 ( 
.A(n_4772),
.B(n_4214),
.Y(n_5044)
);

INVx2_ASAP7_75t_SL g5045 ( 
.A(n_4644),
.Y(n_5045)
);

OAI21xp5_ASAP7_75t_L g5046 ( 
.A1(n_4592),
.A2(n_4396),
.B(n_4325),
.Y(n_5046)
);

INVxp67_ASAP7_75t_L g5047 ( 
.A(n_4687),
.Y(n_5047)
);

INVx3_ASAP7_75t_L g5048 ( 
.A(n_4437),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_L g5049 ( 
.A(n_4728),
.B(n_4367),
.Y(n_5049)
);

AO21x2_ASAP7_75t_L g5050 ( 
.A1(n_4777),
.A2(n_3928),
.B(n_3931),
.Y(n_5050)
);

AND2x2_ASAP7_75t_L g5051 ( 
.A(n_4480),
.B(n_4214),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_4439),
.Y(n_5052)
);

OR2x2_ASAP7_75t_L g5053 ( 
.A(n_4729),
.B(n_3928),
.Y(n_5053)
);

INVx2_ASAP7_75t_L g5054 ( 
.A(n_4864),
.Y(n_5054)
);

INVx2_ASAP7_75t_L g5055 ( 
.A(n_4864),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4445),
.Y(n_5056)
);

BUFx2_ASAP7_75t_L g5057 ( 
.A(n_4649),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4445),
.Y(n_5058)
);

AND2x2_ASAP7_75t_L g5059 ( 
.A(n_4480),
.B(n_4214),
.Y(n_5059)
);

INVx2_ASAP7_75t_L g5060 ( 
.A(n_4556),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4451),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_4451),
.Y(n_5062)
);

OA21x2_ASAP7_75t_L g5063 ( 
.A1(n_4717),
.A2(n_3931),
.B(n_3929),
.Y(n_5063)
);

AO21x2_ASAP7_75t_L g5064 ( 
.A1(n_4542),
.A2(n_3935),
.B(n_3929),
.Y(n_5064)
);

OR2x2_ASAP7_75t_L g5065 ( 
.A(n_4729),
.B(n_4304),
.Y(n_5065)
);

OR2x2_ASAP7_75t_L g5066 ( 
.A(n_4711),
.B(n_4512),
.Y(n_5066)
);

INVx2_ASAP7_75t_SL g5067 ( 
.A(n_4649),
.Y(n_5067)
);

OA21x2_ASAP7_75t_L g5068 ( 
.A1(n_4717),
.A2(n_4705),
.B(n_4671),
.Y(n_5068)
);

INVx2_ASAP7_75t_L g5069 ( 
.A(n_4556),
.Y(n_5069)
);

OA21x2_ASAP7_75t_L g5070 ( 
.A1(n_4671),
.A2(n_3946),
.B(n_3935),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_4454),
.Y(n_5071)
);

NOR3xp33_ASAP7_75t_L g5072 ( 
.A(n_4699),
.B(n_4001),
.C(n_3982),
.Y(n_5072)
);

OR2x2_ASAP7_75t_L g5073 ( 
.A(n_4711),
.B(n_4305),
.Y(n_5073)
);

AND2x2_ASAP7_75t_L g5074 ( 
.A(n_4571),
.B(n_4215),
.Y(n_5074)
);

INVx1_ASAP7_75t_L g5075 ( 
.A(n_4454),
.Y(n_5075)
);

INVx2_ASAP7_75t_SL g5076 ( 
.A(n_4649),
.Y(n_5076)
);

INVx3_ASAP7_75t_L g5077 ( 
.A(n_4440),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_L g5078 ( 
.A(n_4744),
.B(n_4367),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_4462),
.Y(n_5079)
);

AND2x2_ASAP7_75t_L g5080 ( 
.A(n_4571),
.B(n_4215),
.Y(n_5080)
);

HB1xp67_ASAP7_75t_L g5081 ( 
.A(n_4470),
.Y(n_5081)
);

AND2x4_ASAP7_75t_L g5082 ( 
.A(n_4812),
.B(n_4874),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_4462),
.Y(n_5083)
);

AND2x2_ASAP7_75t_L g5084 ( 
.A(n_4812),
.B(n_4215),
.Y(n_5084)
);

NAND2xp5_ASAP7_75t_L g5085 ( 
.A(n_4572),
.B(n_4633),
.Y(n_5085)
);

OAI21x1_ASAP7_75t_L g5086 ( 
.A1(n_4440),
.A2(n_3934),
.B(n_3912),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4463),
.Y(n_5087)
);

OR2x2_ASAP7_75t_L g5088 ( 
.A(n_4522),
.B(n_4305),
.Y(n_5088)
);

NAND2x1_ASAP7_75t_L g5089 ( 
.A(n_4440),
.B(n_4407),
.Y(n_5089)
);

OAI21x1_ASAP7_75t_L g5090 ( 
.A1(n_4440),
.A2(n_4066),
.B(n_4065),
.Y(n_5090)
);

AO21x1_ASAP7_75t_SL g5091 ( 
.A1(n_4898),
.A2(n_4285),
.B(n_4282),
.Y(n_5091)
);

AND2x2_ASAP7_75t_L g5092 ( 
.A(n_4812),
.B(n_4215),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4463),
.Y(n_5093)
);

HB1xp67_ASAP7_75t_L g5094 ( 
.A(n_4490),
.Y(n_5094)
);

BUFx2_ASAP7_75t_L g5095 ( 
.A(n_4651),
.Y(n_5095)
);

INVx2_ASAP7_75t_L g5096 ( 
.A(n_4556),
.Y(n_5096)
);

HB1xp67_ASAP7_75t_L g5097 ( 
.A(n_4494),
.Y(n_5097)
);

AND2x2_ASAP7_75t_L g5098 ( 
.A(n_4812),
.B(n_4407),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4464),
.Y(n_5099)
);

AND2x2_ASAP7_75t_L g5100 ( 
.A(n_4874),
.B(n_4407),
.Y(n_5100)
);

OR2x2_ASAP7_75t_L g5101 ( 
.A(n_4573),
.B(n_4311),
.Y(n_5101)
);

AND2x2_ASAP7_75t_L g5102 ( 
.A(n_4874),
.B(n_4407),
.Y(n_5102)
);

OA21x2_ASAP7_75t_L g5103 ( 
.A1(n_4705),
.A2(n_3958),
.B(n_3946),
.Y(n_5103)
);

AO21x2_ASAP7_75t_L g5104 ( 
.A1(n_4542),
.A2(n_3959),
.B(n_3958),
.Y(n_5104)
);

INVx2_ASAP7_75t_L g5105 ( 
.A(n_4557),
.Y(n_5105)
);

INVx2_ASAP7_75t_L g5106 ( 
.A(n_4557),
.Y(n_5106)
);

AND2x2_ASAP7_75t_L g5107 ( 
.A(n_4874),
.B(n_4067),
.Y(n_5107)
);

INVx2_ASAP7_75t_L g5108 ( 
.A(n_4557),
.Y(n_5108)
);

INVx2_ASAP7_75t_L g5109 ( 
.A(n_4559),
.Y(n_5109)
);

INVx2_ASAP7_75t_L g5110 ( 
.A(n_4559),
.Y(n_5110)
);

INVx2_ASAP7_75t_L g5111 ( 
.A(n_4559),
.Y(n_5111)
);

OR2x2_ASAP7_75t_L g5112 ( 
.A(n_4593),
.B(n_4311),
.Y(n_5112)
);

AO31x2_ASAP7_75t_L g5113 ( 
.A1(n_4618),
.A2(n_3959),
.A3(n_4131),
.B(n_4124),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_4637),
.B(n_4188),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4464),
.Y(n_5115)
);

AND2x2_ASAP7_75t_L g5116 ( 
.A(n_4687),
.B(n_4067),
.Y(n_5116)
);

AO21x2_ASAP7_75t_L g5117 ( 
.A1(n_4542),
.A2(n_4004),
.B(n_4002),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_4467),
.Y(n_5118)
);

AO21x2_ASAP7_75t_L g5119 ( 
.A1(n_4720),
.A2(n_4004),
.B(n_4002),
.Y(n_5119)
);

AO21x2_ASAP7_75t_L g5120 ( 
.A1(n_4720),
.A2(n_4006),
.B(n_4162),
.Y(n_5120)
);

INVx3_ASAP7_75t_L g5121 ( 
.A(n_4450),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4467),
.Y(n_5122)
);

INVx1_ASAP7_75t_L g5123 ( 
.A(n_4476),
.Y(n_5123)
);

INVx3_ASAP7_75t_L g5124 ( 
.A(n_4450),
.Y(n_5124)
);

HB1xp67_ASAP7_75t_L g5125 ( 
.A(n_4498),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_4476),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_4478),
.Y(n_5127)
);

INVx2_ASAP7_75t_L g5128 ( 
.A(n_4566),
.Y(n_5128)
);

HB1xp67_ASAP7_75t_L g5129 ( 
.A(n_4569),
.Y(n_5129)
);

INVx2_ASAP7_75t_L g5130 ( 
.A(n_4566),
.Y(n_5130)
);

HB1xp67_ASAP7_75t_L g5131 ( 
.A(n_4839),
.Y(n_5131)
);

BUFx3_ASAP7_75t_L g5132 ( 
.A(n_4424),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_4478),
.Y(n_5133)
);

AO21x2_ASAP7_75t_L g5134 ( 
.A1(n_4720),
.A2(n_4006),
.B(n_4162),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_4479),
.Y(n_5135)
);

INVx2_ASAP7_75t_L g5136 ( 
.A(n_4566),
.Y(n_5136)
);

HB1xp67_ASAP7_75t_SL g5137 ( 
.A(n_4548),
.Y(n_5137)
);

OR2x2_ASAP7_75t_L g5138 ( 
.A(n_4785),
.B(n_4313),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_4479),
.Y(n_5139)
);

NOR2xp33_ASAP7_75t_L g5140 ( 
.A(n_4709),
.B(n_4819),
.Y(n_5140)
);

INVx1_ASAP7_75t_SL g5141 ( 
.A(n_4485),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_4488),
.Y(n_5142)
);

INVx3_ASAP7_75t_L g5143 ( 
.A(n_4450),
.Y(n_5143)
);

AND2x2_ASAP7_75t_L g5144 ( 
.A(n_4554),
.B(n_4069),
.Y(n_5144)
);

OA21x2_ASAP7_75t_L g5145 ( 
.A1(n_4524),
.A2(n_4395),
.B(n_3977),
.Y(n_5145)
);

OAI21xp5_ASAP7_75t_L g5146 ( 
.A1(n_4701),
.A2(n_4758),
.B(n_4703),
.Y(n_5146)
);

INVx2_ASAP7_75t_L g5147 ( 
.A(n_4567),
.Y(n_5147)
);

INVx2_ASAP7_75t_L g5148 ( 
.A(n_4567),
.Y(n_5148)
);

INVx2_ASAP7_75t_L g5149 ( 
.A(n_4567),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_4488),
.Y(n_5150)
);

OA21x2_ASAP7_75t_L g5151 ( 
.A1(n_4524),
.A2(n_4395),
.B(n_3977),
.Y(n_5151)
);

AOI21xp5_ASAP7_75t_L g5152 ( 
.A1(n_4497),
.A2(n_4853),
.B(n_4916),
.Y(n_5152)
);

INVx3_ASAP7_75t_L g5153 ( 
.A(n_4450),
.Y(n_5153)
);

BUFx2_ASAP7_75t_L g5154 ( 
.A(n_4651),
.Y(n_5154)
);

NOR2xp33_ASAP7_75t_L g5155 ( 
.A(n_4709),
.B(n_4239),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4489),
.Y(n_5156)
);

AO21x2_ASAP7_75t_L g5157 ( 
.A1(n_4568),
.A2(n_4296),
.B(n_4344),
.Y(n_5157)
);

AND2x2_ASAP7_75t_L g5158 ( 
.A(n_4554),
.B(n_4069),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_4489),
.Y(n_5159)
);

INVx3_ASAP7_75t_L g5160 ( 
.A(n_4461),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_4492),
.Y(n_5161)
);

INVxp67_ASAP7_75t_SL g5162 ( 
.A(n_4877),
.Y(n_5162)
);

BUFx2_ASAP7_75t_L g5163 ( 
.A(n_4651),
.Y(n_5163)
);

INVx2_ASAP7_75t_L g5164 ( 
.A(n_4568),
.Y(n_5164)
);

INVx2_ASAP7_75t_L g5165 ( 
.A(n_4568),
.Y(n_5165)
);

OR2x2_ASAP7_75t_L g5166 ( 
.A(n_4629),
.B(n_4313),
.Y(n_5166)
);

BUFx2_ASAP7_75t_L g5167 ( 
.A(n_4677),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_4560),
.B(n_4111),
.Y(n_5168)
);

INVx2_ASAP7_75t_L g5169 ( 
.A(n_4433),
.Y(n_5169)
);

OA21x2_ASAP7_75t_L g5170 ( 
.A1(n_4506),
.A2(n_3962),
.B(n_4303),
.Y(n_5170)
);

BUFx2_ASAP7_75t_L g5171 ( 
.A(n_4677),
.Y(n_5171)
);

INVx1_ASAP7_75t_SL g5172 ( 
.A(n_4541),
.Y(n_5172)
);

HB1xp67_ASAP7_75t_L g5173 ( 
.A(n_4617),
.Y(n_5173)
);

INVx2_ASAP7_75t_L g5174 ( 
.A(n_4433),
.Y(n_5174)
);

INVx1_ASAP7_75t_L g5175 ( 
.A(n_4492),
.Y(n_5175)
);

AO21x2_ASAP7_75t_L g5176 ( 
.A1(n_4576),
.A2(n_4344),
.B(n_4319),
.Y(n_5176)
);

OAI21x1_ASAP7_75t_L g5177 ( 
.A1(n_4461),
.A2(n_4066),
.B(n_4065),
.Y(n_5177)
);

HB1xp67_ASAP7_75t_L g5178 ( 
.A(n_4660),
.Y(n_5178)
);

HB1xp67_ASAP7_75t_L g5179 ( 
.A(n_4665),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_4495),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_4802),
.B(n_4188),
.Y(n_5181)
);

OR2x2_ASAP7_75t_L g5182 ( 
.A(n_4876),
.B(n_4320),
.Y(n_5182)
);

INVx3_ASAP7_75t_L g5183 ( 
.A(n_4461),
.Y(n_5183)
);

BUFx6f_ASAP7_75t_L g5184 ( 
.A(n_4481),
.Y(n_5184)
);

AO21x2_ASAP7_75t_L g5185 ( 
.A1(n_4576),
.A2(n_4319),
.B(n_4303),
.Y(n_5185)
);

AND2x2_ASAP7_75t_L g5186 ( 
.A(n_4560),
.B(n_4111),
.Y(n_5186)
);

INVx3_ASAP7_75t_L g5187 ( 
.A(n_4461),
.Y(n_5187)
);

HB1xp67_ASAP7_75t_L g5188 ( 
.A(n_4692),
.Y(n_5188)
);

AND2x2_ASAP7_75t_L g5189 ( 
.A(n_4596),
.B(n_4127),
.Y(n_5189)
);

HB1xp67_ASAP7_75t_L g5190 ( 
.A(n_4544),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_4495),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_4496),
.Y(n_5192)
);

INVx2_ASAP7_75t_L g5193 ( 
.A(n_4433),
.Y(n_5193)
);

INVx2_ASAP7_75t_L g5194 ( 
.A(n_4443),
.Y(n_5194)
);

INVx2_ASAP7_75t_L g5195 ( 
.A(n_4443),
.Y(n_5195)
);

AND2x4_ASAP7_75t_L g5196 ( 
.A(n_4503),
.B(n_4074),
.Y(n_5196)
);

AO21x2_ASAP7_75t_L g5197 ( 
.A1(n_4576),
.A2(n_4339),
.B(n_4403),
.Y(n_5197)
);

INVx3_ASAP7_75t_L g5198 ( 
.A(n_4491),
.Y(n_5198)
);

BUFx2_ASAP7_75t_L g5199 ( 
.A(n_4677),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_4643),
.B(n_4227),
.Y(n_5200)
);

INVx2_ASAP7_75t_L g5201 ( 
.A(n_4443),
.Y(n_5201)
);

AND2x2_ASAP7_75t_L g5202 ( 
.A(n_4596),
.B(n_4127),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_4496),
.Y(n_5203)
);

HB1xp67_ASAP7_75t_L g5204 ( 
.A(n_4544),
.Y(n_5204)
);

OR2x2_ASAP7_75t_L g5205 ( 
.A(n_4810),
.B(n_4320),
.Y(n_5205)
);

INVx3_ASAP7_75t_L g5206 ( 
.A(n_4491),
.Y(n_5206)
);

INVx3_ASAP7_75t_L g5207 ( 
.A(n_4491),
.Y(n_5207)
);

OA21x2_ASAP7_75t_L g5208 ( 
.A1(n_4506),
.A2(n_3962),
.B(n_4339),
.Y(n_5208)
);

AND2x2_ASAP7_75t_L g5209 ( 
.A(n_4602),
.B(n_4135),
.Y(n_5209)
);

OR2x2_ASAP7_75t_L g5210 ( 
.A(n_4810),
.B(n_4878),
.Y(n_5210)
);

INVx4_ASAP7_75t_SL g5211 ( 
.A(n_4713),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_4500),
.Y(n_5212)
);

INVx5_ASAP7_75t_L g5213 ( 
.A(n_4491),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_4458),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_4500),
.Y(n_5215)
);

AOI22xp33_ASAP7_75t_L g5216 ( 
.A1(n_4453),
.A2(n_4316),
.B1(n_3926),
.B2(n_3825),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_4643),
.B(n_4227),
.Y(n_5217)
);

INVx2_ASAP7_75t_L g5218 ( 
.A(n_4458),
.Y(n_5218)
);

INVx1_ASAP7_75t_L g5219 ( 
.A(n_4510),
.Y(n_5219)
);

OAI21x1_ASAP7_75t_L g5220 ( 
.A1(n_4518),
.A2(n_4066),
.B(n_4065),
.Y(n_5220)
);

INVx2_ASAP7_75t_SL g5221 ( 
.A(n_4713),
.Y(n_5221)
);

AND2x4_ASAP7_75t_L g5222 ( 
.A(n_4503),
.B(n_4074),
.Y(n_5222)
);

AO21x2_ASAP7_75t_L g5223 ( 
.A1(n_4701),
.A2(n_4410),
.B(n_4403),
.Y(n_5223)
);

INVx2_ASAP7_75t_L g5224 ( 
.A(n_4458),
.Y(n_5224)
);

INVx2_ASAP7_75t_L g5225 ( 
.A(n_4459),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_4510),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_4511),
.Y(n_5227)
);

INVx2_ASAP7_75t_L g5228 ( 
.A(n_4459),
.Y(n_5228)
);

AO21x2_ASAP7_75t_L g5229 ( 
.A1(n_4751),
.A2(n_4411),
.B(n_4410),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_L g5230 ( 
.A(n_4793),
.B(n_4237),
.Y(n_5230)
);

AO21x2_ASAP7_75t_L g5231 ( 
.A1(n_4751),
.A2(n_4412),
.B(n_4411),
.Y(n_5231)
);

OR2x6_ASAP7_75t_L g5232 ( 
.A(n_4694),
.B(n_4399),
.Y(n_5232)
);

INVx2_ASAP7_75t_L g5233 ( 
.A(n_4459),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_4511),
.Y(n_5234)
);

NAND2xp5_ASAP7_75t_L g5235 ( 
.A(n_4793),
.B(n_4237),
.Y(n_5235)
);

HB1xp67_ASAP7_75t_L g5236 ( 
.A(n_4578),
.Y(n_5236)
);

AO21x2_ASAP7_75t_L g5237 ( 
.A1(n_4545),
.A2(n_4412),
.B(n_4131),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_4420),
.Y(n_5238)
);

AND2x2_ASAP7_75t_L g5239 ( 
.A(n_4602),
.B(n_4135),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_4516),
.Y(n_5240)
);

OA21x2_ASAP7_75t_L g5241 ( 
.A1(n_4527),
.A2(n_4131),
.B(n_4124),
.Y(n_5241)
);

AO21x2_ASAP7_75t_L g5242 ( 
.A1(n_4545),
.A2(n_4138),
.B(n_4124),
.Y(n_5242)
);

INVxp67_ASAP7_75t_SL g5243 ( 
.A(n_4646),
.Y(n_5243)
);

INVx2_ASAP7_75t_L g5244 ( 
.A(n_4420),
.Y(n_5244)
);

INVx2_ASAP7_75t_SL g5245 ( 
.A(n_4713),
.Y(n_5245)
);

INVx2_ASAP7_75t_SL g5246 ( 
.A(n_4548),
.Y(n_5246)
);

AND2x2_ASAP7_75t_L g5247 ( 
.A(n_4604),
.B(n_4023),
.Y(n_5247)
);

INVx2_ASAP7_75t_L g5248 ( 
.A(n_4426),
.Y(n_5248)
);

OR2x6_ASAP7_75t_L g5249 ( 
.A(n_4694),
.B(n_4399),
.Y(n_5249)
);

INVx2_ASAP7_75t_L g5250 ( 
.A(n_4426),
.Y(n_5250)
);

AND2x2_ASAP7_75t_L g5251 ( 
.A(n_4604),
.B(n_4627),
.Y(n_5251)
);

OR2x6_ASAP7_75t_L g5252 ( 
.A(n_4694),
.B(n_4263),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_4840),
.B(n_4326),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_4516),
.Y(n_5254)
);

AO21x2_ASAP7_75t_L g5255 ( 
.A1(n_4550),
.A2(n_4146),
.B(n_4138),
.Y(n_5255)
);

BUFx3_ASAP7_75t_L g5256 ( 
.A(n_4548),
.Y(n_5256)
);

INVx2_ASAP7_75t_L g5257 ( 
.A(n_4427),
.Y(n_5257)
);

AND2x4_ASAP7_75t_L g5258 ( 
.A(n_4503),
.B(n_4611),
.Y(n_5258)
);

INVx2_ASAP7_75t_L g5259 ( 
.A(n_4427),
.Y(n_5259)
);

INVx1_ASAP7_75t_L g5260 ( 
.A(n_4517),
.Y(n_5260)
);

INVx1_ASAP7_75t_SL g5261 ( 
.A(n_4466),
.Y(n_5261)
);

NAND2xp5_ASAP7_75t_L g5262 ( 
.A(n_4840),
.B(n_4326),
.Y(n_5262)
);

AO21x2_ASAP7_75t_L g5263 ( 
.A1(n_4550),
.A2(n_4553),
.B(n_4435),
.Y(n_5263)
);

AND2x2_ASAP7_75t_L g5264 ( 
.A(n_4627),
.B(n_4023),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_4517),
.Y(n_5265)
);

BUFx6f_ASAP7_75t_L g5266 ( 
.A(n_4481),
.Y(n_5266)
);

OR2x6_ASAP7_75t_L g5267 ( 
.A(n_4763),
.B(n_4263),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_4520),
.Y(n_5268)
);

INVx2_ASAP7_75t_L g5269 ( 
.A(n_4429),
.Y(n_5269)
);

INVx2_ASAP7_75t_L g5270 ( 
.A(n_4429),
.Y(n_5270)
);

AO21x2_ASAP7_75t_L g5271 ( 
.A1(n_4553),
.A2(n_4146),
.B(n_4138),
.Y(n_5271)
);

BUFx3_ASAP7_75t_L g5272 ( 
.A(n_4548),
.Y(n_5272)
);

INVx1_ASAP7_75t_L g5273 ( 
.A(n_4520),
.Y(n_5273)
);

INVx2_ASAP7_75t_L g5274 ( 
.A(n_4435),
.Y(n_5274)
);

OAI21xp5_ASAP7_75t_L g5275 ( 
.A1(n_4776),
.A2(n_3925),
.B(n_4360),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_4525),
.Y(n_5276)
);

INVx3_ASAP7_75t_L g5277 ( 
.A(n_4518),
.Y(n_5277)
);

INVx2_ASAP7_75t_L g5278 ( 
.A(n_4455),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_4525),
.Y(n_5279)
);

INVx2_ASAP7_75t_L g5280 ( 
.A(n_4455),
.Y(n_5280)
);

INVx2_ASAP7_75t_L g5281 ( 
.A(n_4474),
.Y(n_5281)
);

INVx2_ASAP7_75t_L g5282 ( 
.A(n_4474),
.Y(n_5282)
);

INVx2_ASAP7_75t_L g5283 ( 
.A(n_4477),
.Y(n_5283)
);

AND2x2_ASAP7_75t_L g5284 ( 
.A(n_4695),
.B(n_4028),
.Y(n_5284)
);

AND2x2_ASAP7_75t_L g5285 ( 
.A(n_4695),
.B(n_4028),
.Y(n_5285)
);

INVxp67_ASAP7_75t_L g5286 ( 
.A(n_4436),
.Y(n_5286)
);

INVx2_ASAP7_75t_L g5287 ( 
.A(n_4477),
.Y(n_5287)
);

NAND2xp5_ASAP7_75t_L g5288 ( 
.A(n_4878),
.B(n_4329),
.Y(n_5288)
);

INVx3_ASAP7_75t_L g5289 ( 
.A(n_4518),
.Y(n_5289)
);

OR2x6_ASAP7_75t_L g5290 ( 
.A(n_4763),
.B(n_4263),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_4714),
.B(n_4063),
.Y(n_5291)
);

INVx2_ASAP7_75t_L g5292 ( 
.A(n_4672),
.Y(n_5292)
);

OR2x2_ASAP7_75t_L g5293 ( 
.A(n_4907),
.B(n_4329),
.Y(n_5293)
);

AO21x2_ASAP7_75t_L g5294 ( 
.A1(n_4469),
.A2(n_4789),
.B(n_4672),
.Y(n_5294)
);

INVx2_ASAP7_75t_L g5295 ( 
.A(n_4672),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_4529),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_4529),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_4530),
.Y(n_5298)
);

OAI21xp5_ASAP7_75t_L g5299 ( 
.A1(n_4518),
.A2(n_4253),
.B(n_4086),
.Y(n_5299)
);

OAI21x1_ASAP7_75t_L g5300 ( 
.A1(n_4531),
.A2(n_4086),
.B(n_4066),
.Y(n_5300)
);

INVx2_ASAP7_75t_L g5301 ( 
.A(n_4789),
.Y(n_5301)
);

INVx1_ASAP7_75t_SL g5302 ( 
.A(n_4499),
.Y(n_5302)
);

BUFx2_ASAP7_75t_L g5303 ( 
.A(n_4523),
.Y(n_5303)
);

AO21x2_ASAP7_75t_L g5304 ( 
.A1(n_4469),
.A2(n_4164),
.B(n_4146),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4530),
.Y(n_5305)
);

OR2x2_ASAP7_75t_L g5306 ( 
.A(n_4907),
.B(n_4330),
.Y(n_5306)
);

NOR2xp33_ASAP7_75t_L g5307 ( 
.A(n_4697),
.B(n_4168),
.Y(n_5307)
);

AND2x4_ASAP7_75t_L g5308 ( 
.A(n_4503),
.B(n_4074),
.Y(n_5308)
);

INVx2_ASAP7_75t_L g5309 ( 
.A(n_4789),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_4533),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_4533),
.Y(n_5311)
);

OR2x2_ASAP7_75t_L g5312 ( 
.A(n_4534),
.B(n_4330),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_4534),
.Y(n_5313)
);

AOI222xp33_ASAP7_75t_L g5314 ( 
.A1(n_4668),
.A2(n_4382),
.B1(n_4371),
.B2(n_3826),
.C1(n_3836),
.C2(n_3825),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_4519),
.B(n_4345),
.Y(n_5315)
);

INVx2_ASAP7_75t_L g5316 ( 
.A(n_4794),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_4535),
.Y(n_5317)
);

NAND2xp5_ASAP7_75t_L g5318 ( 
.A(n_4519),
.B(n_4345),
.Y(n_5318)
);

NOR2xp67_ASAP7_75t_L g5319 ( 
.A(n_4442),
.B(n_4086),
.Y(n_5319)
);

OA21x2_ASAP7_75t_L g5320 ( 
.A1(n_4527),
.A2(n_4166),
.B(n_4164),
.Y(n_5320)
);

INVx2_ASAP7_75t_L g5321 ( 
.A(n_4794),
.Y(n_5321)
);

INVx2_ASAP7_75t_L g5322 ( 
.A(n_4794),
.Y(n_5322)
);

AND2x2_ASAP7_75t_L g5323 ( 
.A(n_4714),
.B(n_4063),
.Y(n_5323)
);

INVxp67_ASAP7_75t_SL g5324 ( 
.A(n_4646),
.Y(n_5324)
);

INVxp67_ASAP7_75t_SL g5325 ( 
.A(n_4646),
.Y(n_5325)
);

INVx2_ASAP7_75t_L g5326 ( 
.A(n_4798),
.Y(n_5326)
);

HB1xp67_ASAP7_75t_L g5327 ( 
.A(n_4578),
.Y(n_5327)
);

AND2x2_ASAP7_75t_L g5328 ( 
.A(n_4716),
.B(n_4310),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_4519),
.B(n_4349),
.Y(n_5329)
);

OR2x2_ASAP7_75t_L g5330 ( 
.A(n_4535),
.B(n_4349),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_4537),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_4537),
.Y(n_5332)
);

INVx2_ASAP7_75t_L g5333 ( 
.A(n_4798),
.Y(n_5333)
);

AO21x2_ASAP7_75t_L g5334 ( 
.A1(n_4469),
.A2(n_4166),
.B(n_4164),
.Y(n_5334)
);

OR2x6_ASAP7_75t_L g5335 ( 
.A(n_4763),
.B(n_3926),
.Y(n_5335)
);

AO21x2_ASAP7_75t_L g5336 ( 
.A1(n_4798),
.A2(n_4170),
.B(n_4166),
.Y(n_5336)
);

INVx2_ASAP7_75t_L g5337 ( 
.A(n_4800),
.Y(n_5337)
);

INVx2_ASAP7_75t_L g5338 ( 
.A(n_4800),
.Y(n_5338)
);

INVx2_ASAP7_75t_SL g5339 ( 
.A(n_4481),
.Y(n_5339)
);

AOI21x1_ASAP7_75t_L g5340 ( 
.A1(n_4787),
.A2(n_4189),
.B(n_4385),
.Y(n_5340)
);

AND2x2_ASAP7_75t_L g5341 ( 
.A(n_4716),
.B(n_4310),
.Y(n_5341)
);

OA21x2_ASAP7_75t_L g5342 ( 
.A1(n_4502),
.A2(n_4172),
.B(n_4170),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_4538),
.Y(n_5343)
);

NAND2xp5_ASAP7_75t_L g5344 ( 
.A(n_4519),
.B(n_4352),
.Y(n_5344)
);

AND2x2_ASAP7_75t_L g5345 ( 
.A(n_4739),
.B(n_4346),
.Y(n_5345)
);

BUFx12f_ASAP7_75t_L g5346 ( 
.A(n_4523),
.Y(n_5346)
);

INVx3_ASAP7_75t_L g5347 ( 
.A(n_4531),
.Y(n_5347)
);

NOR2xp33_ASAP7_75t_L g5348 ( 
.A(n_5043),
.B(n_4745),
.Y(n_5348)
);

INVx2_ASAP7_75t_L g5349 ( 
.A(n_5294),
.Y(n_5349)
);

BUFx6f_ASAP7_75t_L g5350 ( 
.A(n_4927),
.Y(n_5350)
);

INVx2_ASAP7_75t_L g5351 ( 
.A(n_5294),
.Y(n_5351)
);

OR2x2_ASAP7_75t_L g5352 ( 
.A(n_5210),
.B(n_4588),
.Y(n_5352)
);

INVx2_ASAP7_75t_L g5353 ( 
.A(n_5294),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5131),
.Y(n_5354)
);

AOI22xp33_ASAP7_75t_L g5355 ( 
.A1(n_5146),
.A2(n_4536),
.B1(n_4531),
.B2(n_4618),
.Y(n_5355)
);

AND2x2_ASAP7_75t_L g5356 ( 
.A(n_4930),
.B(n_4588),
.Y(n_5356)
);

AND2x2_ASAP7_75t_L g5357 ( 
.A(n_4930),
.B(n_4610),
.Y(n_5357)
);

INVx2_ASAP7_75t_L g5358 ( 
.A(n_5117),
.Y(n_5358)
);

NAND2xp5_ASAP7_75t_L g5359 ( 
.A(n_5162),
.B(n_4519),
.Y(n_5359)
);

AND2x2_ASAP7_75t_L g5360 ( 
.A(n_4933),
.B(n_4610),
.Y(n_5360)
);

HB1xp67_ASAP7_75t_L g5361 ( 
.A(n_5190),
.Y(n_5361)
);

NAND2xp5_ASAP7_75t_L g5362 ( 
.A(n_5173),
.B(n_4519),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_4980),
.Y(n_5363)
);

OR2x2_ASAP7_75t_L g5364 ( 
.A(n_5210),
.B(n_4762),
.Y(n_5364)
);

OR2x2_ASAP7_75t_L g5365 ( 
.A(n_5036),
.B(n_5066),
.Y(n_5365)
);

AND2x2_ASAP7_75t_L g5366 ( 
.A(n_4933),
.B(n_4558),
.Y(n_5366)
);

INVx1_ASAP7_75t_L g5367 ( 
.A(n_4980),
.Y(n_5367)
);

NAND2xp5_ASAP7_75t_L g5368 ( 
.A(n_4954),
.B(n_4558),
.Y(n_5368)
);

INVx1_ASAP7_75t_L g5369 ( 
.A(n_4981),
.Y(n_5369)
);

AOI22xp33_ASAP7_75t_L g5370 ( 
.A1(n_4938),
.A2(n_4536),
.B1(n_4531),
.B2(n_4641),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_4981),
.Y(n_5371)
);

INVx2_ASAP7_75t_L g5372 ( 
.A(n_5117),
.Y(n_5372)
);

BUFx2_ASAP7_75t_SL g5373 ( 
.A(n_4927),
.Y(n_5373)
);

INVx2_ASAP7_75t_SL g5374 ( 
.A(n_4965),
.Y(n_5374)
);

AND2x4_ASAP7_75t_L g5375 ( 
.A(n_4985),
.B(n_4699),
.Y(n_5375)
);

INVx1_ASAP7_75t_L g5376 ( 
.A(n_4982),
.Y(n_5376)
);

OR2x2_ASAP7_75t_L g5377 ( 
.A(n_5036),
.B(n_4431),
.Y(n_5377)
);

INVx1_ASAP7_75t_L g5378 ( 
.A(n_4982),
.Y(n_5378)
);

OR2x2_ASAP7_75t_L g5379 ( 
.A(n_5066),
.B(n_4431),
.Y(n_5379)
);

AND2x2_ASAP7_75t_L g5380 ( 
.A(n_4955),
.B(n_4558),
.Y(n_5380)
);

AND2x4_ASAP7_75t_SL g5381 ( 
.A(n_4994),
.B(n_3982),
.Y(n_5381)
);

INVxp67_ASAP7_75t_L g5382 ( 
.A(n_5303),
.Y(n_5382)
);

AND2x2_ASAP7_75t_L g5383 ( 
.A(n_4955),
.B(n_4966),
.Y(n_5383)
);

AND2x4_ASAP7_75t_SL g5384 ( 
.A(n_4994),
.B(n_4001),
.Y(n_5384)
);

INVx2_ASAP7_75t_L g5385 ( 
.A(n_5117),
.Y(n_5385)
);

BUFx2_ASAP7_75t_L g5386 ( 
.A(n_5346),
.Y(n_5386)
);

INVx2_ASAP7_75t_L g5387 ( 
.A(n_5304),
.Y(n_5387)
);

INVx2_ASAP7_75t_L g5388 ( 
.A(n_5304),
.Y(n_5388)
);

NAND2xp5_ASAP7_75t_L g5389 ( 
.A(n_4935),
.B(n_4558),
.Y(n_5389)
);

NAND2xp33_ASAP7_75t_R g5390 ( 
.A(n_5303),
.B(n_4828),
.Y(n_5390)
);

OR2x2_ASAP7_75t_L g5391 ( 
.A(n_5166),
.B(n_4448),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_4984),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_4984),
.Y(n_5393)
);

AOI22xp5_ASAP7_75t_L g5394 ( 
.A1(n_4938),
.A2(n_4551),
.B1(n_4441),
.B2(n_4885),
.Y(n_5394)
);

INVx2_ASAP7_75t_L g5395 ( 
.A(n_5304),
.Y(n_5395)
);

BUFx2_ASAP7_75t_L g5396 ( 
.A(n_5346),
.Y(n_5396)
);

AND2x2_ASAP7_75t_L g5397 ( 
.A(n_4966),
.B(n_4558),
.Y(n_5397)
);

AND2x2_ASAP7_75t_L g5398 ( 
.A(n_4985),
.B(n_4558),
.Y(n_5398)
);

INVx2_ASAP7_75t_L g5399 ( 
.A(n_5334),
.Y(n_5399)
);

AND2x2_ASAP7_75t_L g5400 ( 
.A(n_5107),
.B(n_4613),
.Y(n_5400)
);

INVx2_ASAP7_75t_L g5401 ( 
.A(n_5334),
.Y(n_5401)
);

AND2x2_ASAP7_75t_L g5402 ( 
.A(n_5107),
.B(n_4613),
.Y(n_5402)
);

OR2x2_ASAP7_75t_L g5403 ( 
.A(n_5166),
.B(n_4448),
.Y(n_5403)
);

AND2x2_ASAP7_75t_L g5404 ( 
.A(n_5116),
.B(n_4613),
.Y(n_5404)
);

AND2x2_ASAP7_75t_L g5405 ( 
.A(n_5116),
.B(n_4613),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_4993),
.Y(n_5406)
);

INVx1_ASAP7_75t_L g5407 ( 
.A(n_4993),
.Y(n_5407)
);

INVx5_ASAP7_75t_L g5408 ( 
.A(n_4965),
.Y(n_5408)
);

HB1xp67_ASAP7_75t_L g5409 ( 
.A(n_5204),
.Y(n_5409)
);

CKINVDCx5p33_ASAP7_75t_R g5410 ( 
.A(n_4956),
.Y(n_5410)
);

OR2x2_ASAP7_75t_L g5411 ( 
.A(n_5288),
.B(n_4460),
.Y(n_5411)
);

INVx2_ASAP7_75t_L g5412 ( 
.A(n_5334),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_4997),
.Y(n_5413)
);

AND2x2_ASAP7_75t_L g5414 ( 
.A(n_5251),
.B(n_4613),
.Y(n_5414)
);

HB1xp67_ASAP7_75t_L g5415 ( 
.A(n_5236),
.Y(n_5415)
);

AND2x2_ASAP7_75t_L g5416 ( 
.A(n_5251),
.B(n_4613),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_4969),
.Y(n_5417)
);

OR2x2_ASAP7_75t_L g5418 ( 
.A(n_5085),
.B(n_4460),
.Y(n_5418)
);

NOR2x1p5_ASAP7_75t_L g5419 ( 
.A(n_5005),
.B(n_4483),
.Y(n_5419)
);

INVx2_ASAP7_75t_L g5420 ( 
.A(n_4969),
.Y(n_5420)
);

INVxp67_ASAP7_75t_SL g5421 ( 
.A(n_5286),
.Y(n_5421)
);

INVx2_ASAP7_75t_L g5422 ( 
.A(n_4969),
.Y(n_5422)
);

INVx2_ASAP7_75t_L g5423 ( 
.A(n_5014),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_4997),
.Y(n_5424)
);

NAND2xp5_ASAP7_75t_L g5425 ( 
.A(n_4976),
.B(n_4473),
.Y(n_5425)
);

OR2x2_ASAP7_75t_L g5426 ( 
.A(n_4946),
.B(n_4473),
.Y(n_5426)
);

INVx1_ASAP7_75t_L g5427 ( 
.A(n_5000),
.Y(n_5427)
);

AND2x2_ASAP7_75t_L g5428 ( 
.A(n_5082),
.B(n_4699),
.Y(n_5428)
);

OAI22xp5_ASAP7_75t_L g5429 ( 
.A1(n_5152),
.A2(n_4862),
.B1(n_4805),
.B2(n_4891),
.Y(n_5429)
);

INVx3_ASAP7_75t_L g5430 ( 
.A(n_5213),
.Y(n_5430)
);

INVx2_ASAP7_75t_L g5431 ( 
.A(n_5014),
.Y(n_5431)
);

INVx2_ASAP7_75t_L g5432 ( 
.A(n_5014),
.Y(n_5432)
);

NAND2xp5_ASAP7_75t_L g5433 ( 
.A(n_4990),
.B(n_4917),
.Y(n_5433)
);

NAND2xp5_ASAP7_75t_L g5434 ( 
.A(n_4991),
.B(n_4828),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5000),
.Y(n_5435)
);

BUFx2_ASAP7_75t_L g5436 ( 
.A(n_5005),
.Y(n_5436)
);

AND2x2_ASAP7_75t_L g5437 ( 
.A(n_5082),
.B(n_4699),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_5119),
.Y(n_5438)
);

AND2x2_ASAP7_75t_L g5439 ( 
.A(n_5082),
.B(n_4765),
.Y(n_5439)
);

INVx1_ASAP7_75t_L g5440 ( 
.A(n_5002),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_5002),
.Y(n_5441)
);

NOR2xp33_ASAP7_75t_L g5442 ( 
.A(n_4956),
.B(n_4745),
.Y(n_5442)
);

AND2x4_ASAP7_75t_L g5443 ( 
.A(n_5082),
.B(n_4765),
.Y(n_5443)
);

OR2x2_ASAP7_75t_L g5444 ( 
.A(n_4946),
.B(n_4919),
.Y(n_5444)
);

INVx1_ASAP7_75t_L g5445 ( 
.A(n_5008),
.Y(n_5445)
);

INVx1_ASAP7_75t_L g5446 ( 
.A(n_5008),
.Y(n_5446)
);

INVx2_ASAP7_75t_L g5447 ( 
.A(n_5119),
.Y(n_5447)
);

INVxp67_ASAP7_75t_SL g5448 ( 
.A(n_5132),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_5009),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_5009),
.Y(n_5450)
);

BUFx6f_ASAP7_75t_L g5451 ( 
.A(n_4965),
.Y(n_5451)
);

INVx2_ASAP7_75t_SL g5452 ( 
.A(n_4965),
.Y(n_5452)
);

BUFx2_ASAP7_75t_L g5453 ( 
.A(n_5132),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_5011),
.Y(n_5454)
);

NAND2x1_ASAP7_75t_L g5455 ( 
.A(n_5258),
.B(n_5196),
.Y(n_5455)
);

INVx3_ASAP7_75t_L g5456 ( 
.A(n_5213),
.Y(n_5456)
);

NOR2xp33_ASAP7_75t_L g5457 ( 
.A(n_4965),
.B(n_4745),
.Y(n_5457)
);

OAI222xp33_ASAP7_75t_L g5458 ( 
.A1(n_5042),
.A2(n_4796),
.B1(n_4887),
.B2(n_4641),
.C1(n_4664),
.C2(n_4763),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_5144),
.B(n_4765),
.Y(n_5459)
);

AND2x2_ASAP7_75t_L g5460 ( 
.A(n_5144),
.B(n_4765),
.Y(n_5460)
);

AND2x2_ASAP7_75t_L g5461 ( 
.A(n_5158),
.B(n_4842),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_5011),
.Y(n_5462)
);

BUFx2_ASAP7_75t_L g5463 ( 
.A(n_5256),
.Y(n_5463)
);

AND2x2_ASAP7_75t_L g5464 ( 
.A(n_5158),
.B(n_5168),
.Y(n_5464)
);

AND2x4_ASAP7_75t_L g5465 ( 
.A(n_5258),
.B(n_4846),
.Y(n_5465)
);

INVx2_ASAP7_75t_L g5466 ( 
.A(n_5119),
.Y(n_5466)
);

NAND2xp5_ASAP7_75t_L g5467 ( 
.A(n_5004),
.B(n_4842),
.Y(n_5467)
);

INVx2_ASAP7_75t_L g5468 ( 
.A(n_4928),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_5019),
.Y(n_5469)
);

AND2x2_ASAP7_75t_L g5470 ( 
.A(n_5168),
.B(n_4922),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_5019),
.Y(n_5471)
);

OAI21x1_ASAP7_75t_L g5472 ( 
.A1(n_5018),
.A2(n_4755),
.B(n_4547),
.Y(n_5472)
);

AND2x2_ASAP7_75t_L g5473 ( 
.A(n_5186),
.B(n_4922),
.Y(n_5473)
);

INVx4_ASAP7_75t_SL g5474 ( 
.A(n_5256),
.Y(n_5474)
);

INVx2_ASAP7_75t_L g5475 ( 
.A(n_4928),
.Y(n_5475)
);

AOI22xp33_ASAP7_75t_L g5476 ( 
.A1(n_4938),
.A2(n_4664),
.B1(n_4434),
.B2(n_4486),
.Y(n_5476)
);

NAND2xp33_ASAP7_75t_R g5477 ( 
.A(n_4963),
.B(n_4628),
.Y(n_5477)
);

INVx2_ASAP7_75t_L g5478 ( 
.A(n_4929),
.Y(n_5478)
);

INVx1_ASAP7_75t_L g5479 ( 
.A(n_5021),
.Y(n_5479)
);

INVx2_ASAP7_75t_L g5480 ( 
.A(n_4929),
.Y(n_5480)
);

HB1xp67_ASAP7_75t_L g5481 ( 
.A(n_5327),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_5021),
.Y(n_5482)
);

INVx2_ASAP7_75t_L g5483 ( 
.A(n_4934),
.Y(n_5483)
);

INVx2_ASAP7_75t_L g5484 ( 
.A(n_4934),
.Y(n_5484)
);

AND2x2_ASAP7_75t_L g5485 ( 
.A(n_5186),
.B(n_4646),
.Y(n_5485)
);

AND2x4_ASAP7_75t_L g5486 ( 
.A(n_5258),
.B(n_4846),
.Y(n_5486)
);

OR2x2_ASAP7_75t_L g5487 ( 
.A(n_4961),
.B(n_4926),
.Y(n_5487)
);

NAND2xp5_ASAP7_75t_L g5488 ( 
.A(n_5006),
.B(n_4597),
.Y(n_5488)
);

AOI21xp33_ASAP7_75t_L g5489 ( 
.A1(n_5223),
.A2(n_4442),
.B(n_4763),
.Y(n_5489)
);

INVx2_ASAP7_75t_L g5490 ( 
.A(n_4947),
.Y(n_5490)
);

HB1xp67_ASAP7_75t_L g5491 ( 
.A(n_5016),
.Y(n_5491)
);

NAND2xp5_ASAP7_75t_L g5492 ( 
.A(n_5081),
.B(n_4546),
.Y(n_5492)
);

INVx3_ASAP7_75t_L g5493 ( 
.A(n_5213),
.Y(n_5493)
);

OR2x2_ASAP7_75t_L g5494 ( 
.A(n_4961),
.B(n_4909),
.Y(n_5494)
);

AND2x2_ASAP7_75t_L g5495 ( 
.A(n_5189),
.B(n_4646),
.Y(n_5495)
);

INVx3_ASAP7_75t_L g5496 ( 
.A(n_5213),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_5024),
.Y(n_5497)
);

NAND2xp5_ASAP7_75t_L g5498 ( 
.A(n_5094),
.B(n_4449),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5024),
.Y(n_5499)
);

BUFx2_ASAP7_75t_L g5500 ( 
.A(n_5272),
.Y(n_5500)
);

INVx1_ASAP7_75t_L g5501 ( 
.A(n_5030),
.Y(n_5501)
);

NAND2xp5_ASAP7_75t_L g5502 ( 
.A(n_5097),
.B(n_4449),
.Y(n_5502)
);

HB1xp67_ASAP7_75t_L g5503 ( 
.A(n_5125),
.Y(n_5503)
);

OR2x2_ASAP7_75t_L g5504 ( 
.A(n_5205),
.B(n_4909),
.Y(n_5504)
);

OR2x2_ASAP7_75t_L g5505 ( 
.A(n_5205),
.B(n_4919),
.Y(n_5505)
);

INVx1_ASAP7_75t_L g5506 ( 
.A(n_5030),
.Y(n_5506)
);

NAND2x1_ASAP7_75t_L g5507 ( 
.A(n_5258),
.B(n_4679),
.Y(n_5507)
);

BUFx2_ASAP7_75t_L g5508 ( 
.A(n_5272),
.Y(n_5508)
);

NAND2xp5_ASAP7_75t_L g5509 ( 
.A(n_5129),
.B(n_5178),
.Y(n_5509)
);

AND2x2_ASAP7_75t_L g5510 ( 
.A(n_5189),
.B(n_4646),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_5035),
.Y(n_5511)
);

INVxp67_ASAP7_75t_SL g5512 ( 
.A(n_5140),
.Y(n_5512)
);

INVx3_ASAP7_75t_L g5513 ( 
.A(n_5213),
.Y(n_5513)
);

OR2x2_ASAP7_75t_L g5514 ( 
.A(n_5182),
.B(n_4920),
.Y(n_5514)
);

AND2x2_ASAP7_75t_L g5515 ( 
.A(n_5202),
.B(n_4855),
.Y(n_5515)
);

AND2x2_ASAP7_75t_L g5516 ( 
.A(n_5202),
.B(n_4855),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_5035),
.Y(n_5517)
);

INVx2_ASAP7_75t_L g5518 ( 
.A(n_4947),
.Y(n_5518)
);

OAI21xp5_ASAP7_75t_L g5519 ( 
.A1(n_4989),
.A2(n_4799),
.B(n_4755),
.Y(n_5519)
);

INVx2_ASAP7_75t_L g5520 ( 
.A(n_5120),
.Y(n_5520)
);

AND2x2_ASAP7_75t_L g5521 ( 
.A(n_5209),
.B(n_4855),
.Y(n_5521)
);

AND2x2_ASAP7_75t_L g5522 ( 
.A(n_5209),
.B(n_4855),
.Y(n_5522)
);

OR2x2_ASAP7_75t_L g5523 ( 
.A(n_5182),
.B(n_4920),
.Y(n_5523)
);

HB1xp67_ASAP7_75t_L g5524 ( 
.A(n_5179),
.Y(n_5524)
);

INVx2_ASAP7_75t_L g5525 ( 
.A(n_5120),
.Y(n_5525)
);

INVx2_ASAP7_75t_L g5526 ( 
.A(n_5120),
.Y(n_5526)
);

INVx2_ASAP7_75t_L g5527 ( 
.A(n_5134),
.Y(n_5527)
);

OR2x2_ASAP7_75t_L g5528 ( 
.A(n_5026),
.B(n_4926),
.Y(n_5528)
);

OR2x2_ASAP7_75t_L g5529 ( 
.A(n_4940),
.B(n_4945),
.Y(n_5529)
);

AND2x2_ASAP7_75t_L g5530 ( 
.A(n_5239),
.B(n_4855),
.Y(n_5530)
);

NAND2xp5_ASAP7_75t_L g5531 ( 
.A(n_5188),
.B(n_4457),
.Y(n_5531)
);

CKINVDCx5p33_ASAP7_75t_R g5532 ( 
.A(n_5137),
.Y(n_5532)
);

AND2x2_ASAP7_75t_L g5533 ( 
.A(n_5239),
.B(n_4855),
.Y(n_5533)
);

AND2x2_ASAP7_75t_L g5534 ( 
.A(n_5247),
.B(n_4914),
.Y(n_5534)
);

AND2x2_ASAP7_75t_L g5535 ( 
.A(n_5247),
.B(n_4914),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_5040),
.Y(n_5536)
);

AND2x2_ASAP7_75t_L g5537 ( 
.A(n_5264),
.B(n_4914),
.Y(n_5537)
);

BUFx2_ASAP7_75t_L g5538 ( 
.A(n_4942),
.Y(n_5538)
);

AND2x2_ASAP7_75t_L g5539 ( 
.A(n_5264),
.B(n_4914),
.Y(n_5539)
);

INVx1_ASAP7_75t_L g5540 ( 
.A(n_5040),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_5052),
.Y(n_5541)
);

HB1xp67_ASAP7_75t_L g5542 ( 
.A(n_5253),
.Y(n_5542)
);

INVx2_ASAP7_75t_L g5543 ( 
.A(n_5134),
.Y(n_5543)
);

INVx2_ASAP7_75t_L g5544 ( 
.A(n_5134),
.Y(n_5544)
);

INVx2_ASAP7_75t_L g5545 ( 
.A(n_5050),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5052),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_5056),
.Y(n_5547)
);

NAND2xp5_ASAP7_75t_L g5548 ( 
.A(n_5302),
.B(n_4963),
.Y(n_5548)
);

NOR2xp33_ASAP7_75t_L g5549 ( 
.A(n_5261),
.B(n_4754),
.Y(n_5549)
);

NAND2xp5_ASAP7_75t_L g5550 ( 
.A(n_4988),
.B(n_4457),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_5056),
.Y(n_5551)
);

NOR2xp33_ASAP7_75t_L g5552 ( 
.A(n_5246),
.B(n_4754),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5058),
.Y(n_5553)
);

AO221x2_ASAP7_75t_L g5554 ( 
.A1(n_5033),
.A2(n_4598),
.B1(n_4623),
.B2(n_4249),
.C(n_4087),
.Y(n_5554)
);

HB1xp67_ASAP7_75t_L g5555 ( 
.A(n_5262),
.Y(n_5555)
);

AND2x2_ASAP7_75t_L g5556 ( 
.A(n_5284),
.B(n_4914),
.Y(n_5556)
);

INVx2_ASAP7_75t_L g5557 ( 
.A(n_5050),
.Y(n_5557)
);

AND2x2_ASAP7_75t_L g5558 ( 
.A(n_5284),
.B(n_5285),
.Y(n_5558)
);

BUFx3_ASAP7_75t_L g5559 ( 
.A(n_5184),
.Y(n_5559)
);

AND2x2_ASAP7_75t_L g5560 ( 
.A(n_5285),
.B(n_4914),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_5058),
.Y(n_5561)
);

INVx2_ASAP7_75t_L g5562 ( 
.A(n_5050),
.Y(n_5562)
);

INVx2_ASAP7_75t_SL g5563 ( 
.A(n_5184),
.Y(n_5563)
);

AND2x2_ASAP7_75t_L g5564 ( 
.A(n_5291),
.B(n_4915),
.Y(n_5564)
);

AND2x2_ASAP7_75t_L g5565 ( 
.A(n_5291),
.B(n_4915),
.Y(n_5565)
);

INVx2_ASAP7_75t_L g5566 ( 
.A(n_5237),
.Y(n_5566)
);

HB1xp67_ASAP7_75t_L g5567 ( 
.A(n_4931),
.Y(n_5567)
);

INVx2_ASAP7_75t_L g5568 ( 
.A(n_5237),
.Y(n_5568)
);

AND2x2_ASAP7_75t_L g5569 ( 
.A(n_5323),
.B(n_4915),
.Y(n_5569)
);

AND2x4_ASAP7_75t_L g5570 ( 
.A(n_4987),
.B(n_4679),
.Y(n_5570)
);

INVx2_ASAP7_75t_L g5571 ( 
.A(n_5237),
.Y(n_5571)
);

OR2x2_ASAP7_75t_L g5572 ( 
.A(n_4940),
.B(n_4901),
.Y(n_5572)
);

AND2x2_ASAP7_75t_L g5573 ( 
.A(n_5323),
.B(n_4915),
.Y(n_5573)
);

OR2x2_ASAP7_75t_L g5574 ( 
.A(n_4945),
.B(n_4901),
.Y(n_5574)
);

INVx2_ASAP7_75t_L g5575 ( 
.A(n_5064),
.Y(n_5575)
);

AND2x2_ASAP7_75t_L g5576 ( 
.A(n_4996),
.B(n_4915),
.Y(n_5576)
);

OAI211xp5_ASAP7_75t_L g5577 ( 
.A1(n_5275),
.A2(n_4848),
.B(n_4915),
.C(n_4301),
.Y(n_5577)
);

INVxp67_ASAP7_75t_L g5578 ( 
.A(n_4988),
.Y(n_5578)
);

NAND2xp5_ASAP7_75t_L g5579 ( 
.A(n_5057),
.B(n_4468),
.Y(n_5579)
);

INVx2_ASAP7_75t_L g5580 ( 
.A(n_5064),
.Y(n_5580)
);

AND2x2_ASAP7_75t_L g5581 ( 
.A(n_4996),
.B(n_4739),
.Y(n_5581)
);

AND2x2_ASAP7_75t_L g5582 ( 
.A(n_5328),
.B(n_4434),
.Y(n_5582)
);

OR2x2_ASAP7_75t_L g5583 ( 
.A(n_5073),
.B(n_4905),
.Y(n_5583)
);

BUFx3_ASAP7_75t_L g5584 ( 
.A(n_5184),
.Y(n_5584)
);

AND2x2_ASAP7_75t_L g5585 ( 
.A(n_5328),
.B(n_4788),
.Y(n_5585)
);

HB1xp67_ASAP7_75t_L g5586 ( 
.A(n_4931),
.Y(n_5586)
);

INVx2_ASAP7_75t_L g5587 ( 
.A(n_5064),
.Y(n_5587)
);

INVx6_ASAP7_75t_L g5588 ( 
.A(n_4942),
.Y(n_5588)
);

OR2x2_ASAP7_75t_L g5589 ( 
.A(n_5073),
.B(n_4905),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_5061),
.Y(n_5590)
);

INVxp67_ASAP7_75t_SL g5591 ( 
.A(n_5184),
.Y(n_5591)
);

HB1xp67_ASAP7_75t_L g5592 ( 
.A(n_4932),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_5061),
.Y(n_5593)
);

INVx2_ASAP7_75t_L g5594 ( 
.A(n_5104),
.Y(n_5594)
);

NAND2xp5_ASAP7_75t_L g5595 ( 
.A(n_5057),
.B(n_4468),
.Y(n_5595)
);

OR2x2_ASAP7_75t_L g5596 ( 
.A(n_5293),
.B(n_4538),
.Y(n_5596)
);

AND2x2_ASAP7_75t_L g5597 ( 
.A(n_5341),
.B(n_4788),
.Y(n_5597)
);

NAND3xp33_ASAP7_75t_L g5598 ( 
.A(n_5047),
.B(n_4475),
.C(n_4814),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5104),
.Y(n_5599)
);

AND2x2_ASAP7_75t_L g5600 ( 
.A(n_5341),
.B(n_4501),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_5062),
.Y(n_5601)
);

AND2x2_ASAP7_75t_L g5602 ( 
.A(n_5345),
.B(n_4501),
.Y(n_5602)
);

INVx3_ASAP7_75t_L g5603 ( 
.A(n_5213),
.Y(n_5603)
);

HB1xp67_ASAP7_75t_L g5604 ( 
.A(n_4932),
.Y(n_5604)
);

AND2x2_ASAP7_75t_L g5605 ( 
.A(n_5345),
.B(n_4521),
.Y(n_5605)
);

NAND2xp5_ASAP7_75t_L g5606 ( 
.A(n_5095),
.B(n_4475),
.Y(n_5606)
);

BUFx2_ASAP7_75t_L g5607 ( 
.A(n_4942),
.Y(n_5607)
);

INVx2_ASAP7_75t_L g5608 ( 
.A(n_5104),
.Y(n_5608)
);

INVx1_ASAP7_75t_L g5609 ( 
.A(n_5062),
.Y(n_5609)
);

INVx2_ASAP7_75t_L g5610 ( 
.A(n_5263),
.Y(n_5610)
);

BUFx3_ASAP7_75t_L g5611 ( 
.A(n_5184),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_5071),
.Y(n_5612)
);

INVx2_ASAP7_75t_L g5613 ( 
.A(n_5263),
.Y(n_5613)
);

HB1xp67_ASAP7_75t_L g5614 ( 
.A(n_4943),
.Y(n_5614)
);

AND2x2_ASAP7_75t_L g5615 ( 
.A(n_4936),
.B(n_4521),
.Y(n_5615)
);

AND2x2_ASAP7_75t_L g5616 ( 
.A(n_4936),
.B(n_4528),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5071),
.Y(n_5617)
);

INVx2_ASAP7_75t_L g5618 ( 
.A(n_5263),
.Y(n_5618)
);

HB1xp67_ASAP7_75t_L g5619 ( 
.A(n_4943),
.Y(n_5619)
);

BUFx2_ASAP7_75t_L g5620 ( 
.A(n_4942),
.Y(n_5620)
);

OR2x2_ASAP7_75t_L g5621 ( 
.A(n_5293),
.B(n_4540),
.Y(n_5621)
);

NOR2xp33_ASAP7_75t_L g5622 ( 
.A(n_5246),
.B(n_4754),
.Y(n_5622)
);

INVx2_ASAP7_75t_L g5623 ( 
.A(n_5242),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5075),
.Y(n_5624)
);

AND2x2_ASAP7_75t_L g5625 ( 
.A(n_4936),
.B(n_4528),
.Y(n_5625)
);

INVx2_ASAP7_75t_L g5626 ( 
.A(n_5242),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5075),
.Y(n_5627)
);

INVx3_ASAP7_75t_L g5628 ( 
.A(n_5068),
.Y(n_5628)
);

AND2x2_ASAP7_75t_L g5629 ( 
.A(n_4936),
.B(n_4895),
.Y(n_5629)
);

INVx3_ASAP7_75t_SL g5630 ( 
.A(n_5266),
.Y(n_5630)
);

AND2x2_ASAP7_75t_L g5631 ( 
.A(n_4978),
.B(n_4895),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_5242),
.Y(n_5632)
);

OR2x6_ASAP7_75t_L g5633 ( 
.A(n_5335),
.B(n_4001),
.Y(n_5633)
);

INVx2_ASAP7_75t_SL g5634 ( 
.A(n_5266),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_5079),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5079),
.Y(n_5636)
);

INVx1_ASAP7_75t_L g5637 ( 
.A(n_5083),
.Y(n_5637)
);

INVx1_ASAP7_75t_L g5638 ( 
.A(n_5083),
.Y(n_5638)
);

INVx3_ASAP7_75t_L g5639 ( 
.A(n_5068),
.Y(n_5639)
);

AOI22xp33_ASAP7_75t_L g5640 ( 
.A1(n_5223),
.A2(n_4486),
.B1(n_4487),
.B2(n_4482),
.Y(n_5640)
);

INVx2_ASAP7_75t_L g5641 ( 
.A(n_5255),
.Y(n_5641)
);

AND2x2_ASAP7_75t_L g5642 ( 
.A(n_4978),
.B(n_4918),
.Y(n_5642)
);

INVx1_ASAP7_75t_L g5643 ( 
.A(n_5087),
.Y(n_5643)
);

INVx1_ASAP7_75t_L g5644 ( 
.A(n_5087),
.Y(n_5644)
);

NAND2xp5_ASAP7_75t_L g5645 ( 
.A(n_5095),
.B(n_4899),
.Y(n_5645)
);

INVxp67_ASAP7_75t_L g5646 ( 
.A(n_5154),
.Y(n_5646)
);

BUFx3_ASAP7_75t_L g5647 ( 
.A(n_5266),
.Y(n_5647)
);

INVx2_ASAP7_75t_L g5648 ( 
.A(n_5255),
.Y(n_5648)
);

AND2x4_ASAP7_75t_L g5649 ( 
.A(n_4987),
.B(n_4509),
.Y(n_5649)
);

OAI221xp5_ASAP7_75t_L g5650 ( 
.A1(n_4944),
.A2(n_4574),
.B1(n_4086),
.B2(n_4179),
.C(n_4176),
.Y(n_5650)
);

AND2x2_ASAP7_75t_L g5651 ( 
.A(n_4979),
.B(n_4918),
.Y(n_5651)
);

AND2x2_ASAP7_75t_L g5652 ( 
.A(n_4979),
.B(n_4743),
.Y(n_5652)
);

OR2x2_ASAP7_75t_L g5653 ( 
.A(n_5306),
.B(n_4899),
.Y(n_5653)
);

AND2x2_ASAP7_75t_L g5654 ( 
.A(n_5154),
.B(n_4743),
.Y(n_5654)
);

INVx2_ASAP7_75t_L g5655 ( 
.A(n_5255),
.Y(n_5655)
);

NAND2xp5_ASAP7_75t_L g5656 ( 
.A(n_5163),
.B(n_4902),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_5093),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_5163),
.B(n_4743),
.Y(n_5658)
);

BUFx2_ASAP7_75t_L g5659 ( 
.A(n_5266),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_5093),
.Y(n_5660)
);

AND2x2_ASAP7_75t_L g5661 ( 
.A(n_5167),
.B(n_4908),
.Y(n_5661)
);

HB1xp67_ASAP7_75t_L g5662 ( 
.A(n_4948),
.Y(n_5662)
);

AOI22xp33_ASAP7_75t_L g5663 ( 
.A1(n_5223),
.A2(n_5229),
.B1(n_5231),
.B2(n_4959),
.Y(n_5663)
);

AND2x2_ASAP7_75t_L g5664 ( 
.A(n_5167),
.B(n_4908),
.Y(n_5664)
);

AOI222xp33_ASAP7_75t_L g5665 ( 
.A1(n_5046),
.A2(n_4487),
.B1(n_4505),
.B2(n_4513),
.C1(n_4508),
.C2(n_4482),
.Y(n_5665)
);

INVx2_ASAP7_75t_L g5666 ( 
.A(n_5271),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_5099),
.Y(n_5667)
);

INVx1_ASAP7_75t_L g5668 ( 
.A(n_5099),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_5115),
.Y(n_5669)
);

INVx1_ASAP7_75t_L g5670 ( 
.A(n_5115),
.Y(n_5670)
);

INVx2_ASAP7_75t_L g5671 ( 
.A(n_5271),
.Y(n_5671)
);

INVx2_ASAP7_75t_L g5672 ( 
.A(n_5271),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_5118),
.Y(n_5673)
);

NOR2xp33_ASAP7_75t_L g5674 ( 
.A(n_5266),
.B(n_4795),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5118),
.Y(n_5675)
);

HB1xp67_ASAP7_75t_L g5676 ( 
.A(n_4948),
.Y(n_5676)
);

AND2x2_ASAP7_75t_L g5677 ( 
.A(n_5171),
.B(n_4908),
.Y(n_5677)
);

NAND2xp33_ASAP7_75t_R g5678 ( 
.A(n_5171),
.B(n_4813),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_5122),
.Y(n_5679)
);

BUFx2_ASAP7_75t_L g5680 ( 
.A(n_5199),
.Y(n_5680)
);

INVx2_ASAP7_75t_L g5681 ( 
.A(n_4952),
.Y(n_5681)
);

INVx1_ASAP7_75t_SL g5682 ( 
.A(n_5141),
.Y(n_5682)
);

INVx2_ASAP7_75t_L g5683 ( 
.A(n_4952),
.Y(n_5683)
);

INVx2_ASAP7_75t_L g5684 ( 
.A(n_4952),
.Y(n_5684)
);

INVx3_ASAP7_75t_L g5685 ( 
.A(n_5068),
.Y(n_5685)
);

BUFx2_ASAP7_75t_L g5686 ( 
.A(n_5199),
.Y(n_5686)
);

INVx2_ASAP7_75t_L g5687 ( 
.A(n_4968),
.Y(n_5687)
);

AO21x2_ASAP7_75t_L g5688 ( 
.A1(n_4959),
.A2(n_4804),
.B(n_4800),
.Y(n_5688)
);

INVx3_ASAP7_75t_L g5689 ( 
.A(n_5068),
.Y(n_5689)
);

INVx2_ASAP7_75t_L g5690 ( 
.A(n_4968),
.Y(n_5690)
);

AND2x2_ASAP7_75t_L g5691 ( 
.A(n_4971),
.B(n_4419),
.Y(n_5691)
);

AND2x2_ASAP7_75t_L g5692 ( 
.A(n_4971),
.B(n_4419),
.Y(n_5692)
);

OR2x2_ASAP7_75t_L g5693 ( 
.A(n_5306),
.B(n_4540),
.Y(n_5693)
);

NAND2xp5_ASAP7_75t_L g5694 ( 
.A(n_4950),
.B(n_4543),
.Y(n_5694)
);

INVxp67_ASAP7_75t_SL g5695 ( 
.A(n_5307),
.Y(n_5695)
);

INVxp67_ASAP7_75t_SL g5696 ( 
.A(n_5339),
.Y(n_5696)
);

INVx2_ASAP7_75t_L g5697 ( 
.A(n_4968),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_5122),
.Y(n_5698)
);

INVx1_ASAP7_75t_L g5699 ( 
.A(n_5123),
.Y(n_5699)
);

BUFx3_ASAP7_75t_L g5700 ( 
.A(n_5155),
.Y(n_5700)
);

INVxp67_ASAP7_75t_SL g5701 ( 
.A(n_5663),
.Y(n_5701)
);

AND2x2_ASAP7_75t_L g5702 ( 
.A(n_5464),
.B(n_5211),
.Y(n_5702)
);

AND2x2_ASAP7_75t_L g5703 ( 
.A(n_5464),
.B(n_5211),
.Y(n_5703)
);

AND2x2_ASAP7_75t_L g5704 ( 
.A(n_5582),
.B(n_5211),
.Y(n_5704)
);

AND2x2_ASAP7_75t_L g5705 ( 
.A(n_5582),
.B(n_5211),
.Y(n_5705)
);

NAND2xp5_ASAP7_75t_L g5706 ( 
.A(n_5421),
.B(n_5339),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5529),
.Y(n_5707)
);

AND2x4_ASAP7_75t_L g5708 ( 
.A(n_5419),
.B(n_4999),
.Y(n_5708)
);

OR2x2_ASAP7_75t_L g5709 ( 
.A(n_5365),
.B(n_5088),
.Y(n_5709)
);

AND2x2_ASAP7_75t_L g5710 ( 
.A(n_5558),
.B(n_4999),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_5491),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_5503),
.Y(n_5712)
);

AND2x2_ASAP7_75t_L g5713 ( 
.A(n_5558),
.B(n_5038),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_5363),
.Y(n_5714)
);

BUFx3_ASAP7_75t_L g5715 ( 
.A(n_5410),
.Y(n_5715)
);

INVx2_ASAP7_75t_L g5716 ( 
.A(n_5688),
.Y(n_5716)
);

AND2x2_ASAP7_75t_L g5717 ( 
.A(n_5461),
.B(n_5470),
.Y(n_5717)
);

INVx1_ASAP7_75t_L g5718 ( 
.A(n_5367),
.Y(n_5718)
);

INVx2_ASAP7_75t_L g5719 ( 
.A(n_5688),
.Y(n_5719)
);

AND2x2_ASAP7_75t_L g5720 ( 
.A(n_5461),
.B(n_5038),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_5369),
.Y(n_5721)
);

INVx1_ASAP7_75t_SL g5722 ( 
.A(n_5410),
.Y(n_5722)
);

OR2x2_ASAP7_75t_L g5723 ( 
.A(n_5352),
.B(n_5088),
.Y(n_5723)
);

HB1xp67_ASAP7_75t_L g5724 ( 
.A(n_5628),
.Y(n_5724)
);

NAND2xp5_ASAP7_75t_L g5725 ( 
.A(n_5682),
.B(n_5045),
.Y(n_5725)
);

AND2x4_ASAP7_75t_L g5726 ( 
.A(n_5448),
.B(n_5408),
.Y(n_5726)
);

OR2x2_ASAP7_75t_L g5727 ( 
.A(n_5548),
.B(n_5101),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_5371),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_5376),
.Y(n_5729)
);

INVx2_ASAP7_75t_L g5730 ( 
.A(n_5688),
.Y(n_5730)
);

AND2x2_ASAP7_75t_L g5731 ( 
.A(n_5470),
.B(n_5045),
.Y(n_5731)
);

BUFx6f_ASAP7_75t_L g5732 ( 
.A(n_5350),
.Y(n_5732)
);

INVx3_ASAP7_75t_L g5733 ( 
.A(n_5455),
.Y(n_5733)
);

AND2x2_ASAP7_75t_L g5734 ( 
.A(n_5473),
.B(n_5067),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_5378),
.Y(n_5735)
);

NAND2x1_ASAP7_75t_L g5736 ( 
.A(n_5649),
.B(n_5196),
.Y(n_5736)
);

INVx1_ASAP7_75t_L g5737 ( 
.A(n_5392),
.Y(n_5737)
);

OR2x2_ASAP7_75t_L g5738 ( 
.A(n_5364),
.B(n_5101),
.Y(n_5738)
);

NAND2xp5_ASAP7_75t_L g5739 ( 
.A(n_5680),
.B(n_5067),
.Y(n_5739)
);

HB1xp67_ASAP7_75t_L g5740 ( 
.A(n_5628),
.Y(n_5740)
);

BUFx3_ASAP7_75t_L g5741 ( 
.A(n_5588),
.Y(n_5741)
);

AND2x2_ASAP7_75t_L g5742 ( 
.A(n_5473),
.B(n_5076),
.Y(n_5742)
);

BUFx2_ASAP7_75t_L g5743 ( 
.A(n_5538),
.Y(n_5743)
);

AND2x4_ASAP7_75t_L g5744 ( 
.A(n_5408),
.B(n_5076),
.Y(n_5744)
);

AND2x2_ASAP7_75t_L g5745 ( 
.A(n_5400),
.B(n_5221),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5393),
.Y(n_5746)
);

NAND2xp5_ASAP7_75t_L g5747 ( 
.A(n_5686),
.B(n_5221),
.Y(n_5747)
);

INVx2_ASAP7_75t_L g5748 ( 
.A(n_5628),
.Y(n_5748)
);

INVx2_ASAP7_75t_L g5749 ( 
.A(n_5639),
.Y(n_5749)
);

INVx2_ASAP7_75t_L g5750 ( 
.A(n_5639),
.Y(n_5750)
);

AND2x2_ASAP7_75t_L g5751 ( 
.A(n_5400),
.B(n_5245),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_5406),
.Y(n_5752)
);

INVx2_ASAP7_75t_L g5753 ( 
.A(n_5639),
.Y(n_5753)
);

NAND2xp5_ASAP7_75t_L g5754 ( 
.A(n_5578),
.B(n_5245),
.Y(n_5754)
);

AND2x4_ASAP7_75t_L g5755 ( 
.A(n_5408),
.B(n_5072),
.Y(n_5755)
);

AND2x2_ASAP7_75t_L g5756 ( 
.A(n_5402),
.B(n_4483),
.Y(n_5756)
);

OR2x6_ASAP7_75t_L g5757 ( 
.A(n_5588),
.B(n_4483),
.Y(n_5757)
);

BUFx3_ASAP7_75t_L g5758 ( 
.A(n_5588),
.Y(n_5758)
);

OR2x2_ASAP7_75t_L g5759 ( 
.A(n_5433),
.B(n_5112),
.Y(n_5759)
);

OR2x2_ASAP7_75t_L g5760 ( 
.A(n_5488),
.B(n_5112),
.Y(n_5760)
);

OR2x2_ASAP7_75t_L g5761 ( 
.A(n_5509),
.B(n_5065),
.Y(n_5761)
);

BUFx6f_ASAP7_75t_L g5762 ( 
.A(n_5350),
.Y(n_5762)
);

INVx2_ASAP7_75t_SL g5763 ( 
.A(n_5408),
.Y(n_5763)
);

NAND2xp5_ASAP7_75t_L g5764 ( 
.A(n_5646),
.B(n_4950),
.Y(n_5764)
);

AOI22xp33_ASAP7_75t_L g5765 ( 
.A1(n_5355),
.A2(n_5229),
.B1(n_5231),
.B2(n_4959),
.Y(n_5765)
);

INVx3_ASAP7_75t_L g5766 ( 
.A(n_5685),
.Y(n_5766)
);

BUFx2_ASAP7_75t_L g5767 ( 
.A(n_5607),
.Y(n_5767)
);

NOR2x1_ASAP7_75t_SL g5768 ( 
.A(n_5633),
.B(n_4995),
.Y(n_5768)
);

AND2x2_ASAP7_75t_L g5769 ( 
.A(n_5402),
.B(n_4994),
.Y(n_5769)
);

AND2x2_ASAP7_75t_L g5770 ( 
.A(n_5383),
.B(n_4795),
.Y(n_5770)
);

BUFx2_ASAP7_75t_L g5771 ( 
.A(n_5620),
.Y(n_5771)
);

AND2x4_ASAP7_75t_L g5772 ( 
.A(n_5408),
.B(n_5196),
.Y(n_5772)
);

AND2x2_ASAP7_75t_L g5773 ( 
.A(n_5383),
.B(n_4795),
.Y(n_5773)
);

OR2x2_ASAP7_75t_L g5774 ( 
.A(n_5524),
.B(n_5065),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_5407),
.Y(n_5775)
);

NOR2x1p5_ASAP7_75t_L g5776 ( 
.A(n_5532),
.B(n_4001),
.Y(n_5776)
);

HB1xp67_ASAP7_75t_L g5777 ( 
.A(n_5685),
.Y(n_5777)
);

AND2x2_ASAP7_75t_L g5778 ( 
.A(n_5404),
.B(n_4973),
.Y(n_5778)
);

INVx2_ASAP7_75t_L g5779 ( 
.A(n_5685),
.Y(n_5779)
);

INVx1_ASAP7_75t_L g5780 ( 
.A(n_5413),
.Y(n_5780)
);

INVx2_ASAP7_75t_L g5781 ( 
.A(n_5689),
.Y(n_5781)
);

AND2x2_ASAP7_75t_L g5782 ( 
.A(n_5404),
.B(n_4973),
.Y(n_5782)
);

AND2x2_ASAP7_75t_L g5783 ( 
.A(n_5405),
.B(n_5007),
.Y(n_5783)
);

BUFx3_ASAP7_75t_L g5784 ( 
.A(n_5532),
.Y(n_5784)
);

AND2x2_ASAP7_75t_L g5785 ( 
.A(n_5405),
.B(n_5007),
.Y(n_5785)
);

NAND2xp5_ASAP7_75t_L g5786 ( 
.A(n_5436),
.B(n_4951),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_5424),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_5427),
.Y(n_5788)
);

INVx1_ASAP7_75t_L g5789 ( 
.A(n_5435),
.Y(n_5789)
);

AND2x2_ASAP7_75t_L g5790 ( 
.A(n_5414),
.B(n_5023),
.Y(n_5790)
);

INVx3_ASAP7_75t_L g5791 ( 
.A(n_5689),
.Y(n_5791)
);

AOI22xp33_ASAP7_75t_L g5792 ( 
.A1(n_5355),
.A2(n_5231),
.B1(n_5229),
.B2(n_5041),
.Y(n_5792)
);

INVx2_ASAP7_75t_SL g5793 ( 
.A(n_5451),
.Y(n_5793)
);

BUFx2_ASAP7_75t_L g5794 ( 
.A(n_5700),
.Y(n_5794)
);

BUFx2_ASAP7_75t_L g5795 ( 
.A(n_5700),
.Y(n_5795)
);

INVx2_ASAP7_75t_L g5796 ( 
.A(n_5689),
.Y(n_5796)
);

INVx1_ASAP7_75t_L g5797 ( 
.A(n_5440),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5441),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5445),
.Y(n_5799)
);

OR2x2_ASAP7_75t_L g5800 ( 
.A(n_5354),
.B(n_5138),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5387),
.Y(n_5801)
);

INVxp67_ASAP7_75t_SL g5802 ( 
.A(n_5663),
.Y(n_5802)
);

HB1xp67_ASAP7_75t_L g5803 ( 
.A(n_5361),
.Y(n_5803)
);

AND2x2_ASAP7_75t_L g5804 ( 
.A(n_5414),
.B(n_5023),
.Y(n_5804)
);

AND2x4_ASAP7_75t_L g5805 ( 
.A(n_5465),
.B(n_5196),
.Y(n_5805)
);

INVx2_ASAP7_75t_L g5806 ( 
.A(n_5387),
.Y(n_5806)
);

INVx4_ASAP7_75t_L g5807 ( 
.A(n_5350),
.Y(n_5807)
);

INVx4_ASAP7_75t_L g5808 ( 
.A(n_5350),
.Y(n_5808)
);

AND2x4_ASAP7_75t_L g5809 ( 
.A(n_5465),
.B(n_5222),
.Y(n_5809)
);

INVx2_ASAP7_75t_L g5810 ( 
.A(n_5388),
.Y(n_5810)
);

INVx2_ASAP7_75t_L g5811 ( 
.A(n_5388),
.Y(n_5811)
);

INVx2_ASAP7_75t_L g5812 ( 
.A(n_5395),
.Y(n_5812)
);

AND2x2_ASAP7_75t_L g5813 ( 
.A(n_5416),
.B(n_5037),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_5446),
.Y(n_5814)
);

AND2x2_ASAP7_75t_L g5815 ( 
.A(n_5416),
.B(n_5037),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_5449),
.Y(n_5816)
);

HB1xp67_ASAP7_75t_L g5817 ( 
.A(n_5409),
.Y(n_5817)
);

INVx2_ASAP7_75t_L g5818 ( 
.A(n_5395),
.Y(n_5818)
);

INVx2_ASAP7_75t_L g5819 ( 
.A(n_5399),
.Y(n_5819)
);

AND2x2_ASAP7_75t_L g5820 ( 
.A(n_5585),
.B(n_4974),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_5450),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5454),
.Y(n_5822)
);

INVx1_ASAP7_75t_L g5823 ( 
.A(n_5462),
.Y(n_5823)
);

INVx2_ASAP7_75t_L g5824 ( 
.A(n_5399),
.Y(n_5824)
);

INVx4_ASAP7_75t_L g5825 ( 
.A(n_5386),
.Y(n_5825)
);

INVx1_ASAP7_75t_L g5826 ( 
.A(n_5469),
.Y(n_5826)
);

NOR2xp33_ASAP7_75t_SL g5827 ( 
.A(n_5442),
.B(n_5172),
.Y(n_5827)
);

INVx2_ASAP7_75t_L g5828 ( 
.A(n_5401),
.Y(n_5828)
);

AND2x2_ASAP7_75t_L g5829 ( 
.A(n_5585),
.B(n_4974),
.Y(n_5829)
);

INVx2_ASAP7_75t_L g5830 ( 
.A(n_5401),
.Y(n_5830)
);

OR2x2_ASAP7_75t_L g5831 ( 
.A(n_5528),
.B(n_5138),
.Y(n_5831)
);

INVx2_ASAP7_75t_L g5832 ( 
.A(n_5412),
.Y(n_5832)
);

INVx2_ASAP7_75t_L g5833 ( 
.A(n_5412),
.Y(n_5833)
);

AND2x4_ASAP7_75t_L g5834 ( 
.A(n_5465),
.B(n_5486),
.Y(n_5834)
);

NAND2xp5_ASAP7_75t_L g5835 ( 
.A(n_5453),
.B(n_4951),
.Y(n_5835)
);

INVx2_ASAP7_75t_L g5836 ( 
.A(n_5520),
.Y(n_5836)
);

AND2x2_ASAP7_75t_L g5837 ( 
.A(n_5597),
.B(n_4975),
.Y(n_5837)
);

NAND2xp5_ASAP7_75t_L g5838 ( 
.A(n_5696),
.B(n_4960),
.Y(n_5838)
);

INVx3_ASAP7_75t_L g5839 ( 
.A(n_5507),
.Y(n_5839)
);

AOI22xp5_ASAP7_75t_L g5840 ( 
.A1(n_5394),
.A2(n_5319),
.B1(n_5216),
.B2(n_5314),
.Y(n_5840)
);

AOI22xp5_ASAP7_75t_L g5841 ( 
.A1(n_5370),
.A2(n_5319),
.B1(n_5157),
.B2(n_5041),
.Y(n_5841)
);

INVx3_ASAP7_75t_SL g5842 ( 
.A(n_5474),
.Y(n_5842)
);

AND2x2_ASAP7_75t_L g5843 ( 
.A(n_5597),
.B(n_4975),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5471),
.Y(n_5844)
);

AND2x2_ASAP7_75t_L g5845 ( 
.A(n_5380),
.B(n_5039),
.Y(n_5845)
);

AND2x2_ASAP7_75t_L g5846 ( 
.A(n_5380),
.B(n_5039),
.Y(n_5846)
);

AND2x4_ASAP7_75t_L g5847 ( 
.A(n_5486),
.B(n_5222),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_5479),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5482),
.Y(n_5849)
);

INVx3_ASAP7_75t_L g5850 ( 
.A(n_5472),
.Y(n_5850)
);

OR2x2_ASAP7_75t_L g5851 ( 
.A(n_5377),
.B(n_5078),
.Y(n_5851)
);

INVx2_ASAP7_75t_L g5852 ( 
.A(n_5520),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_5497),
.Y(n_5853)
);

INVx1_ASAP7_75t_L g5854 ( 
.A(n_5499),
.Y(n_5854)
);

INVx5_ASAP7_75t_L g5855 ( 
.A(n_5396),
.Y(n_5855)
);

NAND2xp5_ASAP7_75t_L g5856 ( 
.A(n_5415),
.B(n_4960),
.Y(n_5856)
);

INVx2_ASAP7_75t_L g5857 ( 
.A(n_5525),
.Y(n_5857)
);

BUFx6f_ASAP7_75t_L g5858 ( 
.A(n_5451),
.Y(n_5858)
);

NAND2xp5_ASAP7_75t_L g5859 ( 
.A(n_5481),
.B(n_4964),
.Y(n_5859)
);

HB1xp67_ASAP7_75t_L g5860 ( 
.A(n_5382),
.Y(n_5860)
);

INVx2_ASAP7_75t_SL g5861 ( 
.A(n_5451),
.Y(n_5861)
);

INVx1_ASAP7_75t_L g5862 ( 
.A(n_5501),
.Y(n_5862)
);

NAND2xp5_ASAP7_75t_L g5863 ( 
.A(n_5542),
.B(n_4964),
.Y(n_5863)
);

AOI22xp33_ASAP7_75t_L g5864 ( 
.A1(n_5370),
.A2(n_5054),
.B1(n_5055),
.B2(n_5032),
.Y(n_5864)
);

INVx2_ASAP7_75t_L g5865 ( 
.A(n_5525),
.Y(n_5865)
);

INVx2_ASAP7_75t_L g5866 ( 
.A(n_5526),
.Y(n_5866)
);

NAND2xp5_ASAP7_75t_L g5867 ( 
.A(n_5555),
.B(n_4967),
.Y(n_5867)
);

AND2x4_ASAP7_75t_L g5868 ( 
.A(n_5486),
.B(n_5222),
.Y(n_5868)
);

INVx2_ASAP7_75t_L g5869 ( 
.A(n_5526),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_5506),
.Y(n_5870)
);

INVx2_ASAP7_75t_L g5871 ( 
.A(n_5527),
.Y(n_5871)
);

AND2x2_ASAP7_75t_L g5872 ( 
.A(n_5397),
.B(n_5044),
.Y(n_5872)
);

NAND2xp5_ASAP7_75t_L g5873 ( 
.A(n_5379),
.B(n_4967),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5511),
.Y(n_5874)
);

AND2x4_ASAP7_75t_L g5875 ( 
.A(n_5559),
.B(n_5222),
.Y(n_5875)
);

HB1xp67_ASAP7_75t_L g5876 ( 
.A(n_5567),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_5517),
.Y(n_5877)
);

AND2x2_ASAP7_75t_L g5878 ( 
.A(n_5397),
.B(n_5044),
.Y(n_5878)
);

INVx2_ASAP7_75t_L g5879 ( 
.A(n_5527),
.Y(n_5879)
);

CKINVDCx5p33_ASAP7_75t_R g5880 ( 
.A(n_5373),
.Y(n_5880)
);

HB1xp67_ASAP7_75t_L g5881 ( 
.A(n_5586),
.Y(n_5881)
);

INVx2_ASAP7_75t_L g5882 ( 
.A(n_5543),
.Y(n_5882)
);

AND2x2_ASAP7_75t_L g5883 ( 
.A(n_5463),
.B(n_5084),
.Y(n_5883)
);

AND2x2_ASAP7_75t_L g5884 ( 
.A(n_5500),
.B(n_5084),
.Y(n_5884)
);

AND2x2_ASAP7_75t_L g5885 ( 
.A(n_5508),
.B(n_5092),
.Y(n_5885)
);

OR2x2_ASAP7_75t_L g5886 ( 
.A(n_5426),
.B(n_5049),
.Y(n_5886)
);

HB1xp67_ASAP7_75t_L g5887 ( 
.A(n_5592),
.Y(n_5887)
);

INVx2_ASAP7_75t_L g5888 ( 
.A(n_5543),
.Y(n_5888)
);

NAND2xp5_ASAP7_75t_L g5889 ( 
.A(n_5512),
.B(n_5181),
.Y(n_5889)
);

CKINVDCx5p33_ASAP7_75t_R g5890 ( 
.A(n_5390),
.Y(n_5890)
);

INVx3_ASAP7_75t_L g5891 ( 
.A(n_5472),
.Y(n_5891)
);

AND2x2_ASAP7_75t_L g5892 ( 
.A(n_5649),
.B(n_5092),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5536),
.Y(n_5893)
);

INVx1_ASAP7_75t_L g5894 ( 
.A(n_5540),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5541),
.Y(n_5895)
);

INVx3_ASAP7_75t_L g5896 ( 
.A(n_5451),
.Y(n_5896)
);

AND2x2_ASAP7_75t_L g5897 ( 
.A(n_5649),
.B(n_5098),
.Y(n_5897)
);

INVx1_ASAP7_75t_L g5898 ( 
.A(n_5546),
.Y(n_5898)
);

INVx1_ASAP7_75t_L g5899 ( 
.A(n_5547),
.Y(n_5899)
);

NAND2xp5_ASAP7_75t_L g5900 ( 
.A(n_5570),
.B(n_5114),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_5551),
.Y(n_5901)
);

HB1xp67_ASAP7_75t_L g5902 ( 
.A(n_5604),
.Y(n_5902)
);

INVx4_ASAP7_75t_L g5903 ( 
.A(n_5474),
.Y(n_5903)
);

BUFx3_ASAP7_75t_L g5904 ( 
.A(n_5442),
.Y(n_5904)
);

INVx2_ASAP7_75t_SL g5905 ( 
.A(n_5559),
.Y(n_5905)
);

AND2x2_ASAP7_75t_L g5906 ( 
.A(n_5348),
.B(n_5098),
.Y(n_5906)
);

AND2x2_ASAP7_75t_L g5907 ( 
.A(n_5348),
.B(n_5100),
.Y(n_5907)
);

AND2x2_ASAP7_75t_L g5908 ( 
.A(n_5459),
.B(n_5460),
.Y(n_5908)
);

INVx1_ASAP7_75t_L g5909 ( 
.A(n_5553),
.Y(n_5909)
);

NAND2xp5_ASAP7_75t_L g5910 ( 
.A(n_5570),
.B(n_5315),
.Y(n_5910)
);

AND2x2_ASAP7_75t_L g5911 ( 
.A(n_5459),
.B(n_5460),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5561),
.Y(n_5912)
);

INVx2_ASAP7_75t_L g5913 ( 
.A(n_5544),
.Y(n_5913)
);

BUFx2_ASAP7_75t_L g5914 ( 
.A(n_5584),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5590),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5593),
.Y(n_5916)
);

BUFx2_ASAP7_75t_L g5917 ( 
.A(n_5584),
.Y(n_5917)
);

AND2x2_ASAP7_75t_L g5918 ( 
.A(n_5630),
.B(n_5100),
.Y(n_5918)
);

INVx1_ASAP7_75t_L g5919 ( 
.A(n_5601),
.Y(n_5919)
);

HB1xp67_ASAP7_75t_L g5920 ( 
.A(n_5614),
.Y(n_5920)
);

AND2x2_ASAP7_75t_L g5921 ( 
.A(n_5630),
.B(n_5102),
.Y(n_5921)
);

INVx1_ASAP7_75t_L g5922 ( 
.A(n_5609),
.Y(n_5922)
);

AOI21xp5_ASAP7_75t_SL g5923 ( 
.A1(n_5554),
.A2(n_5015),
.B(n_4995),
.Y(n_5923)
);

AND2x2_ASAP7_75t_L g5924 ( 
.A(n_5549),
.B(n_5102),
.Y(n_5924)
);

NAND2x1p5_ASAP7_75t_L g5925 ( 
.A(n_5611),
.B(n_4221),
.Y(n_5925)
);

INVx2_ASAP7_75t_L g5926 ( 
.A(n_5544),
.Y(n_5926)
);

OR2x2_ASAP7_75t_L g5927 ( 
.A(n_5444),
.B(n_5053),
.Y(n_5927)
);

AND2x4_ASAP7_75t_L g5928 ( 
.A(n_5611),
.B(n_5308),
.Y(n_5928)
);

INVx2_ASAP7_75t_L g5929 ( 
.A(n_5438),
.Y(n_5929)
);

OR2x2_ASAP7_75t_L g5930 ( 
.A(n_5487),
.B(n_5053),
.Y(n_5930)
);

INVx1_ASAP7_75t_L g5931 ( 
.A(n_5612),
.Y(n_5931)
);

INVx1_ASAP7_75t_L g5932 ( 
.A(n_5617),
.Y(n_5932)
);

OR2x2_ASAP7_75t_L g5933 ( 
.A(n_5494),
.B(n_5200),
.Y(n_5933)
);

AND2x2_ASAP7_75t_L g5934 ( 
.A(n_5549),
.B(n_5051),
.Y(n_5934)
);

INVxp67_ASAP7_75t_SL g5935 ( 
.A(n_5477),
.Y(n_5935)
);

NAND2xp5_ASAP7_75t_L g5936 ( 
.A(n_5570),
.B(n_5318),
.Y(n_5936)
);

AND2x2_ASAP7_75t_L g5937 ( 
.A(n_5398),
.B(n_5051),
.Y(n_5937)
);

BUFx2_ASAP7_75t_L g5938 ( 
.A(n_5647),
.Y(n_5938)
);

INVx2_ASAP7_75t_L g5939 ( 
.A(n_5438),
.Y(n_5939)
);

OR2x2_ASAP7_75t_L g5940 ( 
.A(n_5572),
.B(n_5574),
.Y(n_5940)
);

INVx2_ASAP7_75t_L g5941 ( 
.A(n_5447),
.Y(n_5941)
);

INVx2_ASAP7_75t_L g5942 ( 
.A(n_5447),
.Y(n_5942)
);

NOR2xp33_ASAP7_75t_L g5943 ( 
.A(n_5457),
.B(n_4622),
.Y(n_5943)
);

INVx2_ASAP7_75t_L g5944 ( 
.A(n_5466),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5624),
.Y(n_5945)
);

NOR2xp67_ASAP7_75t_L g5946 ( 
.A(n_5374),
.B(n_5308),
.Y(n_5946)
);

INVx1_ASAP7_75t_L g5947 ( 
.A(n_5627),
.Y(n_5947)
);

AND2x2_ASAP7_75t_L g5948 ( 
.A(n_5398),
.B(n_5366),
.Y(n_5948)
);

AND2x2_ASAP7_75t_L g5949 ( 
.A(n_5366),
.B(n_5059),
.Y(n_5949)
);

INVx2_ASAP7_75t_L g5950 ( 
.A(n_5466),
.Y(n_5950)
);

NAND2xp5_ASAP7_75t_SL g5951 ( 
.A(n_5476),
.B(n_5340),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5635),
.Y(n_5952)
);

NAND2xp5_ASAP7_75t_L g5953 ( 
.A(n_5591),
.B(n_5329),
.Y(n_5953)
);

AND2x2_ASAP7_75t_L g5954 ( 
.A(n_5428),
.B(n_5059),
.Y(n_5954)
);

BUFx2_ASAP7_75t_L g5955 ( 
.A(n_5647),
.Y(n_5955)
);

INVx2_ASAP7_75t_L g5956 ( 
.A(n_5358),
.Y(n_5956)
);

AND2x2_ASAP7_75t_L g5957 ( 
.A(n_5428),
.B(n_5074),
.Y(n_5957)
);

INVx1_ASAP7_75t_L g5958 ( 
.A(n_5636),
.Y(n_5958)
);

INVx1_ASAP7_75t_L g5959 ( 
.A(n_5637),
.Y(n_5959)
);

INVx1_ASAP7_75t_L g5960 ( 
.A(n_5638),
.Y(n_5960)
);

INVxp67_ASAP7_75t_L g5961 ( 
.A(n_5390),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5643),
.Y(n_5962)
);

AND2x4_ASAP7_75t_L g5963 ( 
.A(n_5374),
.B(n_5308),
.Y(n_5963)
);

OR2x2_ASAP7_75t_L g5964 ( 
.A(n_5391),
.B(n_5217),
.Y(n_5964)
);

BUFx3_ASAP7_75t_L g5965 ( 
.A(n_5457),
.Y(n_5965)
);

INVx1_ASAP7_75t_L g5966 ( 
.A(n_5644),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_5657),
.Y(n_5967)
);

INVx3_ASAP7_75t_L g5968 ( 
.A(n_5430),
.Y(n_5968)
);

HB1xp67_ASAP7_75t_L g5969 ( 
.A(n_5619),
.Y(n_5969)
);

INVx2_ASAP7_75t_L g5970 ( 
.A(n_5358),
.Y(n_5970)
);

INVx2_ASAP7_75t_L g5971 ( 
.A(n_5372),
.Y(n_5971)
);

BUFx2_ASAP7_75t_L g5972 ( 
.A(n_5695),
.Y(n_5972)
);

NAND2xp5_ASAP7_75t_L g5973 ( 
.A(n_5662),
.B(n_5344),
.Y(n_5973)
);

NAND2xp5_ASAP7_75t_L g5974 ( 
.A(n_5676),
.B(n_5123),
.Y(n_5974)
);

NAND2xp5_ASAP7_75t_L g5975 ( 
.A(n_5452),
.B(n_5126),
.Y(n_5975)
);

NOR2xp33_ASAP7_75t_L g5976 ( 
.A(n_5674),
.B(n_4580),
.Y(n_5976)
);

INVx2_ASAP7_75t_SL g5977 ( 
.A(n_5381),
.Y(n_5977)
);

AND2x2_ASAP7_75t_L g5978 ( 
.A(n_5654),
.B(n_4995),
.Y(n_5978)
);

INVx2_ASAP7_75t_L g5979 ( 
.A(n_5372),
.Y(n_5979)
);

INVx2_ASAP7_75t_L g5980 ( 
.A(n_5385),
.Y(n_5980)
);

INVx1_ASAP7_75t_L g5981 ( 
.A(n_5660),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_5667),
.Y(n_5982)
);

INVx2_ASAP7_75t_L g5983 ( 
.A(n_5385),
.Y(n_5983)
);

BUFx3_ASAP7_75t_L g5984 ( 
.A(n_5674),
.Y(n_5984)
);

CKINVDCx5p33_ASAP7_75t_R g5985 ( 
.A(n_5477),
.Y(n_5985)
);

OR2x2_ASAP7_75t_L g5986 ( 
.A(n_5403),
.B(n_5230),
.Y(n_5986)
);

BUFx3_ASAP7_75t_L g5987 ( 
.A(n_5552),
.Y(n_5987)
);

BUFx3_ASAP7_75t_L g5988 ( 
.A(n_5552),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5545),
.Y(n_5989)
);

HB1xp67_ASAP7_75t_L g5990 ( 
.A(n_5468),
.Y(n_5990)
);

INVx1_ASAP7_75t_L g5991 ( 
.A(n_5668),
.Y(n_5991)
);

INVxp67_ASAP7_75t_SL g5992 ( 
.A(n_5678),
.Y(n_5992)
);

INVx1_ASAP7_75t_L g5993 ( 
.A(n_5669),
.Y(n_5993)
);

INVx2_ASAP7_75t_L g5994 ( 
.A(n_5545),
.Y(n_5994)
);

HB1xp67_ASAP7_75t_L g5995 ( 
.A(n_5468),
.Y(n_5995)
);

OR2x6_ASAP7_75t_L g5996 ( 
.A(n_5633),
.B(n_5335),
.Y(n_5996)
);

HB1xp67_ASAP7_75t_L g5997 ( 
.A(n_5475),
.Y(n_5997)
);

INVx1_ASAP7_75t_L g5998 ( 
.A(n_5670),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_5673),
.Y(n_5999)
);

INVx2_ASAP7_75t_L g6000 ( 
.A(n_5557),
.Y(n_6000)
);

INVx4_ASAP7_75t_L g6001 ( 
.A(n_5474),
.Y(n_6001)
);

AND2x4_ASAP7_75t_L g6002 ( 
.A(n_5452),
.B(n_5308),
.Y(n_6002)
);

INVxp67_ASAP7_75t_SL g6003 ( 
.A(n_5678),
.Y(n_6003)
);

BUFx2_ASAP7_75t_L g6004 ( 
.A(n_5659),
.Y(n_6004)
);

INVx1_ASAP7_75t_L g6005 ( 
.A(n_5675),
.Y(n_6005)
);

BUFx3_ASAP7_75t_L g6006 ( 
.A(n_5622),
.Y(n_6006)
);

AND2x4_ASAP7_75t_L g6007 ( 
.A(n_5563),
.B(n_4995),
.Y(n_6007)
);

INVx2_ASAP7_75t_L g6008 ( 
.A(n_5557),
.Y(n_6008)
);

HB1xp67_ASAP7_75t_L g6009 ( 
.A(n_5475),
.Y(n_6009)
);

INVx2_ASAP7_75t_L g6010 ( 
.A(n_5562),
.Y(n_6010)
);

INVx1_ASAP7_75t_L g6011 ( 
.A(n_5679),
.Y(n_6011)
);

NAND2xp5_ASAP7_75t_L g6012 ( 
.A(n_5645),
.B(n_5126),
.Y(n_6012)
);

INVx3_ASAP7_75t_L g6013 ( 
.A(n_5430),
.Y(n_6013)
);

INVx4_ASAP7_75t_R g6014 ( 
.A(n_5563),
.Y(n_6014)
);

INVxp67_ASAP7_75t_L g6015 ( 
.A(n_5622),
.Y(n_6015)
);

AND2x2_ASAP7_75t_L g6016 ( 
.A(n_5437),
.B(n_5074),
.Y(n_6016)
);

OR2x2_ASAP7_75t_L g6017 ( 
.A(n_5434),
.B(n_5235),
.Y(n_6017)
);

AND2x2_ASAP7_75t_L g6018 ( 
.A(n_5437),
.B(n_5080),
.Y(n_6018)
);

NAND2xp5_ASAP7_75t_L g6019 ( 
.A(n_5656),
.B(n_5127),
.Y(n_6019)
);

AND2x2_ASAP7_75t_L g6020 ( 
.A(n_5439),
.B(n_5080),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5698),
.Y(n_6021)
);

INVx2_ASAP7_75t_L g6022 ( 
.A(n_5562),
.Y(n_6022)
);

HB1xp67_ASAP7_75t_L g6023 ( 
.A(n_5478),
.Y(n_6023)
);

INVx1_ASAP7_75t_L g6024 ( 
.A(n_5699),
.Y(n_6024)
);

NAND2xp5_ASAP7_75t_L g6025 ( 
.A(n_5634),
.B(n_5127),
.Y(n_6025)
);

AND2x2_ASAP7_75t_L g6026 ( 
.A(n_5439),
.B(n_4221),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_5652),
.B(n_4221),
.Y(n_6027)
);

INVx1_ASAP7_75t_L g6028 ( 
.A(n_5694),
.Y(n_6028)
);

NAND2xp5_ASAP7_75t_L g6029 ( 
.A(n_5634),
.B(n_5467),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5478),
.Y(n_6030)
);

INVx1_ASAP7_75t_L g6031 ( 
.A(n_5480),
.Y(n_6031)
);

AND2x2_ASAP7_75t_L g6032 ( 
.A(n_5652),
.B(n_4221),
.Y(n_6032)
);

INVx2_ASAP7_75t_L g6033 ( 
.A(n_5575),
.Y(n_6033)
);

NOR2xp33_ASAP7_75t_L g6034 ( 
.A(n_5577),
.B(n_4248),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5480),
.Y(n_6035)
);

AND2x2_ASAP7_75t_L g6036 ( 
.A(n_5356),
.B(n_4301),
.Y(n_6036)
);

AND2x2_ASAP7_75t_L g6037 ( 
.A(n_5356),
.B(n_4301),
.Y(n_6037)
);

AO21x2_ASAP7_75t_L g6038 ( 
.A1(n_5519),
.A2(n_5299),
.B(n_5018),
.Y(n_6038)
);

NAND2xp5_ASAP7_75t_L g6039 ( 
.A(n_5425),
.B(n_5133),
.Y(n_6039)
);

OR2x2_ASAP7_75t_L g6040 ( 
.A(n_5359),
.B(n_4972),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5483),
.Y(n_6041)
);

INVx2_ASAP7_75t_L g6042 ( 
.A(n_5575),
.Y(n_6042)
);

INVx2_ASAP7_75t_L g6043 ( 
.A(n_5580),
.Y(n_6043)
);

OR2x2_ASAP7_75t_L g6044 ( 
.A(n_5972),
.B(n_5709),
.Y(n_6044)
);

INVxp67_ASAP7_75t_SL g6045 ( 
.A(n_5943),
.Y(n_6045)
);

INVx1_ASAP7_75t_L g6046 ( 
.A(n_5990),
.Y(n_6046)
);

NAND2xp5_ASAP7_75t_L g6047 ( 
.A(n_5701),
.B(n_5483),
.Y(n_6047)
);

INVx1_ASAP7_75t_L g6048 ( 
.A(n_5990),
.Y(n_6048)
);

NAND4xp25_ASAP7_75t_L g6049 ( 
.A(n_5904),
.B(n_5961),
.C(n_5988),
.D(n_5987),
.Y(n_6049)
);

AND2x2_ASAP7_75t_L g6050 ( 
.A(n_5717),
.B(n_5357),
.Y(n_6050)
);

NAND2xp5_ASAP7_75t_L g6051 ( 
.A(n_5701),
.B(n_5484),
.Y(n_6051)
);

INVx1_ASAP7_75t_SL g6052 ( 
.A(n_5842),
.Y(n_6052)
);

HB1xp67_ASAP7_75t_L g6053 ( 
.A(n_5794),
.Y(n_6053)
);

INVx1_ASAP7_75t_L g6054 ( 
.A(n_5995),
.Y(n_6054)
);

INVx2_ASAP7_75t_L g6055 ( 
.A(n_5858),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5995),
.Y(n_6056)
);

INVx2_ASAP7_75t_L g6057 ( 
.A(n_5858),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_5997),
.Y(n_6058)
);

NAND2xp5_ASAP7_75t_L g6059 ( 
.A(n_5802),
.B(n_5484),
.Y(n_6059)
);

OR2x6_ASAP7_75t_L g6060 ( 
.A(n_5732),
.B(n_5633),
.Y(n_6060)
);

INVx2_ASAP7_75t_L g6061 ( 
.A(n_5858),
.Y(n_6061)
);

AND2x6_ASAP7_75t_SL g6062 ( 
.A(n_5943),
.B(n_5633),
.Y(n_6062)
);

INVx1_ASAP7_75t_L g6063 ( 
.A(n_5997),
.Y(n_6063)
);

INVx2_ASAP7_75t_L g6064 ( 
.A(n_5858),
.Y(n_6064)
);

HB1xp67_ASAP7_75t_L g6065 ( 
.A(n_5795),
.Y(n_6065)
);

INVx1_ASAP7_75t_L g6066 ( 
.A(n_6009),
.Y(n_6066)
);

NAND3xp33_ASAP7_75t_L g6067 ( 
.A(n_5961),
.B(n_5476),
.C(n_5640),
.Y(n_6067)
);

OAI211xp5_ASAP7_75t_L g6068 ( 
.A1(n_5923),
.A2(n_5489),
.B(n_5357),
.C(n_5360),
.Y(n_6068)
);

INVx1_ASAP7_75t_L g6069 ( 
.A(n_6009),
.Y(n_6069)
);

INVx1_ASAP7_75t_L g6070 ( 
.A(n_6023),
.Y(n_6070)
);

A2O1A1Ixp33_ASAP7_75t_L g6071 ( 
.A1(n_5951),
.A2(n_5429),
.B(n_5640),
.C(n_5650),
.Y(n_6071)
);

NAND4xp25_ASAP7_75t_L g6072 ( 
.A(n_5904),
.B(n_5360),
.C(n_5362),
.D(n_5598),
.Y(n_6072)
);

OR2x6_ASAP7_75t_SL g6073 ( 
.A(n_5985),
.B(n_5880),
.Y(n_6073)
);

INVx1_ASAP7_75t_L g6074 ( 
.A(n_6023),
.Y(n_6074)
);

INVx2_ASAP7_75t_SL g6075 ( 
.A(n_5855),
.Y(n_6075)
);

INVx1_ASAP7_75t_L g6076 ( 
.A(n_5724),
.Y(n_6076)
);

INVx1_ASAP7_75t_L g6077 ( 
.A(n_5724),
.Y(n_6077)
);

OR2x2_ASAP7_75t_L g6078 ( 
.A(n_5940),
.B(n_5492),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5740),
.Y(n_6079)
);

INVx2_ASAP7_75t_L g6080 ( 
.A(n_5732),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_5740),
.Y(n_6081)
);

CKINVDCx20_ASAP7_75t_R g6082 ( 
.A(n_5880),
.Y(n_6082)
);

INVx2_ASAP7_75t_L g6083 ( 
.A(n_5732),
.Y(n_6083)
);

CKINVDCx20_ASAP7_75t_R g6084 ( 
.A(n_5784),
.Y(n_6084)
);

AND2x2_ASAP7_75t_L g6085 ( 
.A(n_5704),
.B(n_5705),
.Y(n_6085)
);

INVx2_ASAP7_75t_L g6086 ( 
.A(n_5732),
.Y(n_6086)
);

INVx1_ASAP7_75t_L g6087 ( 
.A(n_5777),
.Y(n_6087)
);

INVx2_ASAP7_75t_L g6088 ( 
.A(n_5762),
.Y(n_6088)
);

AND2x4_ASAP7_75t_SL g6089 ( 
.A(n_5770),
.B(n_4321),
.Y(n_6089)
);

BUFx2_ASAP7_75t_L g6090 ( 
.A(n_5757),
.Y(n_6090)
);

INVx1_ASAP7_75t_SL g6091 ( 
.A(n_5842),
.Y(n_6091)
);

OA21x2_ASAP7_75t_L g6092 ( 
.A1(n_5765),
.A2(n_5587),
.B(n_5580),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_5777),
.Y(n_6093)
);

OAI21xp33_ASAP7_75t_L g6094 ( 
.A1(n_5951),
.A2(n_5890),
.B(n_5935),
.Y(n_6094)
);

AND2x2_ASAP7_75t_L g6095 ( 
.A(n_5702),
.B(n_5381),
.Y(n_6095)
);

OR2x2_ASAP7_75t_L g6096 ( 
.A(n_5738),
.B(n_5411),
.Y(n_6096)
);

INVxp67_ASAP7_75t_L g6097 ( 
.A(n_5827),
.Y(n_6097)
);

INVx1_ASAP7_75t_L g6098 ( 
.A(n_5860),
.Y(n_6098)
);

INVx2_ASAP7_75t_L g6099 ( 
.A(n_5762),
.Y(n_6099)
);

BUFx3_ASAP7_75t_L g6100 ( 
.A(n_5784),
.Y(n_6100)
);

AO21x2_ASAP7_75t_L g6101 ( 
.A1(n_5802),
.A2(n_5420),
.B(n_5417),
.Y(n_6101)
);

INVx1_ASAP7_75t_SL g6102 ( 
.A(n_5985),
.Y(n_6102)
);

INVx4_ASAP7_75t_SL g6103 ( 
.A(n_5715),
.Y(n_6103)
);

INVx2_ASAP7_75t_L g6104 ( 
.A(n_5762),
.Y(n_6104)
);

NAND2xp5_ASAP7_75t_L g6105 ( 
.A(n_5876),
.B(n_5490),
.Y(n_6105)
);

OAI211xp5_ASAP7_75t_L g6106 ( 
.A1(n_5923),
.A2(n_5456),
.B(n_5493),
.C(n_5430),
.Y(n_6106)
);

INVx2_ASAP7_75t_SL g6107 ( 
.A(n_5855),
.Y(n_6107)
);

NOR2xp33_ASAP7_75t_L g6108 ( 
.A(n_5903),
.B(n_6001),
.Y(n_6108)
);

A2O1A1Ixp33_ASAP7_75t_L g6109 ( 
.A1(n_5765),
.A2(n_5086),
.B(n_5012),
.C(n_5490),
.Y(n_6109)
);

NOR2xp33_ASAP7_75t_L g6110 ( 
.A(n_5903),
.B(n_6001),
.Y(n_6110)
);

INVx1_ASAP7_75t_L g6111 ( 
.A(n_5860),
.Y(n_6111)
);

OR2x6_ASAP7_75t_L g6112 ( 
.A(n_5762),
.B(n_4248),
.Y(n_6112)
);

A2O1A1Ixp33_ASAP7_75t_L g6113 ( 
.A1(n_5792),
.A2(n_5086),
.B(n_5012),
.C(n_5518),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_5803),
.Y(n_6114)
);

HB1xp67_ASAP7_75t_L g6115 ( 
.A(n_5743),
.Y(n_6115)
);

AND2x2_ASAP7_75t_L g6116 ( 
.A(n_5703),
.B(n_5384),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5803),
.Y(n_6117)
);

OA21x2_ASAP7_75t_L g6118 ( 
.A1(n_5792),
.A2(n_5594),
.B(n_5587),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5817),
.Y(n_6119)
);

NOR2xp33_ASAP7_75t_L g6120 ( 
.A(n_5903),
.B(n_5384),
.Y(n_6120)
);

INVx2_ASAP7_75t_L g6121 ( 
.A(n_5834),
.Y(n_6121)
);

OA21x2_ASAP7_75t_L g6122 ( 
.A1(n_5890),
.A2(n_5599),
.B(n_5594),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_5817),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_5876),
.Y(n_6124)
);

A2O1A1Ixp33_ASAP7_75t_L g6125 ( 
.A1(n_5840),
.A2(n_5518),
.B(n_5054),
.C(n_5055),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5881),
.Y(n_6126)
);

INVxp67_ASAP7_75t_L g6127 ( 
.A(n_5976),
.Y(n_6127)
);

INVx2_ASAP7_75t_L g6128 ( 
.A(n_5834),
.Y(n_6128)
);

CKINVDCx16_ASAP7_75t_R g6129 ( 
.A(n_5715),
.Y(n_6129)
);

INVx2_ASAP7_75t_L g6130 ( 
.A(n_5834),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_5881),
.Y(n_6131)
);

AND2x4_ASAP7_75t_L g6132 ( 
.A(n_5773),
.B(n_5443),
.Y(n_6132)
);

INVx2_ASAP7_75t_SL g6133 ( 
.A(n_5855),
.Y(n_6133)
);

OAI21x1_ASAP7_75t_L g6134 ( 
.A1(n_5850),
.A2(n_5493),
.B(n_5456),
.Y(n_6134)
);

AND2x4_ASAP7_75t_L g6135 ( 
.A(n_5741),
.B(n_5443),
.Y(n_6135)
);

NAND2xp5_ASAP7_75t_SL g6136 ( 
.A(n_5772),
.B(n_5443),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_5887),
.Y(n_6137)
);

BUFx3_ASAP7_75t_L g6138 ( 
.A(n_5987),
.Y(n_6138)
);

OAI21xp5_ASAP7_75t_SL g6139 ( 
.A1(n_5935),
.A2(n_5458),
.B(n_5340),
.Y(n_6139)
);

INVx4_ASAP7_75t_SL g6140 ( 
.A(n_5757),
.Y(n_6140)
);

OAI21xp33_ASAP7_75t_L g6141 ( 
.A1(n_5992),
.A2(n_5502),
.B(n_5498),
.Y(n_6141)
);

BUFx3_ASAP7_75t_L g6142 ( 
.A(n_5988),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_5887),
.Y(n_6143)
);

A2O1A1Ixp33_ASAP7_75t_L g6144 ( 
.A1(n_5992),
.A2(n_5032),
.B(n_4962),
.C(n_4977),
.Y(n_6144)
);

OAI21xp5_ASAP7_75t_L g6145 ( 
.A1(n_6003),
.A2(n_5368),
.B(n_5665),
.Y(n_6145)
);

NAND2xp5_ASAP7_75t_SL g6146 ( 
.A(n_5772),
.B(n_5375),
.Y(n_6146)
);

AOI21xp5_ASAP7_75t_L g6147 ( 
.A1(n_6003),
.A2(n_5554),
.B(n_5550),
.Y(n_6147)
);

OA21x2_ASAP7_75t_L g6148 ( 
.A1(n_5716),
.A2(n_5608),
.B(n_5599),
.Y(n_6148)
);

HB1xp67_ASAP7_75t_L g6149 ( 
.A(n_5767),
.Y(n_6149)
);

AOI21x1_ASAP7_75t_L g6150 ( 
.A1(n_5914),
.A2(n_5389),
.B(n_5610),
.Y(n_6150)
);

INVx4_ASAP7_75t_L g6151 ( 
.A(n_5855),
.Y(n_6151)
);

INVx2_ASAP7_75t_L g6152 ( 
.A(n_5963),
.Y(n_6152)
);

O2A1O1Ixp33_ASAP7_75t_L g6153 ( 
.A1(n_5902),
.A2(n_5920),
.B(n_5969),
.C(n_6015),
.Y(n_6153)
);

AOI21x1_ASAP7_75t_L g6154 ( 
.A1(n_5917),
.A2(n_5613),
.B(n_5610),
.Y(n_6154)
);

BUFx2_ASAP7_75t_L g6155 ( 
.A(n_5757),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_5902),
.Y(n_6156)
);

AND2x2_ASAP7_75t_L g6157 ( 
.A(n_5710),
.B(n_5654),
.Y(n_6157)
);

A2O1A1Ixp33_ASAP7_75t_L g6158 ( 
.A1(n_5841),
.A2(n_4962),
.B(n_4977),
.C(n_4958),
.Y(n_6158)
);

OAI21x1_ASAP7_75t_L g6159 ( 
.A1(n_5850),
.A2(n_5891),
.B(n_5839),
.Y(n_6159)
);

NAND2xp5_ASAP7_75t_L g6160 ( 
.A(n_5920),
.B(n_5504),
.Y(n_6160)
);

INVx1_ASAP7_75t_L g6161 ( 
.A(n_5969),
.Y(n_6161)
);

INVx2_ASAP7_75t_L g6162 ( 
.A(n_5963),
.Y(n_6162)
);

AND2x2_ASAP7_75t_L g6163 ( 
.A(n_5710),
.B(n_5658),
.Y(n_6163)
);

NOR2x1_ASAP7_75t_L g6164 ( 
.A(n_6001),
.B(n_5456),
.Y(n_6164)
);

INVx3_ASAP7_75t_L g6165 ( 
.A(n_5805),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_5707),
.Y(n_6166)
);

AND2x2_ASAP7_75t_L g6167 ( 
.A(n_5713),
.B(n_5658),
.Y(n_6167)
);

OAI21x1_ASAP7_75t_L g6168 ( 
.A1(n_5850),
.A2(n_5496),
.B(n_5493),
.Y(n_6168)
);

INVx2_ASAP7_75t_L g6169 ( 
.A(n_5963),
.Y(n_6169)
);

HB1xp67_ASAP7_75t_L g6170 ( 
.A(n_5771),
.Y(n_6170)
);

INVx2_ASAP7_75t_L g6171 ( 
.A(n_6002),
.Y(n_6171)
);

INVx1_ASAP7_75t_L g6172 ( 
.A(n_5748),
.Y(n_6172)
);

AND2x4_ASAP7_75t_L g6173 ( 
.A(n_5741),
.B(n_5758),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_5748),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_5749),
.Y(n_6175)
);

INVx4_ASAP7_75t_L g6176 ( 
.A(n_5807),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_5749),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_5750),
.Y(n_6178)
);

OAI21xp5_ASAP7_75t_L g6179 ( 
.A1(n_6015),
.A2(n_5595),
.B(n_5579),
.Y(n_6179)
);

INVx1_ASAP7_75t_SL g6180 ( 
.A(n_5722),
.Y(n_6180)
);

AND2x2_ASAP7_75t_L g6181 ( 
.A(n_5713),
.B(n_5661),
.Y(n_6181)
);

INVx3_ASAP7_75t_L g6182 ( 
.A(n_5805),
.Y(n_6182)
);

OAI211xp5_ASAP7_75t_L g6183 ( 
.A1(n_5736),
.A2(n_5513),
.B(n_5603),
.C(n_5496),
.Y(n_6183)
);

INVx1_ASAP7_75t_L g6184 ( 
.A(n_5750),
.Y(n_6184)
);

AO21x2_ASAP7_75t_L g6185 ( 
.A1(n_5716),
.A2(n_5420),
.B(n_5417),
.Y(n_6185)
);

AND2x4_ASAP7_75t_L g6186 ( 
.A(n_5758),
.B(n_5661),
.Y(n_6186)
);

NAND2xp5_ASAP7_75t_L g6187 ( 
.A(n_5711),
.B(n_5505),
.Y(n_6187)
);

INVx1_ASAP7_75t_L g6188 ( 
.A(n_5753),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_5753),
.Y(n_6189)
);

INVx2_ASAP7_75t_L g6190 ( 
.A(n_6002),
.Y(n_6190)
);

CKINVDCx20_ASAP7_75t_R g6191 ( 
.A(n_6006),
.Y(n_6191)
);

AND2x4_ASAP7_75t_L g6192 ( 
.A(n_5805),
.B(n_5809),
.Y(n_6192)
);

INVx1_ASAP7_75t_L g6193 ( 
.A(n_5779),
.Y(n_6193)
);

NAND2xp5_ASAP7_75t_L g6194 ( 
.A(n_5712),
.B(n_5514),
.Y(n_6194)
);

INVx1_ASAP7_75t_L g6195 ( 
.A(n_5779),
.Y(n_6195)
);

NAND2xp5_ASAP7_75t_L g6196 ( 
.A(n_6030),
.B(n_5523),
.Y(n_6196)
);

HB1xp67_ASAP7_75t_L g6197 ( 
.A(n_5938),
.Y(n_6197)
);

INVx2_ASAP7_75t_L g6198 ( 
.A(n_6002),
.Y(n_6198)
);

AOI21xp5_ASAP7_75t_L g6199 ( 
.A1(n_6038),
.A2(n_5554),
.B(n_5606),
.Y(n_6199)
);

NAND2xp5_ASAP7_75t_L g6200 ( 
.A(n_6031),
.B(n_5583),
.Y(n_6200)
);

OR2x2_ASAP7_75t_SL g6201 ( 
.A(n_5725),
.B(n_5418),
.Y(n_6201)
);

NAND2xp5_ASAP7_75t_L g6202 ( 
.A(n_6035),
.B(n_6041),
.Y(n_6202)
);

OA21x2_ASAP7_75t_L g6203 ( 
.A1(n_5719),
.A2(n_5608),
.B(n_5423),
.Y(n_6203)
);

NAND2xp5_ASAP7_75t_L g6204 ( 
.A(n_6028),
.B(n_5589),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_5781),
.Y(n_6205)
);

INVx2_ASAP7_75t_L g6206 ( 
.A(n_5733),
.Y(n_6206)
);

INVxp67_ASAP7_75t_SL g6207 ( 
.A(n_5976),
.Y(n_6207)
);

AND2x4_ASAP7_75t_L g6208 ( 
.A(n_5809),
.B(n_5664),
.Y(n_6208)
);

INVx2_ASAP7_75t_SL g6209 ( 
.A(n_5809),
.Y(n_6209)
);

INVx2_ASAP7_75t_L g6210 ( 
.A(n_5733),
.Y(n_6210)
);

OA21x2_ASAP7_75t_L g6211 ( 
.A1(n_5719),
.A2(n_5423),
.B(n_5422),
.Y(n_6211)
);

NAND2xp5_ASAP7_75t_L g6212 ( 
.A(n_5774),
.B(n_5596),
.Y(n_6212)
);

INVx2_ASAP7_75t_L g6213 ( 
.A(n_5733),
.Y(n_6213)
);

OAI21x1_ASAP7_75t_L g6214 ( 
.A1(n_5891),
.A2(n_5513),
.B(n_5496),
.Y(n_6214)
);

INVx4_ASAP7_75t_SL g6215 ( 
.A(n_5965),
.Y(n_6215)
);

INVxp67_ASAP7_75t_SL g6216 ( 
.A(n_6006),
.Y(n_6216)
);

NAND2xp5_ASAP7_75t_L g6217 ( 
.A(n_5714),
.B(n_5621),
.Y(n_6217)
);

INVx1_ASAP7_75t_L g6218 ( 
.A(n_5781),
.Y(n_6218)
);

INVx4_ASAP7_75t_L g6219 ( 
.A(n_5807),
.Y(n_6219)
);

AND2x2_ASAP7_75t_L g6220 ( 
.A(n_5847),
.B(n_5664),
.Y(n_6220)
);

NAND2xp5_ASAP7_75t_L g6221 ( 
.A(n_5718),
.B(n_5653),
.Y(n_6221)
);

AOI21xp5_ASAP7_75t_L g6222 ( 
.A1(n_6038),
.A2(n_5768),
.B(n_5864),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_5796),
.Y(n_6223)
);

A2O1A1Ixp33_ASAP7_75t_L g6224 ( 
.A1(n_6034),
.A2(n_4992),
.B(n_5001),
.C(n_4958),
.Y(n_6224)
);

INVx1_ASAP7_75t_L g6225 ( 
.A(n_5796),
.Y(n_6225)
);

NAND2xp5_ASAP7_75t_L g6226 ( 
.A(n_5721),
.B(n_5693),
.Y(n_6226)
);

BUFx2_ASAP7_75t_L g6227 ( 
.A(n_5847),
.Y(n_6227)
);

BUFx3_ASAP7_75t_L g6228 ( 
.A(n_5965),
.Y(n_6228)
);

BUFx2_ASAP7_75t_L g6229 ( 
.A(n_5847),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_5800),
.Y(n_6230)
);

AND2x4_ASAP7_75t_L g6231 ( 
.A(n_5868),
.B(n_5677),
.Y(n_6231)
);

AOI21xp5_ASAP7_75t_L g6232 ( 
.A1(n_5864),
.A2(n_5531),
.B(n_5677),
.Y(n_6232)
);

INVx2_ASAP7_75t_L g6233 ( 
.A(n_5807),
.Y(n_6233)
);

OAI211xp5_ASAP7_75t_L g6234 ( 
.A1(n_6034),
.A2(n_5825),
.B(n_5839),
.C(n_5946),
.Y(n_6234)
);

INVx1_ASAP7_75t_L g6235 ( 
.A(n_5836),
.Y(n_6235)
);

NAND2xp33_ASAP7_75t_SL g6236 ( 
.A(n_5720),
.B(n_5731),
.Y(n_6236)
);

BUFx2_ASAP7_75t_L g6237 ( 
.A(n_5868),
.Y(n_6237)
);

INVx1_ASAP7_75t_L g6238 ( 
.A(n_5836),
.Y(n_6238)
);

AOI21xp33_ASAP7_75t_SL g6239 ( 
.A1(n_5706),
.A2(n_4698),
.B(n_4683),
.Y(n_6239)
);

INVx1_ASAP7_75t_SL g6240 ( 
.A(n_5984),
.Y(n_6240)
);

HB1xp67_ASAP7_75t_L g6241 ( 
.A(n_5955),
.Y(n_6241)
);

INVx2_ASAP7_75t_L g6242 ( 
.A(n_5808),
.Y(n_6242)
);

BUFx6f_ASAP7_75t_L g6243 ( 
.A(n_5808),
.Y(n_6243)
);

AOI21xp5_ASAP7_75t_L g6244 ( 
.A1(n_5839),
.A2(n_5375),
.B(n_5089),
.Y(n_6244)
);

INVx2_ASAP7_75t_L g6245 ( 
.A(n_5808),
.Y(n_6245)
);

INVx1_ASAP7_75t_L g6246 ( 
.A(n_5852),
.Y(n_6246)
);

INVx2_ASAP7_75t_L g6247 ( 
.A(n_5896),
.Y(n_6247)
);

INVx3_ASAP7_75t_L g6248 ( 
.A(n_5868),
.Y(n_6248)
);

OA21x2_ASAP7_75t_L g6249 ( 
.A1(n_5730),
.A2(n_5431),
.B(n_5422),
.Y(n_6249)
);

INVx1_ASAP7_75t_L g6250 ( 
.A(n_5852),
.Y(n_6250)
);

INVx2_ASAP7_75t_SL g6251 ( 
.A(n_5875),
.Y(n_6251)
);

NAND4xp25_ASAP7_75t_L g6252 ( 
.A(n_5825),
.B(n_5513),
.C(n_5603),
.D(n_5375),
.Y(n_6252)
);

NAND4xp25_ASAP7_75t_L g6253 ( 
.A(n_5825),
.B(n_5603),
.C(n_4998),
.D(n_5048),
.Y(n_6253)
);

AND2x2_ASAP7_75t_L g6254 ( 
.A(n_5734),
.B(n_5581),
.Y(n_6254)
);

NOR2xp33_ASAP7_75t_R g6255 ( 
.A(n_5984),
.B(n_4342),
.Y(n_6255)
);

AOI21xp5_ASAP7_75t_L g6256 ( 
.A1(n_5772),
.A2(n_5089),
.B(n_5001),
.Y(n_6256)
);

INVx1_ASAP7_75t_L g6257 ( 
.A(n_5857),
.Y(n_6257)
);

HB1xp67_ASAP7_75t_L g6258 ( 
.A(n_6004),
.Y(n_6258)
);

HB1xp67_ASAP7_75t_L g6259 ( 
.A(n_5742),
.Y(n_6259)
);

INVx2_ASAP7_75t_L g6260 ( 
.A(n_5896),
.Y(n_6260)
);

NAND3xp33_ASAP7_75t_L g6261 ( 
.A(n_5730),
.B(n_5351),
.C(n_5349),
.Y(n_6261)
);

INVxp67_ASAP7_75t_SL g6262 ( 
.A(n_5776),
.Y(n_6262)
);

INVx2_ASAP7_75t_L g6263 ( 
.A(n_5896),
.Y(n_6263)
);

AO21x2_ASAP7_75t_L g6264 ( 
.A1(n_5857),
.A2(n_5432),
.B(n_5431),
.Y(n_6264)
);

A2O1A1Ixp33_ASAP7_75t_L g6265 ( 
.A1(n_5891),
.A2(n_5010),
.B(n_5013),
.C(n_4992),
.Y(n_6265)
);

NAND2xp33_ASAP7_75t_SL g6266 ( 
.A(n_5934),
.B(n_5485),
.Y(n_6266)
);

INVx2_ASAP7_75t_L g6267 ( 
.A(n_5875),
.Y(n_6267)
);

INVx2_ASAP7_75t_L g6268 ( 
.A(n_5875),
.Y(n_6268)
);

AOI21xp5_ASAP7_75t_L g6269 ( 
.A1(n_5974),
.A2(n_5013),
.B(n_5010),
.Y(n_6269)
);

NAND2xp5_ASAP7_75t_L g6270 ( 
.A(n_5728),
.B(n_5133),
.Y(n_6270)
);

INVx2_ASAP7_75t_L g6271 ( 
.A(n_5928),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_5865),
.Y(n_6272)
);

AND2x2_ASAP7_75t_L g6273 ( 
.A(n_5948),
.B(n_5581),
.Y(n_6273)
);

AND2x4_ASAP7_75t_L g6274 ( 
.A(n_5756),
.B(n_5629),
.Y(n_6274)
);

INVx4_ASAP7_75t_L g6275 ( 
.A(n_5726),
.Y(n_6275)
);

NAND2xp5_ASAP7_75t_L g6276 ( 
.A(n_5729),
.B(n_5135),
.Y(n_6276)
);

AO21x2_ASAP7_75t_L g6277 ( 
.A1(n_5865),
.A2(n_5432),
.B(n_5351),
.Y(n_6277)
);

OR2x2_ASAP7_75t_L g6278 ( 
.A(n_5723),
.B(n_5600),
.Y(n_6278)
);

INVx1_ASAP7_75t_L g6279 ( 
.A(n_5866),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_5866),
.Y(n_6280)
);

A2O1A1Ixp33_ASAP7_75t_L g6281 ( 
.A1(n_5766),
.A2(n_5025),
.B(n_5028),
.C(n_5022),
.Y(n_6281)
);

INVx2_ASAP7_75t_L g6282 ( 
.A(n_5928),
.Y(n_6282)
);

AND2x2_ASAP7_75t_L g6283 ( 
.A(n_5924),
.B(n_5629),
.Y(n_6283)
);

INVx1_ASAP7_75t_SL g6284 ( 
.A(n_5726),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_5869),
.Y(n_6285)
);

BUFx2_ASAP7_75t_L g6286 ( 
.A(n_5928),
.Y(n_6286)
);

INVx2_ASAP7_75t_L g6287 ( 
.A(n_5968),
.Y(n_6287)
);

INVx2_ASAP7_75t_L g6288 ( 
.A(n_5968),
.Y(n_6288)
);

AOI21xp5_ASAP7_75t_L g6289 ( 
.A1(n_5856),
.A2(n_5025),
.B(n_5022),
.Y(n_6289)
);

AOI22xp5_ASAP7_75t_L g6290 ( 
.A1(n_5766),
.A2(n_5568),
.B1(n_5571),
.B2(n_5566),
.Y(n_6290)
);

INVx4_ASAP7_75t_SL g6291 ( 
.A(n_5726),
.Y(n_6291)
);

INVx4_ASAP7_75t_L g6292 ( 
.A(n_5744),
.Y(n_6292)
);

OAI21xp33_ASAP7_75t_L g6293 ( 
.A1(n_5838),
.A2(n_4986),
.B(n_4970),
.Y(n_6293)
);

A2O1A1Ixp33_ASAP7_75t_L g6294 ( 
.A1(n_5766),
.A2(n_5029),
.B(n_5031),
.C(n_5028),
.Y(n_6294)
);

INVx2_ASAP7_75t_L g6295 ( 
.A(n_5968),
.Y(n_6295)
);

INVx2_ASAP7_75t_L g6296 ( 
.A(n_6013),
.Y(n_6296)
);

INVxp67_ASAP7_75t_SL g6297 ( 
.A(n_5925),
.Y(n_6297)
);

NAND2xp5_ASAP7_75t_L g6298 ( 
.A(n_5735),
.B(n_5135),
.Y(n_6298)
);

AND2x2_ASAP7_75t_L g6299 ( 
.A(n_5892),
.B(n_5631),
.Y(n_6299)
);

AND2x2_ASAP7_75t_L g6300 ( 
.A(n_5897),
.B(n_5631),
.Y(n_6300)
);

A2O1A1Ixp33_ASAP7_75t_L g6301 ( 
.A1(n_5791),
.A2(n_5031),
.B(n_5029),
.C(n_4799),
.Y(n_6301)
);

INVx3_ASAP7_75t_L g6302 ( 
.A(n_5744),
.Y(n_6302)
);

INVxp67_ASAP7_75t_L g6303 ( 
.A(n_5769),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_5869),
.Y(n_6304)
);

NAND2xp5_ASAP7_75t_L g6305 ( 
.A(n_5737),
.B(n_5139),
.Y(n_6305)
);

INVx2_ASAP7_75t_L g6306 ( 
.A(n_6013),
.Y(n_6306)
);

INVx2_ASAP7_75t_L g6307 ( 
.A(n_6013),
.Y(n_6307)
);

AND2x2_ASAP7_75t_L g6308 ( 
.A(n_5820),
.B(n_5642),
.Y(n_6308)
);

OR2x6_ASAP7_75t_L g6309 ( 
.A(n_5996),
.B(n_5335),
.Y(n_6309)
);

AND2x2_ASAP7_75t_L g6310 ( 
.A(n_5820),
.B(n_5642),
.Y(n_6310)
);

AOI21xp5_ASAP7_75t_L g6311 ( 
.A1(n_5859),
.A2(n_5015),
.B(n_4995),
.Y(n_6311)
);

NOR2xp33_ASAP7_75t_L g6312 ( 
.A(n_5708),
.B(n_4194),
.Y(n_6312)
);

INVx4_ASAP7_75t_L g6313 ( 
.A(n_5744),
.Y(n_6313)
);

BUFx2_ASAP7_75t_L g6314 ( 
.A(n_5708),
.Y(n_6314)
);

AND2x4_ASAP7_75t_L g6315 ( 
.A(n_5708),
.B(n_5651),
.Y(n_6315)
);

AOI21xp5_ASAP7_75t_L g6316 ( 
.A1(n_6012),
.A2(n_5015),
.B(n_5566),
.Y(n_6316)
);

INVx2_ASAP7_75t_L g6317 ( 
.A(n_5763),
.Y(n_6317)
);

INVx2_ASAP7_75t_L g6318 ( 
.A(n_5763),
.Y(n_6318)
);

INVx3_ASAP7_75t_L g6319 ( 
.A(n_6007),
.Y(n_6319)
);

AND2x2_ASAP7_75t_L g6320 ( 
.A(n_5829),
.B(n_5651),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_5871),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_5871),
.Y(n_6322)
);

AND2x2_ASAP7_75t_L g6323 ( 
.A(n_5829),
.B(n_5485),
.Y(n_6323)
);

INVx2_ASAP7_75t_SL g6324 ( 
.A(n_6014),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_5879),
.Y(n_6325)
);

NAND2xp5_ASAP7_75t_L g6326 ( 
.A(n_5746),
.B(n_5139),
.Y(n_6326)
);

OAI21x1_ASAP7_75t_L g6327 ( 
.A1(n_5791),
.A2(n_5683),
.B(n_5681),
.Y(n_6327)
);

AND2x4_ASAP7_75t_L g6328 ( 
.A(n_5883),
.B(n_5495),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_5879),
.Y(n_6329)
);

O2A1O1Ixp33_ASAP7_75t_L g6330 ( 
.A1(n_5764),
.A2(n_4986),
.B(n_4998),
.C(n_4970),
.Y(n_6330)
);

INVx2_ASAP7_75t_L g6331 ( 
.A(n_5837),
.Y(n_6331)
);

INVx1_ASAP7_75t_L g6332 ( 
.A(n_5882),
.Y(n_6332)
);

INVx5_ASAP7_75t_L g6333 ( 
.A(n_5793),
.Y(n_6333)
);

INVx3_ASAP7_75t_L g6334 ( 
.A(n_6007),
.Y(n_6334)
);

BUFx3_ASAP7_75t_L g6335 ( 
.A(n_5739),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_5882),
.Y(n_6336)
);

AND2x2_ASAP7_75t_L g6337 ( 
.A(n_5837),
.B(n_5843),
.Y(n_6337)
);

INVx2_ASAP7_75t_L g6338 ( 
.A(n_5843),
.Y(n_6338)
);

AND2x2_ASAP7_75t_L g6339 ( 
.A(n_5884),
.B(n_5495),
.Y(n_6339)
);

INVx2_ASAP7_75t_L g6340 ( 
.A(n_5791),
.Y(n_6340)
);

AND2x2_ASAP7_75t_L g6341 ( 
.A(n_5885),
.B(n_5510),
.Y(n_6341)
);

INVx1_ASAP7_75t_L g6342 ( 
.A(n_6053),
.Y(n_6342)
);

NOR2x1_ASAP7_75t_L g6343 ( 
.A(n_6191),
.B(n_5747),
.Y(n_6343)
);

NAND2xp5_ASAP7_75t_SL g6344 ( 
.A(n_6255),
.B(n_6007),
.Y(n_6344)
);

AND2x2_ASAP7_75t_L g6345 ( 
.A(n_6089),
.B(n_5745),
.Y(n_6345)
);

NAND2xp5_ASAP7_75t_L g6346 ( 
.A(n_6207),
.B(n_5905),
.Y(n_6346)
);

INVx2_ASAP7_75t_L g6347 ( 
.A(n_6215),
.Y(n_6347)
);

NAND2xp5_ASAP7_75t_L g6348 ( 
.A(n_6240),
.B(n_5905),
.Y(n_6348)
);

AO21x2_ASAP7_75t_L g6349 ( 
.A1(n_6094),
.A2(n_5913),
.B(n_5888),
.Y(n_6349)
);

NAND2xp5_ASAP7_75t_L g6350 ( 
.A(n_6240),
.B(n_5889),
.Y(n_6350)
);

NAND2xp5_ASAP7_75t_L g6351 ( 
.A(n_6216),
.B(n_5727),
.Y(n_6351)
);

AOI22xp33_ASAP7_75t_L g6352 ( 
.A1(n_6094),
.A2(n_6047),
.B1(n_6059),
.B2(n_6051),
.Y(n_6352)
);

INVx3_ASAP7_75t_L g6353 ( 
.A(n_6192),
.Y(n_6353)
);

AND2x2_ASAP7_75t_L g6354 ( 
.A(n_6337),
.B(n_5751),
.Y(n_6354)
);

AO21x2_ASAP7_75t_L g6355 ( 
.A1(n_6067),
.A2(n_5913),
.B(n_5888),
.Y(n_6355)
);

INVx1_ASAP7_75t_L g6356 ( 
.A(n_6065),
.Y(n_6356)
);

OR2x2_ASAP7_75t_L g6357 ( 
.A(n_6044),
.B(n_5831),
.Y(n_6357)
);

NAND3xp33_ASAP7_75t_L g6358 ( 
.A(n_6139),
.B(n_5861),
.C(n_5793),
.Y(n_6358)
);

OAI21xp5_ASAP7_75t_L g6359 ( 
.A1(n_6139),
.A2(n_5835),
.B(n_5786),
.Y(n_6359)
);

INVx1_ASAP7_75t_L g6360 ( 
.A(n_6258),
.Y(n_6360)
);

NOR3xp33_ASAP7_75t_L g6361 ( 
.A(n_6129),
.B(n_5861),
.C(n_6029),
.Y(n_6361)
);

INVx2_ASAP7_75t_L g6362 ( 
.A(n_6215),
.Y(n_6362)
);

INVx1_ASAP7_75t_L g6363 ( 
.A(n_6115),
.Y(n_6363)
);

AND2x2_ASAP7_75t_L g6364 ( 
.A(n_6050),
.B(n_5906),
.Y(n_6364)
);

AOI22xp33_ASAP7_75t_L g6365 ( 
.A1(n_6047),
.A2(n_5091),
.B1(n_5926),
.B2(n_5929),
.Y(n_6365)
);

OR2x2_ASAP7_75t_L g6366 ( 
.A(n_6180),
.B(n_5761),
.Y(n_6366)
);

AOI22xp33_ASAP7_75t_L g6367 ( 
.A1(n_6051),
.A2(n_5091),
.B1(n_5926),
.B2(n_5929),
.Y(n_6367)
);

INVx1_ASAP7_75t_L g6368 ( 
.A(n_6149),
.Y(n_6368)
);

AO21x2_ASAP7_75t_L g6369 ( 
.A1(n_6067),
.A2(n_5941),
.B(n_5939),
.Y(n_6369)
);

NOR3xp33_ASAP7_75t_L g6370 ( 
.A(n_6102),
.B(n_5977),
.C(n_5754),
.Y(n_6370)
);

NAND3xp33_ASAP7_75t_L g6371 ( 
.A(n_6071),
.B(n_5977),
.C(n_5953),
.Y(n_6371)
);

AOI221xp5_ASAP7_75t_L g6372 ( 
.A1(n_6222),
.A2(n_6039),
.B1(n_6019),
.B2(n_5867),
.C(n_5863),
.Y(n_6372)
);

NAND3xp33_ASAP7_75t_L g6373 ( 
.A(n_6199),
.B(n_5755),
.C(n_5975),
.Y(n_6373)
);

NAND4xp75_ASAP7_75t_L g6374 ( 
.A(n_6147),
.B(n_5978),
.C(n_5918),
.D(n_5921),
.Y(n_6374)
);

OR2x2_ASAP7_75t_L g6375 ( 
.A(n_6180),
.B(n_5759),
.Y(n_6375)
);

AND2x4_ASAP7_75t_L g6376 ( 
.A(n_6291),
.B(n_5907),
.Y(n_6376)
);

INVx2_ASAP7_75t_L g6377 ( 
.A(n_6319),
.Y(n_6377)
);

AOI221xp5_ASAP7_75t_L g6378 ( 
.A1(n_6125),
.A2(n_5775),
.B1(n_5787),
.B2(n_5780),
.C(n_5752),
.Y(n_6378)
);

INVx1_ASAP7_75t_L g6379 ( 
.A(n_6170),
.Y(n_6379)
);

AOI22xp5_ASAP7_75t_L g6380 ( 
.A1(n_6059),
.A2(n_5789),
.B1(n_5797),
.B2(n_5788),
.Y(n_6380)
);

AND2x2_ASAP7_75t_L g6381 ( 
.A(n_6308),
.B(n_6036),
.Y(n_6381)
);

NOR2xp33_ASAP7_75t_L g6382 ( 
.A(n_6082),
.B(n_5760),
.Y(n_6382)
);

AOI221xp5_ASAP7_75t_L g6383 ( 
.A1(n_6109),
.A2(n_6024),
.B1(n_6021),
.B2(n_5814),
.C(n_5816),
.Y(n_6383)
);

NAND2xp5_ASAP7_75t_L g6384 ( 
.A(n_6045),
.B(n_6310),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_6076),
.Y(n_6385)
);

AND2x2_ASAP7_75t_L g6386 ( 
.A(n_6320),
.B(n_6037),
.Y(n_6386)
);

BUFx3_ASAP7_75t_L g6387 ( 
.A(n_6084),
.Y(n_6387)
);

AND2x2_ASAP7_75t_L g6388 ( 
.A(n_6273),
.B(n_6254),
.Y(n_6388)
);

NOR3xp33_ASAP7_75t_L g6389 ( 
.A(n_6102),
.B(n_5873),
.C(n_5939),
.Y(n_6389)
);

AND2x2_ASAP7_75t_L g6390 ( 
.A(n_6085),
.B(n_6027),
.Y(n_6390)
);

OAI211xp5_ASAP7_75t_SL g6391 ( 
.A1(n_6068),
.A2(n_5900),
.B(n_6017),
.C(n_5973),
.Y(n_6391)
);

NAND3xp33_ASAP7_75t_L g6392 ( 
.A(n_6097),
.B(n_5755),
.C(n_6025),
.Y(n_6392)
);

AOI22xp33_ASAP7_75t_L g6393 ( 
.A1(n_6118),
.A2(n_5942),
.B1(n_5944),
.B2(n_5941),
.Y(n_6393)
);

OR2x2_ASAP7_75t_L g6394 ( 
.A(n_6278),
.B(n_5927),
.Y(n_6394)
);

OAI21xp5_ASAP7_75t_L g6395 ( 
.A1(n_6113),
.A2(n_5921),
.B(n_5918),
.Y(n_6395)
);

INVx1_ASAP7_75t_L g6396 ( 
.A(n_6077),
.Y(n_6396)
);

OAI31xp33_ASAP7_75t_L g6397 ( 
.A1(n_6301),
.A2(n_5571),
.A3(n_5568),
.B(n_5930),
.Y(n_6397)
);

NOR2xp33_ASAP7_75t_L g6398 ( 
.A(n_6127),
.B(n_6032),
.Y(n_6398)
);

AND2x2_ASAP7_75t_L g6399 ( 
.A(n_6299),
.B(n_6300),
.Y(n_6399)
);

NAND3xp33_ASAP7_75t_L g6400 ( 
.A(n_6153),
.B(n_5755),
.C(n_6011),
.Y(n_6400)
);

INVxp67_ASAP7_75t_L g6401 ( 
.A(n_6073),
.Y(n_6401)
);

OR2x2_ASAP7_75t_L g6402 ( 
.A(n_6078),
.B(n_5886),
.Y(n_6402)
);

AND2x2_ASAP7_75t_L g6403 ( 
.A(n_6157),
.B(n_6163),
.Y(n_6403)
);

AND2x4_ASAP7_75t_L g6404 ( 
.A(n_6291),
.B(n_5908),
.Y(n_6404)
);

AND2x2_ASAP7_75t_L g6405 ( 
.A(n_6167),
.B(n_5911),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_6079),
.Y(n_6406)
);

NOR3xp33_ASAP7_75t_L g6407 ( 
.A(n_6049),
.B(n_5944),
.C(n_5942),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_6081),
.Y(n_6408)
);

NAND3xp33_ASAP7_75t_L g6409 ( 
.A(n_6049),
.B(n_6145),
.C(n_6197),
.Y(n_6409)
);

AND2x4_ASAP7_75t_SL g6410 ( 
.A(n_6112),
.B(n_4784),
.Y(n_6410)
);

NOR2xp33_ASAP7_75t_L g6411 ( 
.A(n_6275),
.B(n_5851),
.Y(n_6411)
);

INVx1_ASAP7_75t_L g6412 ( 
.A(n_6087),
.Y(n_6412)
);

AOI22xp33_ASAP7_75t_L g6413 ( 
.A1(n_6118),
.A2(n_5956),
.B1(n_5970),
.B2(n_5950),
.Y(n_6413)
);

NAND3xp33_ASAP7_75t_L g6414 ( 
.A(n_6145),
.B(n_5799),
.C(n_5798),
.Y(n_6414)
);

AOI221xp5_ASAP7_75t_L g6415 ( 
.A1(n_6232),
.A2(n_5823),
.B1(n_5826),
.B2(n_5822),
.C(n_5821),
.Y(n_6415)
);

NAND3xp33_ASAP7_75t_L g6416 ( 
.A(n_6241),
.B(n_6005),
.C(n_5848),
.Y(n_6416)
);

NOR3xp33_ASAP7_75t_L g6417 ( 
.A(n_6052),
.B(n_6091),
.C(n_6234),
.Y(n_6417)
);

AND2x2_ASAP7_75t_L g6418 ( 
.A(n_6181),
.B(n_6026),
.Y(n_6418)
);

AND2x2_ASAP7_75t_L g6419 ( 
.A(n_6283),
.B(n_5978),
.Y(n_6419)
);

OAI22xp33_ASAP7_75t_L g6420 ( 
.A1(n_6105),
.A2(n_5996),
.B1(n_5252),
.B2(n_5249),
.Y(n_6420)
);

NAND2xp5_ASAP7_75t_L g6421 ( 
.A(n_6259),
.B(n_5964),
.Y(n_6421)
);

AND2x2_ASAP7_75t_L g6422 ( 
.A(n_6339),
.B(n_5778),
.Y(n_6422)
);

INVx2_ASAP7_75t_L g6423 ( 
.A(n_6319),
.Y(n_6423)
);

AND2x2_ASAP7_75t_L g6424 ( 
.A(n_6341),
.B(n_5782),
.Y(n_6424)
);

AO21x2_ASAP7_75t_L g6425 ( 
.A1(n_6154),
.A2(n_5956),
.B(n_5950),
.Y(n_6425)
);

NAND4xp75_ASAP7_75t_L g6426 ( 
.A(n_6092),
.B(n_5806),
.C(n_5810),
.D(n_5801),
.Y(n_6426)
);

AND2x2_ASAP7_75t_L g6427 ( 
.A(n_6323),
.B(n_5845),
.Y(n_6427)
);

AOI22xp5_ASAP7_75t_L g6428 ( 
.A1(n_6122),
.A2(n_5849),
.B1(n_5853),
.B2(n_5844),
.Y(n_6428)
);

OR2x2_ASAP7_75t_L g6429 ( 
.A(n_6331),
.B(n_5933),
.Y(n_6429)
);

NAND3xp33_ASAP7_75t_L g6430 ( 
.A(n_6098),
.B(n_5999),
.C(n_5998),
.Y(n_6430)
);

NAND3xp33_ASAP7_75t_L g6431 ( 
.A(n_6111),
.B(n_5862),
.C(n_5854),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_6093),
.Y(n_6432)
);

AOI22xp33_ASAP7_75t_L g6433 ( 
.A1(n_6092),
.A2(n_5971),
.B1(n_5979),
.B2(n_5970),
.Y(n_6433)
);

NAND2xp5_ASAP7_75t_L g6434 ( 
.A(n_6228),
.B(n_5986),
.Y(n_6434)
);

NAND2xp5_ASAP7_75t_SL g6435 ( 
.A(n_6173),
.B(n_5949),
.Y(n_6435)
);

NOR3xp33_ASAP7_75t_L g6436 ( 
.A(n_6052),
.B(n_5979),
.C(n_5971),
.Y(n_6436)
);

OR2x2_ASAP7_75t_L g6437 ( 
.A(n_6338),
.B(n_6040),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_6114),
.Y(n_6438)
);

INVx2_ASAP7_75t_L g6439 ( 
.A(n_6334),
.Y(n_6439)
);

AOI22xp33_ASAP7_75t_L g6440 ( 
.A1(n_6101),
.A2(n_5983),
.B1(n_5989),
.B2(n_5980),
.Y(n_6440)
);

NAND2xp5_ASAP7_75t_L g6441 ( 
.A(n_6138),
.B(n_5870),
.Y(n_6441)
);

AND2x2_ASAP7_75t_L g6442 ( 
.A(n_6274),
.B(n_6315),
.Y(n_6442)
);

OR2x2_ASAP7_75t_L g6443 ( 
.A(n_6212),
.B(n_5910),
.Y(n_6443)
);

NOR2xp33_ASAP7_75t_L g6444 ( 
.A(n_6275),
.B(n_5925),
.Y(n_6444)
);

OR2x2_ASAP7_75t_L g6445 ( 
.A(n_6212),
.B(n_5936),
.Y(n_6445)
);

AOI22xp33_ASAP7_75t_SL g6446 ( 
.A1(n_6122),
.A2(n_5996),
.B1(n_5208),
.B2(n_5170),
.Y(n_6446)
);

AND2x2_ASAP7_75t_L g6447 ( 
.A(n_6274),
.B(n_5846),
.Y(n_6447)
);

NOR2xp33_ASAP7_75t_L g6448 ( 
.A(n_6292),
.B(n_6016),
.Y(n_6448)
);

OR2x2_ASAP7_75t_L g6449 ( 
.A(n_6096),
.B(n_5874),
.Y(n_6449)
);

AOI22xp33_ASAP7_75t_SL g6450 ( 
.A1(n_6334),
.A2(n_6105),
.B1(n_6048),
.B2(n_6054),
.Y(n_6450)
);

INVxp67_ASAP7_75t_L g6451 ( 
.A(n_6286),
.Y(n_6451)
);

OAI22xp5_ASAP7_75t_L g6452 ( 
.A1(n_6201),
.A2(n_5878),
.B1(n_5872),
.B2(n_5937),
.Y(n_6452)
);

OR2x2_ASAP7_75t_L g6453 ( 
.A(n_6230),
.B(n_5877),
.Y(n_6453)
);

NOR3xp33_ASAP7_75t_L g6454 ( 
.A(n_6091),
.B(n_5983),
.C(n_5980),
.Y(n_6454)
);

NOR3xp33_ASAP7_75t_L g6455 ( 
.A(n_6090),
.B(n_5994),
.C(n_5989),
.Y(n_6455)
);

AND2x4_ASAP7_75t_L g6456 ( 
.A(n_6140),
.B(n_5954),
.Y(n_6456)
);

OR2x2_ASAP7_75t_L g6457 ( 
.A(n_6194),
.B(n_5893),
.Y(n_6457)
);

NAND3xp33_ASAP7_75t_L g6458 ( 
.A(n_6117),
.B(n_5895),
.C(n_5894),
.Y(n_6458)
);

AOI22xp5_ASAP7_75t_L g6459 ( 
.A1(n_6141),
.A2(n_5899),
.B1(n_5901),
.B2(n_5898),
.Y(n_6459)
);

AOI211xp5_ASAP7_75t_L g6460 ( 
.A1(n_6141),
.A2(n_5912),
.B(n_5915),
.C(n_5909),
.Y(n_6460)
);

NAND4xp75_ASAP7_75t_L g6461 ( 
.A(n_6324),
.B(n_5806),
.C(n_5810),
.D(n_5801),
.Y(n_6461)
);

AOI22xp33_ASAP7_75t_L g6462 ( 
.A1(n_6101),
.A2(n_6000),
.B1(n_6008),
.B2(n_5994),
.Y(n_6462)
);

OA211x2_ASAP7_75t_L g6463 ( 
.A1(n_6146),
.A2(n_4370),
.B(n_3674),
.C(n_5015),
.Y(n_6463)
);

BUFx2_ASAP7_75t_SL g6464 ( 
.A(n_6142),
.Y(n_6464)
);

AND2x2_ASAP7_75t_L g6465 ( 
.A(n_6315),
.B(n_5957),
.Y(n_6465)
);

NOR3xp33_ASAP7_75t_L g6466 ( 
.A(n_6155),
.B(n_6083),
.C(n_6080),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_6119),
.Y(n_6467)
);

OR2x2_ASAP7_75t_L g6468 ( 
.A(n_6194),
.B(n_5916),
.Y(n_6468)
);

NOR3xp33_ASAP7_75t_L g6469 ( 
.A(n_6086),
.B(n_6008),
.C(n_6000),
.Y(n_6469)
);

AND2x2_ASAP7_75t_SL g6470 ( 
.A(n_6173),
.B(n_4301),
.Y(n_6470)
);

OR2x2_ASAP7_75t_L g6471 ( 
.A(n_6187),
.B(n_5919),
.Y(n_6471)
);

NAND4xp75_ASAP7_75t_L g6472 ( 
.A(n_6164),
.B(n_5812),
.C(n_5818),
.D(n_5811),
.Y(n_6472)
);

OAI211xp5_ASAP7_75t_SL g6473 ( 
.A1(n_6179),
.A2(n_5931),
.B(n_5932),
.C(n_5922),
.Y(n_6473)
);

INVx2_ASAP7_75t_SL g6474 ( 
.A(n_6192),
.Y(n_6474)
);

AO21x2_ASAP7_75t_L g6475 ( 
.A1(n_6123),
.A2(n_6022),
.B(n_6010),
.Y(n_6475)
);

AND2x2_ASAP7_75t_L g6476 ( 
.A(n_6103),
.B(n_6018),
.Y(n_6476)
);

NOR2xp33_ASAP7_75t_SL g6477 ( 
.A(n_6292),
.B(n_4041),
.Y(n_6477)
);

AND2x2_ASAP7_75t_L g6478 ( 
.A(n_6103),
.B(n_6020),
.Y(n_6478)
);

NOR2x1_ASAP7_75t_R g6479 ( 
.A(n_6100),
.B(n_4324),
.Y(n_6479)
);

NAND2xp5_ASAP7_75t_L g6480 ( 
.A(n_6284),
.B(n_5945),
.Y(n_6480)
);

NOR2xp33_ASAP7_75t_L g6481 ( 
.A(n_6313),
.B(n_5783),
.Y(n_6481)
);

NOR3xp33_ASAP7_75t_L g6482 ( 
.A(n_6088),
.B(n_6022),
.C(n_6010),
.Y(n_6482)
);

AOI221xp5_ASAP7_75t_L g6483 ( 
.A1(n_6289),
.A2(n_6158),
.B1(n_6269),
.B2(n_6144),
.C(n_6224),
.Y(n_6483)
);

AND2x2_ASAP7_75t_L g6484 ( 
.A(n_6220),
.B(n_5785),
.Y(n_6484)
);

NAND2xp5_ASAP7_75t_L g6485 ( 
.A(n_6284),
.B(n_5947),
.Y(n_6485)
);

NAND2xp33_ASAP7_75t_SL g6486 ( 
.A(n_6314),
.B(n_5790),
.Y(n_6486)
);

OAI21xp5_ASAP7_75t_L g6487 ( 
.A1(n_6150),
.A2(n_5324),
.B(n_5243),
.Y(n_6487)
);

NOR2xp33_ASAP7_75t_L g6488 ( 
.A(n_6313),
.B(n_5804),
.Y(n_6488)
);

INVx2_ASAP7_75t_L g6489 ( 
.A(n_6302),
.Y(n_6489)
);

NOR3xp33_ASAP7_75t_L g6490 ( 
.A(n_6099),
.B(n_6042),
.C(n_6033),
.Y(n_6490)
);

AND2x2_ASAP7_75t_L g6491 ( 
.A(n_6328),
.B(n_5813),
.Y(n_6491)
);

NAND3xp33_ASAP7_75t_L g6492 ( 
.A(n_6333),
.B(n_5958),
.C(n_5952),
.Y(n_6492)
);

AND2x2_ASAP7_75t_L g6493 ( 
.A(n_6328),
.B(n_5815),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_6046),
.Y(n_6494)
);

AND2x2_ASAP7_75t_L g6495 ( 
.A(n_6227),
.B(n_5510),
.Y(n_6495)
);

OR2x6_ASAP7_75t_L g6496 ( 
.A(n_6112),
.B(n_6033),
.Y(n_6496)
);

NAND3xp33_ASAP7_75t_L g6497 ( 
.A(n_6333),
.B(n_5962),
.C(n_5960),
.Y(n_6497)
);

NAND4xp75_ASAP7_75t_L g6498 ( 
.A(n_6316),
.B(n_5812),
.C(n_5818),
.D(n_5811),
.Y(n_6498)
);

INVxp67_ASAP7_75t_SL g6499 ( 
.A(n_6302),
.Y(n_6499)
);

AND2x2_ASAP7_75t_L g6500 ( 
.A(n_6229),
.B(n_5515),
.Y(n_6500)
);

NAND3xp33_ASAP7_75t_L g6501 ( 
.A(n_6333),
.B(n_5991),
.C(n_5982),
.Y(n_6501)
);

NOR3xp33_ASAP7_75t_L g6502 ( 
.A(n_6104),
.B(n_6043),
.C(n_6042),
.Y(n_6502)
);

NOR3xp33_ASAP7_75t_L g6503 ( 
.A(n_6055),
.B(n_6043),
.C(n_5824),
.Y(n_6503)
);

NAND2xp5_ASAP7_75t_L g6504 ( 
.A(n_6237),
.B(n_5959),
.Y(n_6504)
);

AND2x2_ASAP7_75t_L g6505 ( 
.A(n_6112),
.B(n_5515),
.Y(n_6505)
);

AOI22xp33_ASAP7_75t_L g6506 ( 
.A1(n_6235),
.A2(n_5824),
.B1(n_5828),
.B2(n_5819),
.Y(n_6506)
);

INVx1_ASAP7_75t_L g6507 ( 
.A(n_6056),
.Y(n_6507)
);

NAND3xp33_ASAP7_75t_L g6508 ( 
.A(n_6058),
.B(n_5967),
.C(n_5966),
.Y(n_6508)
);

OA21x2_ASAP7_75t_L g6509 ( 
.A1(n_6159),
.A2(n_6327),
.B(n_6066),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_6063),
.Y(n_6510)
);

NAND2xp5_ASAP7_75t_L g6511 ( 
.A(n_6251),
.B(n_6165),
.Y(n_6511)
);

OR2x2_ASAP7_75t_L g6512 ( 
.A(n_6187),
.B(n_5981),
.Y(n_6512)
);

NAND2xp5_ASAP7_75t_L g6513 ( 
.A(n_6165),
.B(n_5993),
.Y(n_6513)
);

NAND2xp5_ASAP7_75t_L g6514 ( 
.A(n_6182),
.B(n_5600),
.Y(n_6514)
);

HB1xp67_ASAP7_75t_L g6515 ( 
.A(n_6152),
.Y(n_6515)
);

NAND3xp33_ASAP7_75t_L g6516 ( 
.A(n_6069),
.B(n_5828),
.C(n_5819),
.Y(n_6516)
);

AND2x2_ASAP7_75t_L g6517 ( 
.A(n_6186),
.B(n_6208),
.Y(n_6517)
);

AOI22xp5_ASAP7_75t_L g6518 ( 
.A1(n_6070),
.A2(n_5832),
.B1(n_5833),
.B2(n_5830),
.Y(n_6518)
);

NAND3xp33_ASAP7_75t_L g6519 ( 
.A(n_6151),
.B(n_5832),
.C(n_5830),
.Y(n_6519)
);

NOR3xp33_ASAP7_75t_L g6520 ( 
.A(n_6057),
.B(n_5833),
.C(n_5353),
.Y(n_6520)
);

AOI22xp33_ASAP7_75t_L g6521 ( 
.A1(n_6238),
.A2(n_6250),
.B1(n_6257),
.B2(n_6246),
.Y(n_6521)
);

NAND2xp5_ASAP7_75t_L g6522 ( 
.A(n_6182),
.B(n_5602),
.Y(n_6522)
);

INVx2_ASAP7_75t_L g6523 ( 
.A(n_6248),
.Y(n_6523)
);

INVx1_ASAP7_75t_L g6524 ( 
.A(n_6074),
.Y(n_6524)
);

NOR3xp33_ASAP7_75t_L g6525 ( 
.A(n_6061),
.B(n_5353),
.C(n_5349),
.Y(n_6525)
);

NAND2xp5_ASAP7_75t_SL g6526 ( 
.A(n_6186),
.B(n_5516),
.Y(n_6526)
);

NAND3xp33_ASAP7_75t_L g6527 ( 
.A(n_6151),
.B(n_5618),
.C(n_5613),
.Y(n_6527)
);

AND2x2_ASAP7_75t_L g6528 ( 
.A(n_6208),
.B(n_5516),
.Y(n_6528)
);

NOR2xp33_ASAP7_75t_L g6529 ( 
.A(n_6132),
.B(n_5521),
.Y(n_6529)
);

AND2x2_ASAP7_75t_L g6530 ( 
.A(n_6231),
.B(n_5521),
.Y(n_6530)
);

NOR3xp33_ASAP7_75t_L g6531 ( 
.A(n_6064),
.B(n_5618),
.C(n_5183),
.Y(n_6531)
);

OR2x2_ASAP7_75t_L g6532 ( 
.A(n_6160),
.B(n_5602),
.Y(n_6532)
);

INVx1_ASAP7_75t_L g6533 ( 
.A(n_6172),
.Y(n_6533)
);

NAND2xp5_ASAP7_75t_L g6534 ( 
.A(n_6248),
.B(n_5605),
.Y(n_6534)
);

AOI211xp5_ASAP7_75t_L g6535 ( 
.A1(n_6072),
.A2(n_5692),
.B(n_5691),
.C(n_5615),
.Y(n_6535)
);

INVx2_ASAP7_75t_L g6536 ( 
.A(n_6231),
.Y(n_6536)
);

INVx1_ASAP7_75t_L g6537 ( 
.A(n_6174),
.Y(n_6537)
);

INVx2_ASAP7_75t_SL g6538 ( 
.A(n_6132),
.Y(n_6538)
);

AND2x2_ASAP7_75t_L g6539 ( 
.A(n_6209),
.B(n_5522),
.Y(n_6539)
);

AOI22xp5_ASAP7_75t_L g6540 ( 
.A1(n_6175),
.A2(n_5626),
.B1(n_5632),
.B2(n_5623),
.Y(n_6540)
);

NAND2xp5_ASAP7_75t_SL g6541 ( 
.A(n_6135),
.B(n_5522),
.Y(n_6541)
);

INVx1_ASAP7_75t_L g6542 ( 
.A(n_6177),
.Y(n_6542)
);

AO21x2_ASAP7_75t_L g6543 ( 
.A1(n_6261),
.A2(n_5626),
.B(n_5623),
.Y(n_6543)
);

NAND2xp5_ASAP7_75t_L g6544 ( 
.A(n_6303),
.B(n_5605),
.Y(n_6544)
);

NOR3xp33_ASAP7_75t_SL g6545 ( 
.A(n_6252),
.B(n_6072),
.C(n_6236),
.Y(n_6545)
);

NOR2x1_ASAP7_75t_L g6546 ( 
.A(n_6176),
.B(n_5015),
.Y(n_6546)
);

OR2x2_ASAP7_75t_L g6547 ( 
.A(n_6160),
.B(n_5691),
.Y(n_6547)
);

AOI22xp33_ASAP7_75t_SL g6548 ( 
.A1(n_6178),
.A2(n_5208),
.B1(n_5170),
.B2(n_5151),
.Y(n_6548)
);

OAI211xp5_ASAP7_75t_L g6549 ( 
.A1(n_6106),
.A2(n_4970),
.B(n_4998),
.C(n_4986),
.Y(n_6549)
);

INVx1_ASAP7_75t_L g6550 ( 
.A(n_6184),
.Y(n_6550)
);

NAND3xp33_ASAP7_75t_L g6551 ( 
.A(n_6124),
.B(n_5121),
.C(n_5048),
.Y(n_6551)
);

NOR3xp33_ASAP7_75t_L g6552 ( 
.A(n_6108),
.B(n_5121),
.C(n_5048),
.Y(n_6552)
);

AND2x2_ASAP7_75t_L g6553 ( 
.A(n_6135),
.B(n_5530),
.Y(n_6553)
);

NOR2x1_ASAP7_75t_R g6554 ( 
.A(n_6176),
.B(n_4324),
.Y(n_6554)
);

OAI211xp5_ASAP7_75t_L g6555 ( 
.A1(n_6179),
.A2(n_5003),
.B(n_5121),
.C(n_5077),
.Y(n_6555)
);

AOI211xp5_ASAP7_75t_L g6556 ( 
.A1(n_6188),
.A2(n_5692),
.B(n_5616),
.C(n_5625),
.Y(n_6556)
);

AOI22xp33_ASAP7_75t_L g6557 ( 
.A1(n_6272),
.A2(n_5632),
.B1(n_5648),
.B2(n_5641),
.Y(n_6557)
);

AOI22xp33_ASAP7_75t_L g6558 ( 
.A1(n_6279),
.A2(n_5641),
.B1(n_5655),
.B2(n_5648),
.Y(n_6558)
);

NAND3xp33_ASAP7_75t_L g6559 ( 
.A(n_6206),
.B(n_5683),
.C(n_5681),
.Y(n_6559)
);

NOR3xp33_ASAP7_75t_L g6560 ( 
.A(n_6110),
.B(n_5077),
.C(n_5003),
.Y(n_6560)
);

NAND3xp33_ASAP7_75t_L g6561 ( 
.A(n_6210),
.B(n_6213),
.C(n_6252),
.Y(n_6561)
);

NAND2xp5_ASAP7_75t_L g6562 ( 
.A(n_6121),
.B(n_5530),
.Y(n_6562)
);

NAND4xp75_ASAP7_75t_L g6563 ( 
.A(n_6311),
.B(n_5616),
.C(n_5625),
.D(n_5615),
.Y(n_6563)
);

INVx2_ASAP7_75t_L g6564 ( 
.A(n_6140),
.Y(n_6564)
);

NAND3xp33_ASAP7_75t_L g6565 ( 
.A(n_6128),
.B(n_5687),
.C(n_5684),
.Y(n_6565)
);

AO21x2_ASAP7_75t_L g6566 ( 
.A1(n_6261),
.A2(n_5666),
.B(n_5655),
.Y(n_6566)
);

NAND3xp33_ASAP7_75t_L g6567 ( 
.A(n_6130),
.B(n_5687),
.C(n_5684),
.Y(n_6567)
);

AOI22xp5_ASAP7_75t_L g6568 ( 
.A1(n_6189),
.A2(n_5671),
.B1(n_5672),
.B2(n_5666),
.Y(n_6568)
);

AOI221xp5_ASAP7_75t_L g6569 ( 
.A1(n_6193),
.A2(n_5672),
.B1(n_5671),
.B2(n_5124),
.C(n_5143),
.Y(n_6569)
);

AOI221xp5_ASAP7_75t_L g6570 ( 
.A1(n_6195),
.A2(n_5124),
.B1(n_5143),
.B2(n_5077),
.C(n_5003),
.Y(n_6570)
);

AND2x2_ASAP7_75t_L g6571 ( 
.A(n_6095),
.B(n_6116),
.Y(n_6571)
);

INVx2_ASAP7_75t_L g6572 ( 
.A(n_6243),
.Y(n_6572)
);

AND2x2_ASAP7_75t_L g6573 ( 
.A(n_6162),
.B(n_5533),
.Y(n_6573)
);

HB1xp67_ASAP7_75t_L g6574 ( 
.A(n_6169),
.Y(n_6574)
);

AND2x4_ASAP7_75t_L g6575 ( 
.A(n_6267),
.B(n_5533),
.Y(n_6575)
);

HB1xp67_ASAP7_75t_L g6576 ( 
.A(n_6171),
.Y(n_6576)
);

AND2x2_ASAP7_75t_L g6577 ( 
.A(n_6190),
.B(n_5534),
.Y(n_6577)
);

NOR3xp33_ASAP7_75t_L g6578 ( 
.A(n_6075),
.B(n_5183),
.C(n_5143),
.Y(n_6578)
);

AND2x4_ASAP7_75t_L g6579 ( 
.A(n_6268),
.B(n_5534),
.Y(n_6579)
);

NAND3xp33_ASAP7_75t_L g6580 ( 
.A(n_6271),
.B(n_6282),
.C(n_6131),
.Y(n_6580)
);

INVxp67_ASAP7_75t_SL g6581 ( 
.A(n_6243),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_6205),
.Y(n_6582)
);

AOI22xp33_ASAP7_75t_L g6583 ( 
.A1(n_6280),
.A2(n_5157),
.B1(n_5176),
.B2(n_4949),
.Y(n_6583)
);

AND2x2_ASAP7_75t_L g6584 ( 
.A(n_6198),
.B(n_5535),
.Y(n_6584)
);

AND2x2_ASAP7_75t_L g6585 ( 
.A(n_6335),
.B(n_5535),
.Y(n_6585)
);

OR2x2_ASAP7_75t_L g6586 ( 
.A(n_6166),
.B(n_5537),
.Y(n_6586)
);

OA211x2_ASAP7_75t_L g6587 ( 
.A1(n_6136),
.A2(n_4392),
.B(n_4207),
.C(n_4255),
.Y(n_6587)
);

AOI22xp5_ASAP7_75t_L g6588 ( 
.A1(n_6218),
.A2(n_5124),
.B1(n_5160),
.B2(n_5153),
.Y(n_6588)
);

NAND2xp5_ASAP7_75t_L g6589 ( 
.A(n_6317),
.B(n_5537),
.Y(n_6589)
);

OR2x2_ASAP7_75t_L g6590 ( 
.A(n_6204),
.B(n_5539),
.Y(n_6590)
);

NOR3xp33_ASAP7_75t_L g6591 ( 
.A(n_6107),
.B(n_5207),
.C(n_5160),
.Y(n_6591)
);

NAND4xp75_ASAP7_75t_L g6592 ( 
.A(n_6120),
.B(n_6225),
.C(n_6223),
.D(n_6133),
.Y(n_6592)
);

AND2x2_ASAP7_75t_L g6593 ( 
.A(n_6312),
.B(n_6262),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_6475),
.Y(n_6594)
);

AND2x2_ASAP7_75t_L g6595 ( 
.A(n_6387),
.B(n_6297),
.Y(n_6595)
);

NAND4xp25_ASAP7_75t_L g6596 ( 
.A(n_6409),
.B(n_6126),
.C(n_6143),
.D(n_6137),
.Y(n_6596)
);

NAND2xp5_ASAP7_75t_SL g6597 ( 
.A(n_6376),
.B(n_6243),
.Y(n_6597)
);

OAI211xp5_ASAP7_75t_L g6598 ( 
.A1(n_6352),
.A2(n_6161),
.B(n_6156),
.C(n_6183),
.Y(n_6598)
);

AOI221xp5_ASAP7_75t_L g6599 ( 
.A1(n_6483),
.A2(n_6202),
.B1(n_6265),
.B2(n_6304),
.C(n_6285),
.Y(n_6599)
);

INVx1_ASAP7_75t_SL g6600 ( 
.A(n_6355),
.Y(n_6600)
);

AND2x2_ASAP7_75t_L g6601 ( 
.A(n_6403),
.B(n_6239),
.Y(n_6601)
);

OAI33xp33_ASAP7_75t_L g6602 ( 
.A1(n_6414),
.A2(n_6202),
.A3(n_6318),
.B1(n_6196),
.B2(n_6200),
.B3(n_6204),
.Y(n_6602)
);

AND2x2_ASAP7_75t_L g6603 ( 
.A(n_6388),
.B(n_6239),
.Y(n_6603)
);

OR2x2_ASAP7_75t_L g6604 ( 
.A(n_6375),
.B(n_6196),
.Y(n_6604)
);

INVx2_ASAP7_75t_L g6605 ( 
.A(n_6353),
.Y(n_6605)
);

INVxp67_ASAP7_75t_SL g6606 ( 
.A(n_6382),
.Y(n_6606)
);

OR2x2_ASAP7_75t_L g6607 ( 
.A(n_6402),
.B(n_6200),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6475),
.Y(n_6608)
);

AND2x2_ASAP7_75t_L g6609 ( 
.A(n_6399),
.B(n_6060),
.Y(n_6609)
);

INVx1_ASAP7_75t_SL g6610 ( 
.A(n_6355),
.Y(n_6610)
);

OAI31xp33_ASAP7_75t_L g6611 ( 
.A1(n_6397),
.A2(n_6322),
.A3(n_6325),
.B(n_6321),
.Y(n_6611)
);

AOI32xp33_ASAP7_75t_L g6612 ( 
.A1(n_6391),
.A2(n_6266),
.A3(n_6226),
.B1(n_6221),
.B2(n_6217),
.Y(n_6612)
);

BUFx2_ASAP7_75t_L g6613 ( 
.A(n_6404),
.Y(n_6613)
);

INVx1_ASAP7_75t_L g6614 ( 
.A(n_6369),
.Y(n_6614)
);

OR2x2_ASAP7_75t_L g6615 ( 
.A(n_6366),
.B(n_6217),
.Y(n_6615)
);

INVx1_ASAP7_75t_SL g6616 ( 
.A(n_6369),
.Y(n_6616)
);

NAND2x1_ASAP7_75t_SL g6617 ( 
.A(n_6343),
.B(n_6287),
.Y(n_6617)
);

OR2x2_ASAP7_75t_L g6618 ( 
.A(n_6357),
.B(n_6221),
.Y(n_6618)
);

NOR2xp33_ASAP7_75t_L g6619 ( 
.A(n_6464),
.B(n_6219),
.Y(n_6619)
);

AND2x2_ASAP7_75t_SL g6620 ( 
.A(n_6410),
.B(n_6219),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_6425),
.Y(n_6621)
);

AND2x2_ASAP7_75t_L g6622 ( 
.A(n_6354),
.B(n_6060),
.Y(n_6622)
);

OAI33xp33_ASAP7_75t_L g6623 ( 
.A1(n_6473),
.A2(n_6226),
.A3(n_6336),
.B1(n_6332),
.B2(n_6329),
.B3(n_6245),
.Y(n_6623)
);

INVx1_ASAP7_75t_L g6624 ( 
.A(n_6425),
.Y(n_6624)
);

NOR2xp33_ASAP7_75t_L g6625 ( 
.A(n_6344),
.B(n_6062),
.Y(n_6625)
);

AOI222xp33_ASAP7_75t_L g6626 ( 
.A1(n_6383),
.A2(n_6294),
.B1(n_6281),
.B2(n_6276),
.C1(n_6270),
.C2(n_6298),
.Y(n_6626)
);

AND2x2_ASAP7_75t_L g6627 ( 
.A(n_6419),
.B(n_6405),
.Y(n_6627)
);

AND2x2_ASAP7_75t_L g6628 ( 
.A(n_6422),
.B(n_6060),
.Y(n_6628)
);

NOR2xp33_ASAP7_75t_L g6629 ( 
.A(n_6345),
.B(n_6062),
.Y(n_6629)
);

HB1xp67_ASAP7_75t_L g6630 ( 
.A(n_6472),
.Y(n_6630)
);

INVx1_ASAP7_75t_L g6631 ( 
.A(n_6515),
.Y(n_6631)
);

INVx2_ASAP7_75t_L g6632 ( 
.A(n_6353),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_6574),
.Y(n_6633)
);

AND2x2_ASAP7_75t_L g6634 ( 
.A(n_6424),
.B(n_6233),
.Y(n_6634)
);

HB1xp67_ASAP7_75t_L g6635 ( 
.A(n_6349),
.Y(n_6635)
);

AOI33xp33_ASAP7_75t_L g6636 ( 
.A1(n_6450),
.A2(n_6242),
.A3(n_6260),
.B1(n_6263),
.B2(n_6247),
.B3(n_6288),
.Y(n_6636)
);

INVx2_ASAP7_75t_L g6637 ( 
.A(n_6404),
.Y(n_6637)
);

OAI21xp33_ASAP7_75t_L g6638 ( 
.A1(n_6545),
.A2(n_6253),
.B(n_6293),
.Y(n_6638)
);

INVx2_ASAP7_75t_SL g6639 ( 
.A(n_6376),
.Y(n_6639)
);

INVx1_ASAP7_75t_L g6640 ( 
.A(n_6576),
.Y(n_6640)
);

NAND2xp5_ASAP7_75t_L g6641 ( 
.A(n_6427),
.B(n_6340),
.Y(n_6641)
);

AOI22xp5_ASAP7_75t_L g6642 ( 
.A1(n_6426),
.A2(n_6290),
.B1(n_6264),
.B2(n_6277),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6384),
.Y(n_6643)
);

INVx1_ASAP7_75t_L g6644 ( 
.A(n_6394),
.Y(n_6644)
);

HB1xp67_ASAP7_75t_L g6645 ( 
.A(n_6349),
.Y(n_6645)
);

INVx2_ASAP7_75t_L g6646 ( 
.A(n_6456),
.Y(n_6646)
);

AND2x2_ASAP7_75t_L g6647 ( 
.A(n_6364),
.B(n_5539),
.Y(n_6647)
);

INVx1_ASAP7_75t_L g6648 ( 
.A(n_6499),
.Y(n_6648)
);

INVx2_ASAP7_75t_L g6649 ( 
.A(n_6456),
.Y(n_6649)
);

AND2x2_ASAP7_75t_L g6650 ( 
.A(n_6476),
.B(n_5556),
.Y(n_6650)
);

INVx1_ASAP7_75t_L g6651 ( 
.A(n_6351),
.Y(n_6651)
);

AND2x4_ASAP7_75t_L g6652 ( 
.A(n_6517),
.B(n_6295),
.Y(n_6652)
);

OR2x2_ASAP7_75t_L g6653 ( 
.A(n_6532),
.B(n_6270),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_6437),
.Y(n_6654)
);

NAND2xp5_ASAP7_75t_L g6655 ( 
.A(n_6495),
.B(n_6296),
.Y(n_6655)
);

OR2x2_ASAP7_75t_L g6656 ( 
.A(n_6421),
.B(n_6276),
.Y(n_6656)
);

NAND2xp5_ASAP7_75t_L g6657 ( 
.A(n_6500),
.B(n_6306),
.Y(n_6657)
);

NAND2xp5_ASAP7_75t_L g6658 ( 
.A(n_6585),
.B(n_6307),
.Y(n_6658)
);

INVx2_ASAP7_75t_L g6659 ( 
.A(n_6484),
.Y(n_6659)
);

INVx2_ASAP7_75t_L g6660 ( 
.A(n_6491),
.Y(n_6660)
);

INVx1_ASAP7_75t_L g6661 ( 
.A(n_6429),
.Y(n_6661)
);

AND2x2_ASAP7_75t_L g6662 ( 
.A(n_6478),
.B(n_5556),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_6449),
.Y(n_6663)
);

INVx1_ASAP7_75t_L g6664 ( 
.A(n_6451),
.Y(n_6664)
);

INVx2_ASAP7_75t_L g6665 ( 
.A(n_6493),
.Y(n_6665)
);

OAI22xp5_ASAP7_75t_L g6666 ( 
.A1(n_6371),
.A2(n_6244),
.B1(n_6256),
.B2(n_5564),
.Y(n_6666)
);

AOI31xp33_ASAP7_75t_L g6667 ( 
.A1(n_6581),
.A2(n_6305),
.A3(n_6326),
.B(n_6298),
.Y(n_6667)
);

INVx1_ASAP7_75t_L g6668 ( 
.A(n_6348),
.Y(n_6668)
);

AOI22xp5_ASAP7_75t_L g6669 ( 
.A1(n_6498),
.A2(n_6290),
.B1(n_6264),
.B2(n_6277),
.Y(n_6669)
);

OAI21xp5_ASAP7_75t_SL g6670 ( 
.A1(n_6359),
.A2(n_6253),
.B(n_6330),
.Y(n_6670)
);

AND3x2_ASAP7_75t_L g6671 ( 
.A(n_6466),
.B(n_5325),
.C(n_5576),
.Y(n_6671)
);

INVx2_ASAP7_75t_L g6672 ( 
.A(n_6447),
.Y(n_6672)
);

NOR2xp33_ASAP7_75t_R g6673 ( 
.A(n_6486),
.B(n_4287),
.Y(n_6673)
);

INVx2_ASAP7_75t_L g6674 ( 
.A(n_6442),
.Y(n_6674)
);

OAI31xp33_ASAP7_75t_L g6675 ( 
.A1(n_6358),
.A2(n_6293),
.A3(n_6326),
.B(n_6305),
.Y(n_6675)
);

INVx2_ASAP7_75t_L g6676 ( 
.A(n_6390),
.Y(n_6676)
);

NAND2xp5_ASAP7_75t_L g6677 ( 
.A(n_6474),
.B(n_6575),
.Y(n_6677)
);

OR2x2_ASAP7_75t_L g6678 ( 
.A(n_6547),
.B(n_5573),
.Y(n_6678)
);

BUFx3_ASAP7_75t_L g6679 ( 
.A(n_6538),
.Y(n_6679)
);

AND2x2_ASAP7_75t_L g6680 ( 
.A(n_6465),
.B(n_5573),
.Y(n_6680)
);

OR2x2_ASAP7_75t_L g6681 ( 
.A(n_6544),
.B(n_5560),
.Y(n_6681)
);

INVx2_ASAP7_75t_L g6682 ( 
.A(n_6553),
.Y(n_6682)
);

OAI21xp5_ASAP7_75t_SL g6683 ( 
.A1(n_6380),
.A2(n_5576),
.B(n_5160),
.Y(n_6683)
);

AND2x2_ASAP7_75t_L g6684 ( 
.A(n_6528),
.B(n_5560),
.Y(n_6684)
);

NOR2xp67_ASAP7_75t_L g6685 ( 
.A(n_6580),
.B(n_5690),
.Y(n_6685)
);

NOR2xp33_ASAP7_75t_L g6686 ( 
.A(n_6347),
.B(n_5564),
.Y(n_6686)
);

AOI222xp33_ASAP7_75t_L g6687 ( 
.A1(n_6440),
.A2(n_4957),
.B1(n_4949),
.B2(n_4953),
.C1(n_5069),
.C2(n_5060),
.Y(n_6687)
);

AND2x2_ASAP7_75t_L g6688 ( 
.A(n_6530),
.B(n_5565),
.Y(n_6688)
);

INVx1_ASAP7_75t_L g6689 ( 
.A(n_6480),
.Y(n_6689)
);

AND2x2_ASAP7_75t_L g6690 ( 
.A(n_6381),
.B(n_5565),
.Y(n_6690)
);

AOI211x1_ASAP7_75t_L g6691 ( 
.A1(n_6400),
.A2(n_5569),
.B(n_5150),
.C(n_5156),
.Y(n_6691)
);

INVx4_ASAP7_75t_L g6692 ( 
.A(n_6362),
.Y(n_6692)
);

AND2x2_ASAP7_75t_L g6693 ( 
.A(n_6386),
.B(n_5569),
.Y(n_6693)
);

AND2x2_ASAP7_75t_SL g6694 ( 
.A(n_6470),
.B(n_4509),
.Y(n_6694)
);

INVx2_ASAP7_75t_L g6695 ( 
.A(n_6418),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_6485),
.Y(n_6696)
);

AOI221xp5_ASAP7_75t_L g6697 ( 
.A1(n_6462),
.A2(n_6185),
.B1(n_5187),
.B2(n_5198),
.C(n_5183),
.Y(n_6697)
);

AND2x2_ASAP7_75t_L g6698 ( 
.A(n_6571),
.B(n_6214),
.Y(n_6698)
);

OAI22xp5_ASAP7_75t_L g6699 ( 
.A1(n_6365),
.A2(n_5335),
.B1(n_5290),
.B2(n_5267),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_6360),
.Y(n_6700)
);

INVx1_ASAP7_75t_L g6701 ( 
.A(n_6363),
.Y(n_6701)
);

NOR2xp33_ASAP7_75t_L g6702 ( 
.A(n_6435),
.B(n_6309),
.Y(n_6702)
);

OAI22xp5_ASAP7_75t_L g6703 ( 
.A1(n_6367),
.A2(n_5335),
.B1(n_5290),
.B2(n_5267),
.Y(n_6703)
);

AOI21xp5_ASAP7_75t_L g6704 ( 
.A1(n_6526),
.A2(n_6168),
.B(n_6134),
.Y(n_6704)
);

HB1xp67_ASAP7_75t_L g6705 ( 
.A(n_6509),
.Y(n_6705)
);

INVx1_ASAP7_75t_L g6706 ( 
.A(n_6368),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_6379),
.Y(n_6707)
);

OAI221xp5_ASAP7_75t_L g6708 ( 
.A1(n_6446),
.A2(n_6309),
.B1(n_5198),
.B2(n_5206),
.C(n_5187),
.Y(n_6708)
);

OR2x2_ASAP7_75t_L g6709 ( 
.A(n_6350),
.B(n_5142),
.Y(n_6709)
);

HB1xp67_ASAP7_75t_L g6710 ( 
.A(n_6509),
.Y(n_6710)
);

O2A1O1Ixp33_ASAP7_75t_SL g6711 ( 
.A1(n_6541),
.A2(n_5697),
.B(n_5690),
.C(n_5187),
.Y(n_6711)
);

AND2x2_ASAP7_75t_L g6712 ( 
.A(n_6539),
.B(n_5697),
.Y(n_6712)
);

OAI33xp33_ASAP7_75t_L g6713 ( 
.A1(n_6516),
.A2(n_5150),
.A3(n_5156),
.B1(n_5161),
.B2(n_5159),
.B3(n_5142),
.Y(n_6713)
);

AND2x2_ASAP7_75t_L g6714 ( 
.A(n_6573),
.B(n_4287),
.Y(n_6714)
);

AND2x2_ASAP7_75t_L g6715 ( 
.A(n_6577),
.B(n_4287),
.Y(n_6715)
);

NOR2xp33_ASAP7_75t_L g6716 ( 
.A(n_6479),
.B(n_6309),
.Y(n_6716)
);

INVx1_ASAP7_75t_L g6717 ( 
.A(n_6342),
.Y(n_6717)
);

AND2x4_ASAP7_75t_L g6718 ( 
.A(n_6536),
.B(n_5347),
.Y(n_6718)
);

OAI31xp33_ASAP7_75t_L g6719 ( 
.A1(n_6373),
.A2(n_5347),
.A3(n_5198),
.B(n_5206),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6356),
.Y(n_6720)
);

OAI221xp5_ASAP7_75t_L g6721 ( 
.A1(n_6548),
.A2(n_5207),
.B1(n_5277),
.B2(n_5206),
.C(n_5153),
.Y(n_6721)
);

INVx2_ASAP7_75t_L g6722 ( 
.A(n_6575),
.Y(n_6722)
);

INVx1_ASAP7_75t_L g6723 ( 
.A(n_6346),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_6377),
.Y(n_6724)
);

NOR2xp33_ASAP7_75t_SL g6725 ( 
.A(n_6592),
.B(n_4041),
.Y(n_6725)
);

OR2x2_ASAP7_75t_L g6726 ( 
.A(n_6443),
.B(n_5159),
.Y(n_6726)
);

INVx1_ASAP7_75t_L g6727 ( 
.A(n_6423),
.Y(n_6727)
);

AND2x2_ASAP7_75t_L g6728 ( 
.A(n_6584),
.B(n_4306),
.Y(n_6728)
);

NAND3xp33_ASAP7_75t_SL g6729 ( 
.A(n_6389),
.B(n_6417),
.C(n_6407),
.Y(n_6729)
);

OAI33xp33_ASAP7_75t_L g6730 ( 
.A1(n_6511),
.A2(n_5175),
.A3(n_5180),
.B1(n_5192),
.B2(n_5191),
.B3(n_5161),
.Y(n_6730)
);

OAI33xp33_ASAP7_75t_L g6731 ( 
.A1(n_6458),
.A2(n_6504),
.A3(n_6519),
.B1(n_6408),
.B2(n_6385),
.B3(n_6412),
.Y(n_6731)
);

OAI33xp33_ASAP7_75t_L g6732 ( 
.A1(n_6458),
.A2(n_6519),
.A3(n_6406),
.B1(n_6432),
.B2(n_6396),
.B3(n_6513),
.Y(n_6732)
);

INVx1_ASAP7_75t_L g6733 ( 
.A(n_6439),
.Y(n_6733)
);

NAND2xp5_ASAP7_75t_L g6734 ( 
.A(n_6579),
.B(n_5175),
.Y(n_6734)
);

AOI222xp33_ASAP7_75t_L g6735 ( 
.A1(n_6393),
.A2(n_5060),
.B1(n_5096),
.B2(n_5106),
.C1(n_5105),
.C2(n_5069),
.Y(n_6735)
);

INVx2_ASAP7_75t_L g6736 ( 
.A(n_6579),
.Y(n_6736)
);

OAI31xp33_ASAP7_75t_L g6737 ( 
.A1(n_6455),
.A2(n_5207),
.A3(n_5277),
.B(n_5153),
.Y(n_6737)
);

AOI211xp5_ASAP7_75t_L g6738 ( 
.A1(n_6372),
.A2(n_5277),
.B(n_5347),
.C(n_5289),
.Y(n_6738)
);

INVx2_ASAP7_75t_L g6739 ( 
.A(n_6564),
.Y(n_6739)
);

OAI31xp33_ASAP7_75t_SL g6740 ( 
.A1(n_6546),
.A2(n_5090),
.A3(n_5220),
.B(n_5177),
.Y(n_6740)
);

INVx2_ASAP7_75t_SL g6741 ( 
.A(n_6505),
.Y(n_6741)
);

INVx3_ASAP7_75t_L g6742 ( 
.A(n_6496),
.Y(n_6742)
);

AND2x2_ASAP7_75t_L g6743 ( 
.A(n_6593),
.B(n_4306),
.Y(n_6743)
);

NAND2xp5_ASAP7_75t_L g6744 ( 
.A(n_6411),
.B(n_5180),
.Y(n_6744)
);

INVxp67_ASAP7_75t_SL g6745 ( 
.A(n_6479),
.Y(n_6745)
);

NAND3xp33_ASAP7_75t_L g6746 ( 
.A(n_6436),
.B(n_6148),
.C(n_6203),
.Y(n_6746)
);

INVx2_ASAP7_75t_L g6747 ( 
.A(n_6496),
.Y(n_6747)
);

AND2x4_ASAP7_75t_L g6748 ( 
.A(n_6523),
.B(n_5289),
.Y(n_6748)
);

OR2x2_ASAP7_75t_L g6749 ( 
.A(n_6445),
.B(n_5191),
.Y(n_6749)
);

INVx1_ASAP7_75t_L g6750 ( 
.A(n_6590),
.Y(n_6750)
);

INVxp67_ASAP7_75t_L g6751 ( 
.A(n_6554),
.Y(n_6751)
);

AND2x4_ASAP7_75t_L g6752 ( 
.A(n_6489),
.B(n_5289),
.Y(n_6752)
);

AND2x2_ASAP7_75t_L g6753 ( 
.A(n_6481),
.B(n_6488),
.Y(n_6753)
);

OAI221xp5_ASAP7_75t_SL g6754 ( 
.A1(n_6535),
.A2(n_5249),
.B1(n_5252),
.B2(n_5232),
.C(n_5034),
.Y(n_6754)
);

BUFx2_ASAP7_75t_L g6755 ( 
.A(n_6496),
.Y(n_6755)
);

AND2x2_ASAP7_75t_L g6756 ( 
.A(n_6529),
.B(n_4306),
.Y(n_6756)
);

NAND2xp5_ASAP7_75t_L g6757 ( 
.A(n_6398),
.B(n_5192),
.Y(n_6757)
);

OAI22xp33_ASAP7_75t_L g6758 ( 
.A1(n_6428),
.A2(n_5252),
.B1(n_5249),
.B2(n_5034),
.Y(n_6758)
);

INVx2_ASAP7_75t_L g6759 ( 
.A(n_6461),
.Y(n_6759)
);

AND4x1_ASAP7_75t_L g6760 ( 
.A(n_6370),
.B(n_4285),
.C(n_3922),
.D(n_3936),
.Y(n_6760)
);

AND2x2_ASAP7_75t_L g6761 ( 
.A(n_6448),
.B(n_4324),
.Y(n_6761)
);

INVx1_ASAP7_75t_L g6762 ( 
.A(n_6514),
.Y(n_6762)
);

AND2x2_ASAP7_75t_L g6763 ( 
.A(n_6361),
.B(n_4336),
.Y(n_6763)
);

INVx1_ASAP7_75t_L g6764 ( 
.A(n_6522),
.Y(n_6764)
);

OAI221xp5_ASAP7_75t_L g6765 ( 
.A1(n_6395),
.A2(n_5208),
.B1(n_5170),
.B2(n_5232),
.C(n_5034),
.Y(n_6765)
);

OR2x2_ASAP7_75t_L g6766 ( 
.A(n_6534),
.B(n_5203),
.Y(n_6766)
);

NAND2xp5_ASAP7_75t_L g6767 ( 
.A(n_6572),
.B(n_5203),
.Y(n_6767)
);

HB1xp67_ASAP7_75t_L g6768 ( 
.A(n_6452),
.Y(n_6768)
);

INVx1_ASAP7_75t_L g6769 ( 
.A(n_6457),
.Y(n_6769)
);

OR2x2_ASAP7_75t_L g6770 ( 
.A(n_6586),
.B(n_5215),
.Y(n_6770)
);

AOI31xp33_ASAP7_75t_L g6771 ( 
.A1(n_6401),
.A2(n_4921),
.A3(n_3998),
.B(n_4078),
.Y(n_6771)
);

NAND3xp33_ASAP7_75t_L g6772 ( 
.A(n_6454),
.B(n_6148),
.C(n_6203),
.Y(n_6772)
);

AND2x2_ASAP7_75t_L g6773 ( 
.A(n_6535),
.B(n_4336),
.Y(n_6773)
);

INVx2_ASAP7_75t_L g6774 ( 
.A(n_6453),
.Y(n_6774)
);

INVx1_ASAP7_75t_L g6775 ( 
.A(n_6468),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_6471),
.Y(n_6776)
);

NOR2xp67_ASAP7_75t_L g6777 ( 
.A(n_6561),
.B(n_5212),
.Y(n_6777)
);

HB1xp67_ASAP7_75t_L g6778 ( 
.A(n_6562),
.Y(n_6778)
);

INVx2_ASAP7_75t_SL g6779 ( 
.A(n_6434),
.Y(n_6779)
);

AND2x2_ASAP7_75t_L g6780 ( 
.A(n_6556),
.B(n_4336),
.Y(n_6780)
);

AOI21xp5_ASAP7_75t_L g6781 ( 
.A1(n_6460),
.A2(n_6185),
.B(n_6211),
.Y(n_6781)
);

INVx1_ASAP7_75t_L g6782 ( 
.A(n_6512),
.Y(n_6782)
);

AND2x2_ASAP7_75t_L g6783 ( 
.A(n_6556),
.B(n_4413),
.Y(n_6783)
);

NAND2xp5_ASAP7_75t_L g6784 ( 
.A(n_6380),
.B(n_6521),
.Y(n_6784)
);

INVx1_ASAP7_75t_L g6785 ( 
.A(n_6527),
.Y(n_6785)
);

BUFx3_ASAP7_75t_L g6786 ( 
.A(n_6444),
.Y(n_6786)
);

INVx2_ASAP7_75t_SL g6787 ( 
.A(n_6589),
.Y(n_6787)
);

NOR2xp33_ASAP7_75t_L g6788 ( 
.A(n_6554),
.B(n_4413),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_6527),
.Y(n_6789)
);

INVx1_ASAP7_75t_L g6790 ( 
.A(n_6518),
.Y(n_6790)
);

AOI22xp33_ASAP7_75t_L g6791 ( 
.A1(n_6520),
.A2(n_6211),
.B1(n_6249),
.B2(n_5157),
.Y(n_6791)
);

HB1xp67_ASAP7_75t_L g6792 ( 
.A(n_6374),
.Y(n_6792)
);

INVx1_ASAP7_75t_L g6793 ( 
.A(n_6518),
.Y(n_6793)
);

INVx1_ASAP7_75t_L g6794 ( 
.A(n_6428),
.Y(n_6794)
);

NAND2x1_ASAP7_75t_SL g6795 ( 
.A(n_6459),
.B(n_6438),
.Y(n_6795)
);

AND2x2_ASAP7_75t_L g6796 ( 
.A(n_6563),
.B(n_4413),
.Y(n_6796)
);

NAND4xp25_ASAP7_75t_SL g6797 ( 
.A(n_6378),
.B(n_4863),
.C(n_4865),
.D(n_4860),
.Y(n_6797)
);

AND2x4_ASAP7_75t_L g6798 ( 
.A(n_6392),
.B(n_4856),
.Y(n_6798)
);

AOI221xp5_ASAP7_75t_L g6799 ( 
.A1(n_6525),
.A2(n_4957),
.B1(n_4953),
.B2(n_4941),
.C(n_5096),
.Y(n_6799)
);

NAND2xp5_ASAP7_75t_L g6800 ( 
.A(n_6469),
.B(n_5212),
.Y(n_6800)
);

INVx1_ASAP7_75t_L g6801 ( 
.A(n_6467),
.Y(n_6801)
);

AND2x2_ASAP7_75t_L g6802 ( 
.A(n_6477),
.B(n_4807),
.Y(n_6802)
);

AND2x2_ASAP7_75t_L g6803 ( 
.A(n_6441),
.B(n_4807),
.Y(n_6803)
);

NAND2xp5_ASAP7_75t_L g6804 ( 
.A(n_6482),
.B(n_6490),
.Y(n_6804)
);

AND2x2_ASAP7_75t_L g6805 ( 
.A(n_6494),
.B(n_4346),
.Y(n_6805)
);

INVx2_ASAP7_75t_L g6806 ( 
.A(n_6533),
.Y(n_6806)
);

INVx2_ASAP7_75t_L g6807 ( 
.A(n_6537),
.Y(n_6807)
);

INVx1_ASAP7_75t_L g6808 ( 
.A(n_6507),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_6510),
.Y(n_6809)
);

INVx1_ASAP7_75t_L g6810 ( 
.A(n_6524),
.Y(n_6810)
);

OAI31xp33_ASAP7_75t_L g6811 ( 
.A1(n_6413),
.A2(n_4176),
.A3(n_4179),
.B(n_4102),
.Y(n_6811)
);

OAI221xp5_ASAP7_75t_L g6812 ( 
.A1(n_6433),
.A2(n_6502),
.B1(n_6503),
.B2(n_6583),
.C(n_6506),
.Y(n_6812)
);

OAI321xp33_ASAP7_75t_L g6813 ( 
.A1(n_6459),
.A2(n_5290),
.A3(n_5267),
.B1(n_6249),
.B2(n_5232),
.C(n_5034),
.Y(n_6813)
);

BUFx2_ASAP7_75t_L g6814 ( 
.A(n_6487),
.Y(n_6814)
);

INVx1_ASAP7_75t_L g6815 ( 
.A(n_6540),
.Y(n_6815)
);

AND2x2_ASAP7_75t_L g6816 ( 
.A(n_6542),
.B(n_4363),
.Y(n_6816)
);

NAND2xp5_ASAP7_75t_L g6817 ( 
.A(n_6460),
.B(n_5215),
.Y(n_6817)
);

AND2x2_ASAP7_75t_L g6818 ( 
.A(n_6550),
.B(n_4363),
.Y(n_6818)
);

HB1xp67_ASAP7_75t_L g6819 ( 
.A(n_6582),
.Y(n_6819)
);

AND2x2_ASAP7_75t_L g6820 ( 
.A(n_6552),
.B(n_4218),
.Y(n_6820)
);

NAND2xp5_ASAP7_75t_L g6821 ( 
.A(n_6415),
.B(n_5219),
.Y(n_6821)
);

AOI31xp33_ASAP7_75t_L g6822 ( 
.A1(n_6416),
.A2(n_3998),
.A3(n_3991),
.B(n_4295),
.Y(n_6822)
);

AND2x4_ASAP7_75t_L g6823 ( 
.A(n_6613),
.B(n_6430),
.Y(n_6823)
);

INVx1_ASAP7_75t_L g6824 ( 
.A(n_6635),
.Y(n_6824)
);

AOI22xp33_ASAP7_75t_L g6825 ( 
.A1(n_6794),
.A2(n_6566),
.B1(n_6543),
.B2(n_6558),
.Y(n_6825)
);

OR2x2_ASAP7_75t_L g6826 ( 
.A(n_6618),
.B(n_6431),
.Y(n_6826)
);

INVx2_ASAP7_75t_SL g6827 ( 
.A(n_6617),
.Y(n_6827)
);

INVx1_ASAP7_75t_L g6828 ( 
.A(n_6645),
.Y(n_6828)
);

AND2x2_ASAP7_75t_L g6829 ( 
.A(n_6627),
.B(n_6560),
.Y(n_6829)
);

OR2x2_ASAP7_75t_L g6830 ( 
.A(n_6607),
.B(n_6508),
.Y(n_6830)
);

INVx2_ASAP7_75t_L g6831 ( 
.A(n_6795),
.Y(n_6831)
);

INVx2_ASAP7_75t_L g6832 ( 
.A(n_6679),
.Y(n_6832)
);

INVxp67_ASAP7_75t_L g6833 ( 
.A(n_6755),
.Y(n_6833)
);

OAI21xp33_ASAP7_75t_L g6834 ( 
.A1(n_6625),
.A2(n_6567),
.B(n_6565),
.Y(n_6834)
);

AND2x2_ASAP7_75t_L g6835 ( 
.A(n_6647),
.B(n_6492),
.Y(n_6835)
);

NAND2xp5_ASAP7_75t_L g6836 ( 
.A(n_6606),
.B(n_6497),
.Y(n_6836)
);

INVx1_ASAP7_75t_L g6837 ( 
.A(n_6594),
.Y(n_6837)
);

AND2x2_ASAP7_75t_L g6838 ( 
.A(n_6690),
.B(n_6501),
.Y(n_6838)
);

OR2x2_ASAP7_75t_L g6839 ( 
.A(n_6615),
.B(n_6559),
.Y(n_6839)
);

AND2x2_ASAP7_75t_L g6840 ( 
.A(n_6693),
.B(n_6591),
.Y(n_6840)
);

OR2x2_ASAP7_75t_L g6841 ( 
.A(n_6604),
.B(n_6551),
.Y(n_6841)
);

INVx1_ASAP7_75t_L g6842 ( 
.A(n_6705),
.Y(n_6842)
);

INVx2_ASAP7_75t_L g6843 ( 
.A(n_6742),
.Y(n_6843)
);

AND2x2_ASAP7_75t_L g6844 ( 
.A(n_6609),
.B(n_6578),
.Y(n_6844)
);

OR2x6_ASAP7_75t_L g6845 ( 
.A(n_6739),
.B(n_5249),
.Y(n_6845)
);

INVx1_ASAP7_75t_L g6846 ( 
.A(n_6710),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_6608),
.Y(n_6847)
);

INVxp67_ASAP7_75t_L g6848 ( 
.A(n_6725),
.Y(n_6848)
);

OR2x2_ASAP7_75t_L g6849 ( 
.A(n_6644),
.B(n_6551),
.Y(n_6849)
);

INVx1_ASAP7_75t_L g6850 ( 
.A(n_6614),
.Y(n_6850)
);

AOI22xp5_ASAP7_75t_L g6851 ( 
.A1(n_6600),
.A2(n_6616),
.B1(n_6610),
.B2(n_6746),
.Y(n_6851)
);

AND2x2_ASAP7_75t_L g6852 ( 
.A(n_6650),
.B(n_6662),
.Y(n_6852)
);

INVx1_ASAP7_75t_L g6853 ( 
.A(n_6746),
.Y(n_6853)
);

AND2x2_ASAP7_75t_L g6854 ( 
.A(n_6680),
.B(n_6531),
.Y(n_6854)
);

INVx1_ASAP7_75t_L g6855 ( 
.A(n_6772),
.Y(n_6855)
);

INVx2_ASAP7_75t_L g6856 ( 
.A(n_6742),
.Y(n_6856)
);

AND2x4_ASAP7_75t_L g6857 ( 
.A(n_6639),
.B(n_6588),
.Y(n_6857)
);

NAND2xp5_ASAP7_75t_L g6858 ( 
.A(n_6634),
.B(n_6569),
.Y(n_6858)
);

AND2x4_ASAP7_75t_SL g6859 ( 
.A(n_6595),
.B(n_6588),
.Y(n_6859)
);

INVx1_ASAP7_75t_SL g6860 ( 
.A(n_6603),
.Y(n_6860)
);

INVx1_ASAP7_75t_L g6861 ( 
.A(n_6772),
.Y(n_6861)
);

INVx2_ASAP7_75t_L g6862 ( 
.A(n_6698),
.Y(n_6862)
);

NAND2xp5_ASAP7_75t_SL g6863 ( 
.A(n_6620),
.B(n_6420),
.Y(n_6863)
);

AND2x4_ASAP7_75t_L g6864 ( 
.A(n_6646),
.B(n_5219),
.Y(n_6864)
);

INVx2_ASAP7_75t_SL g6865 ( 
.A(n_6628),
.Y(n_6865)
);

INVx1_ASAP7_75t_L g6866 ( 
.A(n_6621),
.Y(n_6866)
);

AND2x2_ASAP7_75t_L g6867 ( 
.A(n_6622),
.B(n_6570),
.Y(n_6867)
);

INVx1_ASAP7_75t_L g6868 ( 
.A(n_6624),
.Y(n_6868)
);

OR2x2_ASAP7_75t_L g6869 ( 
.A(n_6654),
.B(n_6555),
.Y(n_6869)
);

AND2x2_ASAP7_75t_L g6870 ( 
.A(n_6601),
.B(n_6549),
.Y(n_6870)
);

NAND2xp5_ASAP7_75t_L g6871 ( 
.A(n_6676),
.B(n_6540),
.Y(n_6871)
);

NOR2xp33_ASAP7_75t_L g6872 ( 
.A(n_6692),
.B(n_6568),
.Y(n_6872)
);

INVx3_ASAP7_75t_L g6873 ( 
.A(n_6652),
.Y(n_6873)
);

AND2x2_ASAP7_75t_L g6874 ( 
.A(n_6684),
.B(n_6688),
.Y(n_6874)
);

INVx1_ASAP7_75t_L g6875 ( 
.A(n_6600),
.Y(n_6875)
);

INVx1_ASAP7_75t_L g6876 ( 
.A(n_6610),
.Y(n_6876)
);

NOR3xp33_ASAP7_75t_L g6877 ( 
.A(n_6729),
.B(n_6568),
.C(n_5106),
.Y(n_6877)
);

INVx1_ASAP7_75t_L g6878 ( 
.A(n_6616),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6642),
.Y(n_6879)
);

INVx1_ASAP7_75t_L g6880 ( 
.A(n_6642),
.Y(n_6880)
);

NOR2xp33_ASAP7_75t_L g6881 ( 
.A(n_6692),
.B(n_5226),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_6631),
.Y(n_6882)
);

AND2x2_ASAP7_75t_L g6883 ( 
.A(n_6649),
.B(n_5226),
.Y(n_6883)
);

AND2x2_ASAP7_75t_L g6884 ( 
.A(n_6743),
.B(n_5227),
.Y(n_6884)
);

AND2x2_ASAP7_75t_L g6885 ( 
.A(n_6659),
.B(n_5227),
.Y(n_6885)
);

INVx1_ASAP7_75t_L g6886 ( 
.A(n_6633),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_6640),
.Y(n_6887)
);

INVx2_ASAP7_75t_SL g6888 ( 
.A(n_6652),
.Y(n_6888)
);

INVx3_ASAP7_75t_L g6889 ( 
.A(n_6748),
.Y(n_6889)
);

INVx2_ASAP7_75t_SL g6890 ( 
.A(n_6671),
.Y(n_6890)
);

CKINVDCx8_ASAP7_75t_R g6891 ( 
.A(n_6814),
.Y(n_6891)
);

INVxp67_ASAP7_75t_L g6892 ( 
.A(n_6725),
.Y(n_6892)
);

AND2x2_ASAP7_75t_L g6893 ( 
.A(n_6695),
.B(n_5234),
.Y(n_6893)
);

AND2x2_ASAP7_75t_L g6894 ( 
.A(n_6637),
.B(n_5234),
.Y(n_6894)
);

NAND2xp5_ASAP7_75t_L g6895 ( 
.A(n_6667),
.B(n_6557),
.Y(n_6895)
);

AOI22xp5_ASAP7_75t_L g6896 ( 
.A1(n_6669),
.A2(n_6566),
.B1(n_6543),
.B2(n_6463),
.Y(n_6896)
);

NAND2xp5_ASAP7_75t_SL g6897 ( 
.A(n_6612),
.B(n_4333),
.Y(n_6897)
);

OR2x2_ASAP7_75t_L g6898 ( 
.A(n_6661),
.B(n_5240),
.Y(n_6898)
);

O2A1O1Ixp5_ASAP7_75t_L g6899 ( 
.A1(n_6781),
.A2(n_4582),
.B(n_4603),
.C(n_4564),
.Y(n_6899)
);

INVx1_ASAP7_75t_L g6900 ( 
.A(n_6669),
.Y(n_6900)
);

AND3x2_ASAP7_75t_L g6901 ( 
.A(n_6630),
.B(n_6587),
.C(n_4814),
.Y(n_6901)
);

INVx2_ASAP7_75t_SL g6902 ( 
.A(n_6678),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6778),
.Y(n_6903)
);

AND2x2_ASAP7_75t_L g6904 ( 
.A(n_6714),
.B(n_5331),
.Y(n_6904)
);

INVxp67_ASAP7_75t_L g6905 ( 
.A(n_6619),
.Y(n_6905)
);

INVx1_ASAP7_75t_SL g6906 ( 
.A(n_6673),
.Y(n_6906)
);

INVx1_ASAP7_75t_L g6907 ( 
.A(n_6722),
.Y(n_6907)
);

INVx1_ASAP7_75t_L g6908 ( 
.A(n_6736),
.Y(n_6908)
);

NAND2x1p5_ASAP7_75t_L g6909 ( 
.A(n_6597),
.B(n_4209),
.Y(n_6909)
);

INVxp67_ASAP7_75t_L g6910 ( 
.A(n_6686),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_6605),
.Y(n_6911)
);

INVx1_ASAP7_75t_L g6912 ( 
.A(n_6632),
.Y(n_6912)
);

INVx1_ASAP7_75t_L g6913 ( 
.A(n_6653),
.Y(n_6913)
);

NAND2xp5_ASAP7_75t_L g6914 ( 
.A(n_6667),
.B(n_5240),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_6774),
.Y(n_6915)
);

INVx1_ASAP7_75t_L g6916 ( 
.A(n_6819),
.Y(n_6916)
);

NOR2xp33_ASAP7_75t_L g6917 ( 
.A(n_6602),
.B(n_5254),
.Y(n_6917)
);

NAND2xp5_ASAP7_75t_L g6918 ( 
.A(n_6741),
.B(n_5254),
.Y(n_6918)
);

AND2x2_ASAP7_75t_L g6919 ( 
.A(n_6715),
.B(n_5332),
.Y(n_6919)
);

INVx1_ASAP7_75t_L g6920 ( 
.A(n_6790),
.Y(n_6920)
);

AOI33xp33_ASAP7_75t_L g6921 ( 
.A1(n_6785),
.A2(n_5273),
.A3(n_5265),
.B1(n_5276),
.B2(n_5268),
.B3(n_5260),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6793),
.Y(n_6922)
);

OR2x2_ASAP7_75t_L g6923 ( 
.A(n_6779),
.B(n_6663),
.Y(n_6923)
);

INVx1_ASAP7_75t_L g6924 ( 
.A(n_6789),
.Y(n_6924)
);

INVx2_ASAP7_75t_L g6925 ( 
.A(n_6728),
.Y(n_6925)
);

INVx2_ASAP7_75t_SL g6926 ( 
.A(n_6712),
.Y(n_6926)
);

AND2x4_ASAP7_75t_L g6927 ( 
.A(n_6660),
.B(n_5260),
.Y(n_6927)
);

INVx1_ASAP7_75t_L g6928 ( 
.A(n_6777),
.Y(n_6928)
);

INVx1_ASAP7_75t_L g6929 ( 
.A(n_6777),
.Y(n_6929)
);

OR2x2_ASAP7_75t_L g6930 ( 
.A(n_6656),
.B(n_5265),
.Y(n_6930)
);

INVx1_ASAP7_75t_L g6931 ( 
.A(n_6726),
.Y(n_6931)
);

INVx2_ASAP7_75t_L g6932 ( 
.A(n_6665),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_6685),
.Y(n_6933)
);

INVx1_ASAP7_75t_L g6934 ( 
.A(n_6685),
.Y(n_6934)
);

INVx2_ASAP7_75t_L g6935 ( 
.A(n_6672),
.Y(n_6935)
);

NOR2xp33_ASAP7_75t_L g6936 ( 
.A(n_6731),
.B(n_5268),
.Y(n_6936)
);

NAND2xp5_ASAP7_75t_L g6937 ( 
.A(n_6769),
.B(n_6775),
.Y(n_6937)
);

INVx1_ASAP7_75t_L g6938 ( 
.A(n_6817),
.Y(n_6938)
);

INVx1_ASAP7_75t_L g6939 ( 
.A(n_6784),
.Y(n_6939)
);

INVx1_ASAP7_75t_L g6940 ( 
.A(n_6648),
.Y(n_6940)
);

OR2x2_ASAP7_75t_L g6941 ( 
.A(n_6776),
.B(n_5273),
.Y(n_6941)
);

OR2x2_ASAP7_75t_L g6942 ( 
.A(n_6782),
.B(n_5276),
.Y(n_6942)
);

AND2x4_ASAP7_75t_L g6943 ( 
.A(n_6674),
.B(n_5279),
.Y(n_6943)
);

NOR2x1p5_ASAP7_75t_L g6944 ( 
.A(n_6677),
.B(n_4209),
.Y(n_6944)
);

AND2x2_ASAP7_75t_L g6945 ( 
.A(n_6753),
.B(n_5343),
.Y(n_6945)
);

INVx1_ASAP7_75t_L g6946 ( 
.A(n_6749),
.Y(n_6946)
);

OR2x2_ASAP7_75t_L g6947 ( 
.A(n_6596),
.B(n_5279),
.Y(n_6947)
);

AND2x2_ASAP7_75t_L g6948 ( 
.A(n_6768),
.B(n_5343),
.Y(n_6948)
);

INVx1_ASAP7_75t_L g6949 ( 
.A(n_6750),
.Y(n_6949)
);

OR2x2_ASAP7_75t_L g6950 ( 
.A(n_6596),
.B(n_5296),
.Y(n_6950)
);

INVx1_ASAP7_75t_L g6951 ( 
.A(n_6655),
.Y(n_6951)
);

AND2x2_ASAP7_75t_L g6952 ( 
.A(n_6798),
.B(n_6682),
.Y(n_6952)
);

AND2x4_ASAP7_75t_SL g6953 ( 
.A(n_6761),
.B(n_4333),
.Y(n_6953)
);

INVx1_ASAP7_75t_L g6954 ( 
.A(n_6657),
.Y(n_6954)
);

AND2x2_ASAP7_75t_L g6955 ( 
.A(n_6798),
.B(n_5313),
.Y(n_6955)
);

NOR2xp33_ASAP7_75t_L g6956 ( 
.A(n_6732),
.B(n_5296),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_6770),
.Y(n_6957)
);

INVx2_ASAP7_75t_L g6958 ( 
.A(n_6681),
.Y(n_6958)
);

INVx1_ASAP7_75t_L g6959 ( 
.A(n_6734),
.Y(n_6959)
);

OR2x2_ASAP7_75t_L g6960 ( 
.A(n_6787),
.B(n_5297),
.Y(n_6960)
);

OR2x2_ASAP7_75t_L g6961 ( 
.A(n_6724),
.B(n_5297),
.Y(n_6961)
);

INVx1_ASAP7_75t_L g6962 ( 
.A(n_6641),
.Y(n_6962)
);

NAND2xp5_ASAP7_75t_L g6963 ( 
.A(n_6691),
.B(n_5298),
.Y(n_6963)
);

INVx1_ASAP7_75t_L g6964 ( 
.A(n_6709),
.Y(n_6964)
);

NAND2xp5_ASAP7_75t_L g6965 ( 
.A(n_6691),
.B(n_5298),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6727),
.Y(n_6966)
);

NAND2xp5_ASAP7_75t_L g6967 ( 
.A(n_6747),
.B(n_5305),
.Y(n_6967)
);

NAND2xp5_ASAP7_75t_L g6968 ( 
.A(n_6816),
.B(n_5305),
.Y(n_6968)
);

NAND2xp5_ASAP7_75t_L g6969 ( 
.A(n_6818),
.B(n_5310),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6733),
.Y(n_6970)
);

INVx1_ASAP7_75t_L g6971 ( 
.A(n_6664),
.Y(n_6971)
);

OR2x2_ASAP7_75t_L g6972 ( 
.A(n_6651),
.B(n_5310),
.Y(n_6972)
);

NOR5xp2_ASAP7_75t_L g6973 ( 
.A(n_6598),
.B(n_5317),
.C(n_5331),
.D(n_5313),
.E(n_5311),
.Y(n_6973)
);

AND2x2_ASAP7_75t_L g6974 ( 
.A(n_6796),
.B(n_5332),
.Y(n_6974)
);

INVx1_ASAP7_75t_L g6975 ( 
.A(n_6636),
.Y(n_6975)
);

NAND2xp5_ASAP7_75t_L g6976 ( 
.A(n_6626),
.B(n_5311),
.Y(n_6976)
);

INVx2_ASAP7_75t_L g6977 ( 
.A(n_6786),
.Y(n_6977)
);

AND2x2_ASAP7_75t_L g6978 ( 
.A(n_6756),
.B(n_5317),
.Y(n_6978)
);

INVx1_ASAP7_75t_L g6979 ( 
.A(n_6658),
.Y(n_6979)
);

INVx2_ASAP7_75t_L g6980 ( 
.A(n_6748),
.Y(n_6980)
);

OR2x2_ASAP7_75t_L g6981 ( 
.A(n_6668),
.B(n_5312),
.Y(n_6981)
);

AND2x2_ASAP7_75t_L g6982 ( 
.A(n_6792),
.B(n_4209),
.Y(n_6982)
);

INVx2_ASAP7_75t_L g6983 ( 
.A(n_6752),
.Y(n_6983)
);

NAND2xp5_ASAP7_75t_L g6984 ( 
.A(n_6805),
.B(n_4972),
.Y(n_6984)
);

NOR2x1p5_ASAP7_75t_L g6985 ( 
.A(n_6745),
.B(n_4218),
.Y(n_6985)
);

AND2x4_ASAP7_75t_L g6986 ( 
.A(n_6751),
.B(n_6806),
.Y(n_6986)
);

AND2x2_ASAP7_75t_L g6987 ( 
.A(n_6629),
.B(n_4218),
.Y(n_6987)
);

NAND2xp5_ASAP7_75t_L g6988 ( 
.A(n_6718),
.B(n_4983),
.Y(n_6988)
);

NAND2xp5_ASAP7_75t_L g6989 ( 
.A(n_6718),
.B(n_4983),
.Y(n_6989)
);

AND2x2_ASAP7_75t_L g6990 ( 
.A(n_6773),
.B(n_4222),
.Y(n_6990)
);

OAI21xp33_ASAP7_75t_L g6991 ( 
.A1(n_6702),
.A2(n_4222),
.B(n_4860),
.Y(n_6991)
);

AND2x2_ASAP7_75t_L g6992 ( 
.A(n_6763),
.B(n_4222),
.Y(n_6992)
);

OR2x2_ASAP7_75t_L g6993 ( 
.A(n_6689),
.B(n_5312),
.Y(n_6993)
);

AND2x2_ASAP7_75t_L g6994 ( 
.A(n_6780),
.B(n_3980),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6767),
.Y(n_6995)
);

NAND2x1p5_ASAP7_75t_L g6996 ( 
.A(n_6723),
.B(n_4379),
.Y(n_6996)
);

AND2x2_ASAP7_75t_L g6997 ( 
.A(n_6783),
.B(n_3980),
.Y(n_6997)
);

NAND2x1p5_ASAP7_75t_L g6998 ( 
.A(n_6700),
.B(n_4379),
.Y(n_6998)
);

OAI21xp5_ASAP7_75t_SL g6999 ( 
.A1(n_6670),
.A2(n_4406),
.B(n_4379),
.Y(n_6999)
);

BUFx2_ASAP7_75t_L g7000 ( 
.A(n_6752),
.Y(n_7000)
);

INVx1_ASAP7_75t_L g7001 ( 
.A(n_6800),
.Y(n_7001)
);

AND2x2_ASAP7_75t_L g7002 ( 
.A(n_6643),
.B(n_3932),
.Y(n_7002)
);

AND2x2_ASAP7_75t_L g7003 ( 
.A(n_6694),
.B(n_6803),
.Y(n_7003)
);

OR2x2_ASAP7_75t_L g7004 ( 
.A(n_6696),
.B(n_5330),
.Y(n_7004)
);

HB1xp67_ASAP7_75t_L g7005 ( 
.A(n_6804),
.Y(n_7005)
);

NOR2xp33_ASAP7_75t_L g7006 ( 
.A(n_6638),
.B(n_4379),
.Y(n_7006)
);

BUFx2_ASAP7_75t_L g7007 ( 
.A(n_6759),
.Y(n_7007)
);

NAND2xp5_ASAP7_75t_L g7008 ( 
.A(n_6807),
.B(n_5197),
.Y(n_7008)
);

INVx1_ASAP7_75t_SL g7009 ( 
.A(n_6820),
.Y(n_7009)
);

AOI22xp5_ASAP7_75t_L g7010 ( 
.A1(n_6812),
.A2(n_5252),
.B1(n_5034),
.B2(n_5232),
.Y(n_7010)
);

INVx2_ASAP7_75t_L g7011 ( 
.A(n_6766),
.Y(n_7011)
);

AND2x2_ASAP7_75t_L g7012 ( 
.A(n_6762),
.B(n_3932),
.Y(n_7012)
);

INVx1_ASAP7_75t_L g7013 ( 
.A(n_6815),
.Y(n_7013)
);

NAND2x1_ASAP7_75t_L g7014 ( 
.A(n_6822),
.B(n_4564),
.Y(n_7014)
);

INVx2_ASAP7_75t_L g7015 ( 
.A(n_6802),
.Y(n_7015)
);

AND2x2_ASAP7_75t_L g7016 ( 
.A(n_6764),
.B(n_3996),
.Y(n_7016)
);

NAND2xp5_ASAP7_75t_L g7017 ( 
.A(n_6675),
.B(n_5197),
.Y(n_7017)
);

INVx1_ASAP7_75t_L g7018 ( 
.A(n_6821),
.Y(n_7018)
);

AOI21xp5_ASAP7_75t_L g7019 ( 
.A1(n_6853),
.A2(n_6675),
.B(n_6611),
.Y(n_7019)
);

AND2x2_ASAP7_75t_L g7020 ( 
.A(n_6852),
.B(n_6666),
.Y(n_7020)
);

AND2x2_ASAP7_75t_L g7021 ( 
.A(n_6874),
.B(n_6701),
.Y(n_7021)
);

OAI22xp5_ASAP7_75t_L g7022 ( 
.A1(n_6831),
.A2(n_6754),
.B1(n_6708),
.B2(n_6670),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_6873),
.Y(n_7023)
);

AND2x2_ASAP7_75t_L g7024 ( 
.A(n_6860),
.B(n_6706),
.Y(n_7024)
);

AND2x2_ASAP7_75t_L g7025 ( 
.A(n_6888),
.B(n_6707),
.Y(n_7025)
);

INVxp33_ASAP7_75t_L g7026 ( 
.A(n_6823),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_6873),
.Y(n_7027)
);

INVx1_ASAP7_75t_SL g7028 ( 
.A(n_6823),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_7000),
.Y(n_7029)
);

AOI32xp33_ASAP7_75t_L g7030 ( 
.A1(n_6855),
.A2(n_6599),
.A3(n_6765),
.B1(n_6638),
.B2(n_6738),
.Y(n_7030)
);

NAND2xp5_ASAP7_75t_L g7031 ( 
.A(n_6865),
.B(n_6801),
.Y(n_7031)
);

NAND2xp5_ASAP7_75t_L g7032 ( 
.A(n_6926),
.B(n_6808),
.Y(n_7032)
);

AOI22xp5_ASAP7_75t_L g7033 ( 
.A1(n_6861),
.A2(n_6880),
.B1(n_6879),
.B2(n_6851),
.Y(n_7033)
);

OR2x2_ASAP7_75t_L g7034 ( 
.A(n_6839),
.B(n_6757),
.Y(n_7034)
);

OAI222xp33_ASAP7_75t_L g7035 ( 
.A1(n_6896),
.A2(n_6699),
.B1(n_6703),
.B2(n_6791),
.C1(n_6704),
.C2(n_6758),
.Y(n_7035)
);

AND2x2_ASAP7_75t_L g7036 ( 
.A(n_6952),
.B(n_6717),
.Y(n_7036)
);

AND2x4_ASAP7_75t_SL g7037 ( 
.A(n_6977),
.B(n_6720),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6841),
.Y(n_7038)
);

INVx1_ASAP7_75t_L g7039 ( 
.A(n_6948),
.Y(n_7039)
);

NAND2xp5_ASAP7_75t_L g7040 ( 
.A(n_6857),
.B(n_6809),
.Y(n_7040)
);

AND2x4_ASAP7_75t_L g7041 ( 
.A(n_6827),
.B(n_6810),
.Y(n_7041)
);

INVx1_ASAP7_75t_L g7042 ( 
.A(n_6923),
.Y(n_7042)
);

AOI221xp5_ASAP7_75t_L g7043 ( 
.A1(n_6900),
.A2(n_6611),
.B1(n_6623),
.B2(n_6713),
.C(n_6799),
.Y(n_7043)
);

INVx2_ASAP7_75t_L g7044 ( 
.A(n_6889),
.Y(n_7044)
);

OAI21xp33_ASAP7_75t_L g7045 ( 
.A1(n_6834),
.A2(n_6716),
.B(n_6788),
.Y(n_7045)
);

INVx1_ASAP7_75t_L g7046 ( 
.A(n_6933),
.Y(n_7046)
);

O2A1O1Ixp5_ASAP7_75t_R g7047 ( 
.A1(n_6836),
.A2(n_6744),
.B(n_6719),
.C(n_6738),
.Y(n_7047)
);

INVx1_ASAP7_75t_L g7048 ( 
.A(n_6933),
.Y(n_7048)
);

AND2x4_ASAP7_75t_L g7049 ( 
.A(n_6832),
.B(n_6760),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_6934),
.Y(n_7050)
);

INVx1_ASAP7_75t_L g7051 ( 
.A(n_6934),
.Y(n_7051)
);

INVx1_ASAP7_75t_L g7052 ( 
.A(n_6871),
.Y(n_7052)
);

NOR2x1_ASAP7_75t_L g7053 ( 
.A(n_6889),
.B(n_6683),
.Y(n_7053)
);

NAND4xp25_ASAP7_75t_L g7054 ( 
.A(n_7006),
.B(n_6719),
.C(n_6737),
.D(n_6740),
.Y(n_7054)
);

NAND2xp5_ASAP7_75t_L g7055 ( 
.A(n_6857),
.B(n_6683),
.Y(n_7055)
);

AND2x4_ASAP7_75t_SL g7056 ( 
.A(n_6925),
.B(n_4379),
.Y(n_7056)
);

AND2x2_ASAP7_75t_L g7057 ( 
.A(n_6835),
.B(n_6740),
.Y(n_7057)
);

OAI21xp5_ASAP7_75t_L g7058 ( 
.A1(n_6895),
.A2(n_6797),
.B(n_6697),
.Y(n_7058)
);

INVx1_ASAP7_75t_L g7059 ( 
.A(n_6843),
.Y(n_7059)
);

NAND2xp5_ASAP7_75t_L g7060 ( 
.A(n_6872),
.B(n_6735),
.Y(n_7060)
);

INVx1_ASAP7_75t_L g7061 ( 
.A(n_6856),
.Y(n_7061)
);

INVx1_ASAP7_75t_L g7062 ( 
.A(n_6891),
.Y(n_7062)
);

BUFx3_ASAP7_75t_L g7063 ( 
.A(n_6986),
.Y(n_7063)
);

AOI22xp5_ASAP7_75t_L g7064 ( 
.A1(n_6939),
.A2(n_6735),
.B1(n_6687),
.B2(n_6730),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_6826),
.Y(n_7065)
);

NAND2x1_ASAP7_75t_L g7066 ( 
.A(n_6973),
.B(n_6822),
.Y(n_7066)
);

AOI22xp33_ASAP7_75t_L g7067 ( 
.A1(n_6825),
.A2(n_6811),
.B1(n_4941),
.B2(n_6721),
.Y(n_7067)
);

OAI21xp5_ASAP7_75t_SL g7068 ( 
.A1(n_6901),
.A2(n_6999),
.B(n_6833),
.Y(n_7068)
);

INVx2_ASAP7_75t_L g7069 ( 
.A(n_6845),
.Y(n_7069)
);

NAND2xp5_ASAP7_75t_L g7070 ( 
.A(n_6902),
.B(n_6760),
.Y(n_7070)
);

AND2x2_ASAP7_75t_L g7071 ( 
.A(n_6838),
.B(n_6737),
.Y(n_7071)
);

OAI22xp5_ASAP7_75t_L g7072 ( 
.A1(n_6830),
.A2(n_6771),
.B1(n_5232),
.B2(n_4582),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_6928),
.Y(n_7073)
);

OAI221xp5_ASAP7_75t_L g7074 ( 
.A1(n_6877),
.A2(n_6811),
.B1(n_6771),
.B2(n_6711),
.C(n_6813),
.Y(n_7074)
);

INVx2_ASAP7_75t_L g7075 ( 
.A(n_6845),
.Y(n_7075)
);

OAI22xp33_ASAP7_75t_L g7076 ( 
.A1(n_6939),
.A2(n_6813),
.B1(n_5290),
.B2(n_5267),
.Y(n_7076)
);

XNOR2xp5_ASAP7_75t_L g7077 ( 
.A(n_6944),
.B(n_5267),
.Y(n_7077)
);

AND2x2_ASAP7_75t_L g7078 ( 
.A(n_6862),
.B(n_6932),
.Y(n_7078)
);

AOI22xp5_ASAP7_75t_L g7079 ( 
.A1(n_7007),
.A2(n_5290),
.B1(n_5105),
.B2(n_5109),
.Y(n_7079)
);

NAND3xp33_ASAP7_75t_L g7080 ( 
.A(n_6924),
.B(n_5208),
.C(n_5170),
.Y(n_7080)
);

AND2x4_ASAP7_75t_L g7081 ( 
.A(n_6935),
.B(n_5220),
.Y(n_7081)
);

NAND2xp5_ASAP7_75t_L g7082 ( 
.A(n_6945),
.B(n_5197),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6928),
.Y(n_7083)
);

AOI22xp5_ASAP7_75t_L g7084 ( 
.A1(n_6842),
.A2(n_6846),
.B1(n_7017),
.B2(n_6936),
.Y(n_7084)
);

OAI21xp33_ASAP7_75t_L g7085 ( 
.A1(n_6975),
.A2(n_4863),
.B(n_4860),
.Y(n_7085)
);

AND2x2_ASAP7_75t_L g7086 ( 
.A(n_6870),
.B(n_3996),
.Y(n_7086)
);

NAND2xp5_ASAP7_75t_L g7087 ( 
.A(n_6913),
.B(n_5330),
.Y(n_7087)
);

OAI221xp5_ASAP7_75t_L g7088 ( 
.A1(n_6924),
.A2(n_5151),
.B1(n_5145),
.B2(n_5110),
.C(n_5111),
.Y(n_7088)
);

OAI32xp33_ASAP7_75t_L g7089 ( 
.A1(n_6976),
.A2(n_4603),
.A3(n_4631),
.B1(n_4624),
.B2(n_4564),
.Y(n_7089)
);

INVx2_ASAP7_75t_L g7090 ( 
.A(n_6909),
.Y(n_7090)
);

AOI21xp33_ASAP7_75t_SL g7091 ( 
.A1(n_6890),
.A2(n_5177),
.B(n_5090),
.Y(n_7091)
);

OR2x2_ASAP7_75t_L g7092 ( 
.A(n_6849),
.B(n_5027),
.Y(n_7092)
);

O2A1O1Ixp33_ASAP7_75t_SL g7093 ( 
.A1(n_7014),
.A2(n_4603),
.B(n_4624),
.C(n_4564),
.Y(n_7093)
);

INVxp33_ASAP7_75t_L g7094 ( 
.A(n_6854),
.Y(n_7094)
);

A2O1A1Ixp33_ASAP7_75t_L g7095 ( 
.A1(n_6956),
.A2(n_5300),
.B(n_4547),
.C(n_5109),
.Y(n_7095)
);

INVx1_ASAP7_75t_L g7096 ( 
.A(n_6929),
.Y(n_7096)
);

INVx1_ASAP7_75t_L g7097 ( 
.A(n_6929),
.Y(n_7097)
);

NAND2xp5_ASAP7_75t_L g7098 ( 
.A(n_7011),
.B(n_5027),
.Y(n_7098)
);

INVx1_ASAP7_75t_L g7099 ( 
.A(n_6930),
.Y(n_7099)
);

HB1xp67_ASAP7_75t_L g7100 ( 
.A(n_6958),
.Y(n_7100)
);

OAI222xp33_ASAP7_75t_L g7101 ( 
.A1(n_7013),
.A2(n_4574),
.B1(n_5111),
.B2(n_5128),
.C1(n_5110),
.C2(n_5108),
.Y(n_7101)
);

INVx1_ASAP7_75t_L g7102 ( 
.A(n_6824),
.Y(n_7102)
);

OR2x2_ASAP7_75t_L g7103 ( 
.A(n_6937),
.B(n_4543),
.Y(n_7103)
);

NAND2x1_ASAP7_75t_SL g7104 ( 
.A(n_6840),
.B(n_4582),
.Y(n_7104)
);

INVxp67_ASAP7_75t_SL g7105 ( 
.A(n_6910),
.Y(n_7105)
);

NAND2xp5_ASAP7_75t_L g7106 ( 
.A(n_6964),
.B(n_4549),
.Y(n_7106)
);

AOI22xp33_ASAP7_75t_L g7107 ( 
.A1(n_6875),
.A2(n_4941),
.B1(n_5128),
.B2(n_5108),
.Y(n_7107)
);

OR2x2_ASAP7_75t_L g7108 ( 
.A(n_6915),
.B(n_4549),
.Y(n_7108)
);

AND2x2_ASAP7_75t_L g7109 ( 
.A(n_6982),
.B(n_6844),
.Y(n_7109)
);

INVx1_ASAP7_75t_L g7110 ( 
.A(n_6981),
.Y(n_7110)
);

INVx2_ASAP7_75t_L g7111 ( 
.A(n_6996),
.Y(n_7111)
);

INVx1_ASAP7_75t_L g7112 ( 
.A(n_6993),
.Y(n_7112)
);

AND2x4_ASAP7_75t_L g7113 ( 
.A(n_6980),
.B(n_5300),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_7004),
.Y(n_7114)
);

AOI22xp5_ASAP7_75t_L g7115 ( 
.A1(n_6917),
.A2(n_5136),
.B1(n_5147),
.B2(n_5130),
.Y(n_7115)
);

AND2x4_ASAP7_75t_L g7116 ( 
.A(n_6983),
.B(n_4582),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_6824),
.Y(n_7117)
);

NAND2xp5_ASAP7_75t_L g7118 ( 
.A(n_6931),
.B(n_4552),
.Y(n_7118)
);

AND2x2_ASAP7_75t_L g7119 ( 
.A(n_6829),
.B(n_4856),
.Y(n_7119)
);

OR2x2_ASAP7_75t_L g7120 ( 
.A(n_6984),
.B(n_4552),
.Y(n_7120)
);

NAND3xp33_ASAP7_75t_L g7121 ( 
.A(n_7018),
.B(n_5151),
.C(n_5145),
.Y(n_7121)
);

NAND3xp33_ASAP7_75t_SL g7122 ( 
.A(n_6906),
.B(n_5136),
.C(n_5130),
.Y(n_7122)
);

NAND3xp33_ASAP7_75t_SL g7123 ( 
.A(n_7009),
.B(n_5148),
.C(n_5147),
.Y(n_7123)
);

NOR2xp67_ASAP7_75t_L g7124 ( 
.A(n_6848),
.B(n_4675),
.Y(n_7124)
);

AND2x2_ASAP7_75t_L g7125 ( 
.A(n_6987),
.B(n_4859),
.Y(n_7125)
);

INVx1_ASAP7_75t_SL g7126 ( 
.A(n_6859),
.Y(n_7126)
);

OR2x2_ASAP7_75t_L g7127 ( 
.A(n_6911),
.B(n_4555),
.Y(n_7127)
);

INVxp67_ASAP7_75t_L g7128 ( 
.A(n_6920),
.Y(n_7128)
);

NAND2xp5_ASAP7_75t_L g7129 ( 
.A(n_6946),
.B(n_4555),
.Y(n_7129)
);

OR2x2_ASAP7_75t_L g7130 ( 
.A(n_6912),
.B(n_4561),
.Y(n_7130)
);

NOR2xp33_ASAP7_75t_L g7131 ( 
.A(n_6892),
.B(n_4379),
.Y(n_7131)
);

INVx1_ASAP7_75t_L g7132 ( 
.A(n_6907),
.Y(n_7132)
);

INVx1_ASAP7_75t_L g7133 ( 
.A(n_6908),
.Y(n_7133)
);

OR2x2_ASAP7_75t_L g7134 ( 
.A(n_6903),
.B(n_4561),
.Y(n_7134)
);

NAND3xp33_ASAP7_75t_SL g7135 ( 
.A(n_6858),
.B(n_5149),
.C(n_5148),
.Y(n_7135)
);

OR2x2_ASAP7_75t_L g7136 ( 
.A(n_6916),
.B(n_4563),
.Y(n_7136)
);

INVx1_ASAP7_75t_L g7137 ( 
.A(n_7002),
.Y(n_7137)
);

INVx1_ASAP7_75t_SL g7138 ( 
.A(n_6869),
.Y(n_7138)
);

INVx1_ASAP7_75t_L g7139 ( 
.A(n_7012),
.Y(n_7139)
);

OR2x2_ASAP7_75t_L g7140 ( 
.A(n_6962),
.B(n_4563),
.Y(n_7140)
);

INVxp67_ASAP7_75t_L g7141 ( 
.A(n_6920),
.Y(n_7141)
);

INVx1_ASAP7_75t_L g7142 ( 
.A(n_7016),
.Y(n_7142)
);

INVx1_ASAP7_75t_L g7143 ( 
.A(n_7005),
.Y(n_7143)
);

NAND2xp5_ASAP7_75t_L g7144 ( 
.A(n_6957),
.B(n_4565),
.Y(n_7144)
);

INVxp67_ASAP7_75t_L g7145 ( 
.A(n_6922),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_6960),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_6883),
.Y(n_7147)
);

NAND2xp5_ASAP7_75t_L g7148 ( 
.A(n_6884),
.B(n_4565),
.Y(n_7148)
);

AOI221xp5_ASAP7_75t_L g7149 ( 
.A1(n_7018),
.A2(n_5165),
.B1(n_5169),
.B2(n_5164),
.C(n_5149),
.Y(n_7149)
);

OAI22xp5_ASAP7_75t_L g7150 ( 
.A1(n_6951),
.A2(n_4624),
.B1(n_4631),
.B2(n_4603),
.Y(n_7150)
);

INVxp67_ASAP7_75t_L g7151 ( 
.A(n_6922),
.Y(n_7151)
);

AND2x2_ASAP7_75t_L g7152 ( 
.A(n_7003),
.B(n_6992),
.Y(n_7152)
);

O2A1O1Ixp33_ASAP7_75t_SL g7153 ( 
.A1(n_6897),
.A2(n_4631),
.B(n_4636),
.C(n_4624),
.Y(n_7153)
);

INVx1_ASAP7_75t_L g7154 ( 
.A(n_6894),
.Y(n_7154)
);

OR2x2_ASAP7_75t_L g7155 ( 
.A(n_6988),
.B(n_4570),
.Y(n_7155)
);

OR2x2_ASAP7_75t_L g7156 ( 
.A(n_6989),
.B(n_4570),
.Y(n_7156)
);

NAND2x1p5_ASAP7_75t_L g7157 ( 
.A(n_6986),
.B(n_4406),
.Y(n_7157)
);

AOI32xp33_ASAP7_75t_L g7158 ( 
.A1(n_6938),
.A2(n_4870),
.A3(n_4706),
.B1(n_4675),
.B2(n_4659),
.Y(n_7158)
);

AOI33xp33_ASAP7_75t_L g7159 ( 
.A1(n_6882),
.A2(n_4913),
.A3(n_4865),
.B1(n_4923),
.B2(n_4883),
.B3(n_4863),
.Y(n_7159)
);

OR2x2_ASAP7_75t_L g7160 ( 
.A(n_6949),
.B(n_4575),
.Y(n_7160)
);

AND2x2_ASAP7_75t_L g7161 ( 
.A(n_6867),
.B(n_4859),
.Y(n_7161)
);

AOI33xp33_ASAP7_75t_L g7162 ( 
.A1(n_6886),
.A2(n_4923),
.A3(n_4865),
.B1(n_4925),
.B2(n_4913),
.B3(n_4883),
.Y(n_7162)
);

INVx1_ASAP7_75t_SL g7163 ( 
.A(n_6953),
.Y(n_7163)
);

OAI22xp5_ASAP7_75t_L g7164 ( 
.A1(n_6954),
.A2(n_4636),
.B1(n_4659),
.B2(n_4631),
.Y(n_7164)
);

INVx1_ASAP7_75t_L g7165 ( 
.A(n_6885),
.Y(n_7165)
);

NAND3xp33_ASAP7_75t_L g7166 ( 
.A(n_6863),
.B(n_6970),
.C(n_6966),
.Y(n_7166)
);

INVx2_ASAP7_75t_L g7167 ( 
.A(n_6998),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_6893),
.Y(n_7168)
);

INVxp67_ASAP7_75t_SL g7169 ( 
.A(n_6985),
.Y(n_7169)
);

NAND2xp5_ASAP7_75t_L g7170 ( 
.A(n_6904),
.B(n_4575),
.Y(n_7170)
);

INVx1_ASAP7_75t_L g7171 ( 
.A(n_6968),
.Y(n_7171)
);

NAND2xp5_ASAP7_75t_L g7172 ( 
.A(n_6919),
.B(n_6979),
.Y(n_7172)
);

INVx1_ASAP7_75t_L g7173 ( 
.A(n_6969),
.Y(n_7173)
);

OAI21xp33_ASAP7_75t_L g7174 ( 
.A1(n_6991),
.A2(n_7010),
.B(n_6990),
.Y(n_7174)
);

OR2x6_ASAP7_75t_L g7175 ( 
.A(n_6971),
.B(n_4574),
.Y(n_7175)
);

AOI21xp33_ASAP7_75t_L g7176 ( 
.A1(n_7013),
.A2(n_6914),
.B(n_6938),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_6961),
.Y(n_7177)
);

AOI22xp5_ASAP7_75t_L g7178 ( 
.A1(n_6876),
.A2(n_5165),
.B1(n_5169),
.B2(n_5164),
.Y(n_7178)
);

AND2x2_ASAP7_75t_L g7179 ( 
.A(n_6994),
.B(n_4861),
.Y(n_7179)
);

OAI31xp33_ASAP7_75t_L g7180 ( 
.A1(n_6878),
.A2(n_5193),
.A3(n_5194),
.B(n_5174),
.Y(n_7180)
);

O2A1O1Ixp5_ASAP7_75t_L g7181 ( 
.A1(n_6899),
.A2(n_4659),
.B(n_4675),
.C(n_4636),
.Y(n_7181)
);

INVx2_ASAP7_75t_SL g7182 ( 
.A(n_6978),
.Y(n_7182)
);

AOI32xp33_ASAP7_75t_L g7183 ( 
.A1(n_6828),
.A2(n_4910),
.A3(n_4675),
.B1(n_4696),
.B2(n_4659),
.Y(n_7183)
);

INVx1_ASAP7_75t_L g7184 ( 
.A(n_6941),
.Y(n_7184)
);

INVx1_ASAP7_75t_L g7185 ( 
.A(n_6942),
.Y(n_7185)
);

INVx1_ASAP7_75t_L g7186 ( 
.A(n_6898),
.Y(n_7186)
);

INVx1_ASAP7_75t_L g7187 ( 
.A(n_6955),
.Y(n_7187)
);

NOR2x1p5_ASAP7_75t_L g7188 ( 
.A(n_7015),
.B(n_4406),
.Y(n_7188)
);

NAND3xp33_ASAP7_75t_L g7189 ( 
.A(n_6940),
.B(n_5151),
.C(n_5145),
.Y(n_7189)
);

INVx2_ASAP7_75t_SL g7190 ( 
.A(n_6943),
.Y(n_7190)
);

NAND2xp5_ASAP7_75t_L g7191 ( 
.A(n_6943),
.B(n_4581),
.Y(n_7191)
);

OAI22xp33_ASAP7_75t_L g7192 ( 
.A1(n_6947),
.A2(n_5174),
.B1(n_5194),
.B2(n_5193),
.Y(n_7192)
);

NOR2xp33_ASAP7_75t_L g7193 ( 
.A(n_6905),
.B(n_4406),
.Y(n_7193)
);

AND2x2_ASAP7_75t_L g7194 ( 
.A(n_6997),
.B(n_4861),
.Y(n_7194)
);

NAND2xp5_ASAP7_75t_L g7195 ( 
.A(n_6927),
.B(n_4581),
.Y(n_7195)
);

AND2x2_ASAP7_75t_L g7196 ( 
.A(n_6887),
.B(n_4406),
.Y(n_7196)
);

OAI21xp5_ASAP7_75t_L g7197 ( 
.A1(n_6950),
.A2(n_4502),
.B(n_5195),
.Y(n_7197)
);

NAND2xp5_ASAP7_75t_L g7198 ( 
.A(n_7063),
.B(n_6927),
.Y(n_7198)
);

OR2x2_ASAP7_75t_L g7199 ( 
.A(n_7028),
.B(n_7001),
.Y(n_7199)
);

INVx1_ASAP7_75t_L g7200 ( 
.A(n_7100),
.Y(n_7200)
);

INVx1_ASAP7_75t_SL g7201 ( 
.A(n_7126),
.Y(n_7201)
);

OAI21xp5_ASAP7_75t_L g7202 ( 
.A1(n_7019),
.A2(n_6881),
.B(n_6995),
.Y(n_7202)
);

INVx1_ASAP7_75t_SL g7203 ( 
.A(n_7021),
.Y(n_7203)
);

INVx2_ASAP7_75t_L g7204 ( 
.A(n_7157),
.Y(n_7204)
);

AND2x2_ASAP7_75t_L g7205 ( 
.A(n_7020),
.B(n_6974),
.Y(n_7205)
);

NAND2xp5_ASAP7_75t_L g7206 ( 
.A(n_7049),
.B(n_6864),
.Y(n_7206)
);

INVx2_ASAP7_75t_L g7207 ( 
.A(n_7104),
.Y(n_7207)
);

AND2x2_ASAP7_75t_L g7208 ( 
.A(n_7109),
.B(n_6940),
.Y(n_7208)
);

NAND3x1_ASAP7_75t_SL g7209 ( 
.A(n_7053),
.B(n_6959),
.C(n_6921),
.Y(n_7209)
);

INVx1_ASAP7_75t_L g7210 ( 
.A(n_7040),
.Y(n_7210)
);

INVx1_ASAP7_75t_L g7211 ( 
.A(n_7036),
.Y(n_7211)
);

NAND2xp5_ASAP7_75t_L g7212 ( 
.A(n_7049),
.B(n_6864),
.Y(n_7212)
);

BUFx2_ASAP7_75t_L g7213 ( 
.A(n_7152),
.Y(n_7213)
);

AND2x2_ASAP7_75t_L g7214 ( 
.A(n_7078),
.B(n_6918),
.Y(n_7214)
);

AND2x2_ASAP7_75t_L g7215 ( 
.A(n_7026),
.B(n_6972),
.Y(n_7215)
);

INVx1_ASAP7_75t_L g7216 ( 
.A(n_7024),
.Y(n_7216)
);

CKINVDCx16_ASAP7_75t_R g7217 ( 
.A(n_7138),
.Y(n_7217)
);

NOR2x1_ASAP7_75t_L g7218 ( 
.A(n_7166),
.B(n_6828),
.Y(n_7218)
);

CKINVDCx16_ASAP7_75t_R g7219 ( 
.A(n_7034),
.Y(n_7219)
);

INVx2_ASAP7_75t_SL g7220 ( 
.A(n_7037),
.Y(n_7220)
);

NOR2x1_ASAP7_75t_SL g7221 ( 
.A(n_7190),
.B(n_6967),
.Y(n_7221)
);

AND2x2_ASAP7_75t_L g7222 ( 
.A(n_7119),
.B(n_6963),
.Y(n_7222)
);

INVx1_ASAP7_75t_L g7223 ( 
.A(n_7044),
.Y(n_7223)
);

AND2x2_ASAP7_75t_L g7224 ( 
.A(n_7086),
.B(n_6965),
.Y(n_7224)
);

INVx1_ASAP7_75t_SL g7225 ( 
.A(n_7055),
.Y(n_7225)
);

INVxp67_ASAP7_75t_L g7226 ( 
.A(n_7025),
.Y(n_7226)
);

INVx2_ASAP7_75t_L g7227 ( 
.A(n_7161),
.Y(n_7227)
);

NAND2xp5_ASAP7_75t_L g7228 ( 
.A(n_7057),
.B(n_7008),
.Y(n_7228)
);

INVx1_ASAP7_75t_L g7229 ( 
.A(n_7052),
.Y(n_7229)
);

CKINVDCx16_ASAP7_75t_R g7230 ( 
.A(n_7062),
.Y(n_7230)
);

AND2x4_ASAP7_75t_L g7231 ( 
.A(n_7041),
.B(n_6850),
.Y(n_7231)
);

OAI22xp5_ASAP7_75t_L g7232 ( 
.A1(n_7094),
.A2(n_6868),
.B1(n_6866),
.B2(n_6847),
.Y(n_7232)
);

NAND2xp5_ASAP7_75t_L g7233 ( 
.A(n_7182),
.B(n_7041),
.Y(n_7233)
);

HB1xp67_ASAP7_75t_L g7234 ( 
.A(n_7029),
.Y(n_7234)
);

NAND2xp5_ASAP7_75t_L g7235 ( 
.A(n_7039),
.B(n_6837),
.Y(n_7235)
);

NAND2xp5_ASAP7_75t_L g7236 ( 
.A(n_7147),
.B(n_6837),
.Y(n_7236)
);

OA21x2_ASAP7_75t_L g7237 ( 
.A1(n_7033),
.A2(n_5201),
.B(n_5195),
.Y(n_7237)
);

OR2x2_ASAP7_75t_L g7238 ( 
.A(n_7038),
.B(n_4883),
.Y(n_7238)
);

AND2x2_ASAP7_75t_L g7239 ( 
.A(n_7125),
.B(n_4636),
.Y(n_7239)
);

NOR2x1_ASAP7_75t_L g7240 ( 
.A(n_7042),
.B(n_4696),
.Y(n_7240)
);

AND2x2_ASAP7_75t_L g7241 ( 
.A(n_7071),
.B(n_4696),
.Y(n_7241)
);

INVx1_ASAP7_75t_L g7242 ( 
.A(n_7092),
.Y(n_7242)
);

OR2x2_ASAP7_75t_L g7243 ( 
.A(n_7023),
.B(n_4913),
.Y(n_7243)
);

INVx2_ASAP7_75t_L g7244 ( 
.A(n_7188),
.Y(n_7244)
);

OR2x6_ASAP7_75t_L g7245 ( 
.A(n_7059),
.B(n_4574),
.Y(n_7245)
);

AOI22xp33_ASAP7_75t_L g7246 ( 
.A1(n_7060),
.A2(n_5214),
.B1(n_5218),
.B2(n_5201),
.Y(n_7246)
);

INVx1_ASAP7_75t_L g7247 ( 
.A(n_7027),
.Y(n_7247)
);

INVx1_ASAP7_75t_L g7248 ( 
.A(n_7031),
.Y(n_7248)
);

INVx1_ASAP7_75t_L g7249 ( 
.A(n_7172),
.Y(n_7249)
);

INVx1_ASAP7_75t_L g7250 ( 
.A(n_7102),
.Y(n_7250)
);

AOI22xp33_ASAP7_75t_SL g7251 ( 
.A1(n_7070),
.A2(n_5145),
.B1(n_4939),
.B2(n_4937),
.Y(n_7251)
);

HB1xp67_ASAP7_75t_L g7252 ( 
.A(n_7128),
.Y(n_7252)
);

AND2x2_ASAP7_75t_L g7253 ( 
.A(n_7065),
.B(n_4696),
.Y(n_7253)
);

INVxp67_ASAP7_75t_L g7254 ( 
.A(n_7193),
.Y(n_7254)
);

NOR2x1_ASAP7_75t_L g7255 ( 
.A(n_7061),
.B(n_4844),
.Y(n_7255)
);

INVx3_ASAP7_75t_L g7256 ( 
.A(n_7116),
.Y(n_7256)
);

NAND2xp5_ASAP7_75t_L g7257 ( 
.A(n_7154),
.B(n_5238),
.Y(n_7257)
);

INVx5_ASAP7_75t_SL g7258 ( 
.A(n_7105),
.Y(n_7258)
);

OAI21xp33_ASAP7_75t_SL g7259 ( 
.A1(n_7030),
.A2(n_4844),
.B(n_4706),
.Y(n_7259)
);

AND2x4_ASAP7_75t_L g7260 ( 
.A(n_7132),
.B(n_4706),
.Y(n_7260)
);

OR2x2_ASAP7_75t_L g7261 ( 
.A(n_7110),
.B(n_4923),
.Y(n_7261)
);

INVx1_ASAP7_75t_L g7262 ( 
.A(n_7102),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_7117),
.Y(n_7263)
);

HB1xp67_ASAP7_75t_L g7264 ( 
.A(n_7141),
.Y(n_7264)
);

CKINVDCx16_ASAP7_75t_R g7265 ( 
.A(n_7143),
.Y(n_7265)
);

AOI22xp33_ASAP7_75t_L g7266 ( 
.A1(n_7121),
.A2(n_5218),
.B1(n_5224),
.B2(n_5214),
.Y(n_7266)
);

AND2x2_ASAP7_75t_L g7267 ( 
.A(n_7179),
.B(n_4706),
.Y(n_7267)
);

INVx4_ASAP7_75t_L g7268 ( 
.A(n_7046),
.Y(n_7268)
);

NAND2xp5_ASAP7_75t_L g7269 ( 
.A(n_7112),
.B(n_5244),
.Y(n_7269)
);

NOR2xp33_ASAP7_75t_L g7270 ( 
.A(n_7074),
.B(n_5224),
.Y(n_7270)
);

AND2x2_ASAP7_75t_L g7271 ( 
.A(n_7194),
.B(n_4844),
.Y(n_7271)
);

INVx3_ASAP7_75t_L g7272 ( 
.A(n_7116),
.Y(n_7272)
);

OR2x2_ASAP7_75t_L g7273 ( 
.A(n_7114),
.B(n_4925),
.Y(n_7273)
);

CKINVDCx20_ASAP7_75t_R g7274 ( 
.A(n_7137),
.Y(n_7274)
);

INVx2_ASAP7_75t_L g7275 ( 
.A(n_7113),
.Y(n_7275)
);

OR2x2_ASAP7_75t_L g7276 ( 
.A(n_7133),
.B(n_4925),
.Y(n_7276)
);

AND2x2_ASAP7_75t_L g7277 ( 
.A(n_7139),
.B(n_4844),
.Y(n_7277)
);

INVx1_ASAP7_75t_SL g7278 ( 
.A(n_7196),
.Y(n_7278)
);

AOI222xp33_ASAP7_75t_L g7279 ( 
.A1(n_7043),
.A2(n_5228),
.B1(n_5233),
.B2(n_5225),
.C1(n_5244),
.C2(n_5238),
.Y(n_7279)
);

INVx1_ASAP7_75t_L g7280 ( 
.A(n_7098),
.Y(n_7280)
);

NOR2xp33_ASAP7_75t_L g7281 ( 
.A(n_7145),
.B(n_5225),
.Y(n_7281)
);

INVx1_ASAP7_75t_L g7282 ( 
.A(n_7165),
.Y(n_7282)
);

NAND3xp33_ASAP7_75t_L g7283 ( 
.A(n_7151),
.B(n_5233),
.C(n_5228),
.Y(n_7283)
);

OR2x2_ASAP7_75t_L g7284 ( 
.A(n_7142),
.B(n_4870),
.Y(n_7284)
);

BUFx2_ASAP7_75t_L g7285 ( 
.A(n_7169),
.Y(n_7285)
);

NAND2xp5_ASAP7_75t_L g7286 ( 
.A(n_7168),
.B(n_7177),
.Y(n_7286)
);

NOR2x1p5_ASAP7_75t_L g7287 ( 
.A(n_7032),
.B(n_4406),
.Y(n_7287)
);

AND2x2_ASAP7_75t_L g7288 ( 
.A(n_7090),
.B(n_4870),
.Y(n_7288)
);

INVx1_ASAP7_75t_SL g7289 ( 
.A(n_7056),
.Y(n_7289)
);

INVx2_ASAP7_75t_SL g7290 ( 
.A(n_7099),
.Y(n_7290)
);

AND2x2_ASAP7_75t_L g7291 ( 
.A(n_7163),
.B(n_4870),
.Y(n_7291)
);

INVx1_ASAP7_75t_SL g7292 ( 
.A(n_7087),
.Y(n_7292)
);

OAI21x1_ASAP7_75t_L g7293 ( 
.A1(n_7066),
.A2(n_5250),
.B(n_5248),
.Y(n_7293)
);

NOR2xp33_ASAP7_75t_L g7294 ( 
.A(n_7054),
.B(n_7068),
.Y(n_7294)
);

OR2x2_ASAP7_75t_L g7295 ( 
.A(n_7184),
.B(n_4879),
.Y(n_7295)
);

NAND2xp5_ASAP7_75t_L g7296 ( 
.A(n_7185),
.B(n_5248),
.Y(n_7296)
);

INVx1_ASAP7_75t_L g7297 ( 
.A(n_7117),
.Y(n_7297)
);

AND2x4_ASAP7_75t_L g7298 ( 
.A(n_7186),
.B(n_4879),
.Y(n_7298)
);

INVx2_ASAP7_75t_L g7299 ( 
.A(n_7113),
.Y(n_7299)
);

INVx1_ASAP7_75t_L g7300 ( 
.A(n_7123),
.Y(n_7300)
);

NOR2x1p5_ASAP7_75t_L g7301 ( 
.A(n_7187),
.B(n_4123),
.Y(n_7301)
);

INVx1_ASAP7_75t_L g7302 ( 
.A(n_7096),
.Y(n_7302)
);

NAND2xp5_ASAP7_75t_L g7303 ( 
.A(n_7146),
.B(n_5250),
.Y(n_7303)
);

INVx1_ASAP7_75t_SL g7304 ( 
.A(n_7047),
.Y(n_7304)
);

AOI22xp5_ASAP7_75t_L g7305 ( 
.A1(n_7064),
.A2(n_5257),
.B1(n_5269),
.B2(n_5259),
.Y(n_7305)
);

INVx2_ASAP7_75t_L g7306 ( 
.A(n_7081),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_7096),
.Y(n_7307)
);

OR2x2_ASAP7_75t_L g7308 ( 
.A(n_7171),
.B(n_4879),
.Y(n_7308)
);

INVx1_ASAP7_75t_L g7309 ( 
.A(n_7097),
.Y(n_7309)
);

INVx1_ASAP7_75t_L g7310 ( 
.A(n_7097),
.Y(n_7310)
);

NAND2xp5_ASAP7_75t_L g7311 ( 
.A(n_7173),
.B(n_5257),
.Y(n_7311)
);

AOI31xp33_ASAP7_75t_L g7312 ( 
.A1(n_7176),
.A2(n_3998),
.A3(n_3991),
.B(n_4312),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_7122),
.Y(n_7313)
);

AND2x4_ASAP7_75t_SL g7314 ( 
.A(n_7167),
.B(n_3957),
.Y(n_7314)
);

NAND2xp5_ASAP7_75t_L g7315 ( 
.A(n_7111),
.B(n_5259),
.Y(n_7315)
);

INVx1_ASAP7_75t_L g7316 ( 
.A(n_7103),
.Y(n_7316)
);

INVx1_ASAP7_75t_L g7317 ( 
.A(n_7148),
.Y(n_7317)
);

INVx2_ASAP7_75t_L g7318 ( 
.A(n_7081),
.Y(n_7318)
);

INVx2_ASAP7_75t_L g7319 ( 
.A(n_7175),
.Y(n_7319)
);

AND2x2_ASAP7_75t_L g7320 ( 
.A(n_7131),
.B(n_4879),
.Y(n_7320)
);

AOI222xp33_ASAP7_75t_L g7321 ( 
.A1(n_7080),
.A2(n_7189),
.B1(n_7135),
.B2(n_7067),
.C1(n_7088),
.C2(n_7035),
.Y(n_7321)
);

AND2x2_ASAP7_75t_L g7322 ( 
.A(n_7058),
.B(n_4910),
.Y(n_7322)
);

CKINVDCx20_ASAP7_75t_R g7323 ( 
.A(n_7022),
.Y(n_7323)
);

INVx1_ASAP7_75t_SL g7324 ( 
.A(n_7140),
.Y(n_7324)
);

INVx1_ASAP7_75t_L g7325 ( 
.A(n_7170),
.Y(n_7325)
);

INVx1_ASAP7_75t_L g7326 ( 
.A(n_7127),
.Y(n_7326)
);

INVx2_ASAP7_75t_SL g7327 ( 
.A(n_7120),
.Y(n_7327)
);

OR2x2_ASAP7_75t_L g7328 ( 
.A(n_7108),
.B(n_4910),
.Y(n_7328)
);

AND3x1_ASAP7_75t_L g7329 ( 
.A(n_7045),
.B(n_4910),
.C(n_4176),
.Y(n_7329)
);

INVx2_ASAP7_75t_L g7330 ( 
.A(n_7175),
.Y(n_7330)
);

INVx1_ASAP7_75t_L g7331 ( 
.A(n_7130),
.Y(n_7331)
);

NAND2xp5_ASAP7_75t_L g7332 ( 
.A(n_7115),
.B(n_5269),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_7191),
.Y(n_7333)
);

INVx1_ASAP7_75t_L g7334 ( 
.A(n_7195),
.Y(n_7334)
);

BUFx3_ASAP7_75t_L g7335 ( 
.A(n_7048),
.Y(n_7335)
);

INVx1_ASAP7_75t_SL g7336 ( 
.A(n_7134),
.Y(n_7336)
);

INVx1_ASAP7_75t_L g7337 ( 
.A(n_7050),
.Y(n_7337)
);

INVx2_ASAP7_75t_L g7338 ( 
.A(n_7160),
.Y(n_7338)
);

NOR2xp33_ASAP7_75t_L g7339 ( 
.A(n_7077),
.B(n_7174),
.Y(n_7339)
);

AND2x2_ASAP7_75t_L g7340 ( 
.A(n_7051),
.B(n_4045),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_7073),
.Y(n_7341)
);

INVx1_ASAP7_75t_L g7342 ( 
.A(n_7083),
.Y(n_7342)
);

OR2x2_ASAP7_75t_L g7343 ( 
.A(n_7155),
.B(n_4584),
.Y(n_7343)
);

INVxp67_ASAP7_75t_L g7344 ( 
.A(n_7069),
.Y(n_7344)
);

AND2x2_ASAP7_75t_L g7345 ( 
.A(n_7084),
.B(n_4045),
.Y(n_7345)
);

INVx1_ASAP7_75t_L g7346 ( 
.A(n_7106),
.Y(n_7346)
);

INVx1_ASAP7_75t_L g7347 ( 
.A(n_7213),
.Y(n_7347)
);

AOI322xp5_ASAP7_75t_L g7348 ( 
.A1(n_7305),
.A2(n_7095),
.A3(n_7107),
.B1(n_7076),
.B2(n_7075),
.C1(n_7192),
.C2(n_7085),
.Y(n_7348)
);

OAI22xp5_ASAP7_75t_L g7349 ( 
.A1(n_7217),
.A2(n_7124),
.B1(n_7072),
.B2(n_7091),
.Y(n_7349)
);

INVx1_ASAP7_75t_L g7350 ( 
.A(n_7208),
.Y(n_7350)
);

AOI221x1_ASAP7_75t_L g7351 ( 
.A1(n_7232),
.A2(n_7197),
.B1(n_7129),
.B2(n_7144),
.C(n_7118),
.Y(n_7351)
);

INVx2_ASAP7_75t_L g7352 ( 
.A(n_7219),
.Y(n_7352)
);

INVx2_ASAP7_75t_L g7353 ( 
.A(n_7258),
.Y(n_7353)
);

HB1xp67_ASAP7_75t_L g7354 ( 
.A(n_7205),
.Y(n_7354)
);

OR2x6_ASAP7_75t_L g7355 ( 
.A(n_7285),
.B(n_7200),
.Y(n_7355)
);

AND2x2_ASAP7_75t_L g7356 ( 
.A(n_7201),
.B(n_7156),
.Y(n_7356)
);

INVx1_ASAP7_75t_L g7357 ( 
.A(n_7200),
.Y(n_7357)
);

INVx1_ASAP7_75t_L g7358 ( 
.A(n_7237),
.Y(n_7358)
);

INVx2_ASAP7_75t_L g7359 ( 
.A(n_7258),
.Y(n_7359)
);

INVxp67_ASAP7_75t_L g7360 ( 
.A(n_7221),
.Y(n_7360)
);

OAI21xp33_ASAP7_75t_L g7361 ( 
.A1(n_7304),
.A2(n_7079),
.B(n_7159),
.Y(n_7361)
);

AND2x2_ASAP7_75t_SL g7362 ( 
.A(n_7230),
.B(n_7136),
.Y(n_7362)
);

INVx1_ASAP7_75t_L g7363 ( 
.A(n_7237),
.Y(n_7363)
);

OAI21xp5_ASAP7_75t_L g7364 ( 
.A1(n_7218),
.A2(n_7226),
.B(n_7203),
.Y(n_7364)
);

INVx1_ASAP7_75t_L g7365 ( 
.A(n_7234),
.Y(n_7365)
);

AOI221xp5_ASAP7_75t_L g7366 ( 
.A1(n_7313),
.A2(n_7082),
.B1(n_7180),
.B2(n_7089),
.C(n_7101),
.Y(n_7366)
);

XOR2xp5_ASAP7_75t_L g7367 ( 
.A(n_7323),
.B(n_7178),
.Y(n_7367)
);

AOI22xp5_ASAP7_75t_L g7368 ( 
.A1(n_7225),
.A2(n_7149),
.B1(n_7153),
.B2(n_7150),
.Y(n_7368)
);

O2A1O1Ixp5_ASAP7_75t_L g7369 ( 
.A1(n_7268),
.A2(n_7181),
.B(n_7164),
.C(n_7093),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_7233),
.Y(n_7370)
);

INVx1_ASAP7_75t_L g7371 ( 
.A(n_7199),
.Y(n_7371)
);

AOI22xp5_ASAP7_75t_L g7372 ( 
.A1(n_7279),
.A2(n_5274),
.B1(n_5278),
.B2(n_5270),
.Y(n_7372)
);

AND2x4_ASAP7_75t_L g7373 ( 
.A(n_7220),
.B(n_5270),
.Y(n_7373)
);

NAND2xp5_ASAP7_75t_L g7374 ( 
.A(n_7265),
.B(n_7231),
.Y(n_7374)
);

OR2x2_ASAP7_75t_L g7375 ( 
.A(n_7227),
.B(n_7211),
.Y(n_7375)
);

AND2x2_ASAP7_75t_L g7376 ( 
.A(n_7214),
.B(n_7162),
.Y(n_7376)
);

NOR2xp33_ASAP7_75t_L g7377 ( 
.A(n_7268),
.B(n_5274),
.Y(n_7377)
);

INVx1_ASAP7_75t_L g7378 ( 
.A(n_7231),
.Y(n_7378)
);

AOI211xp5_ASAP7_75t_L g7379 ( 
.A1(n_7202),
.A2(n_4291),
.B(n_7158),
.C(n_7183),
.Y(n_7379)
);

AOI222xp33_ASAP7_75t_L g7380 ( 
.A1(n_7300),
.A2(n_7262),
.B1(n_7263),
.B2(n_7250),
.C1(n_7228),
.C2(n_7270),
.Y(n_7380)
);

AOI222xp33_ASAP7_75t_L g7381 ( 
.A1(n_7250),
.A2(n_5282),
.B1(n_5280),
.B2(n_5283),
.C1(n_5281),
.C2(n_5278),
.Y(n_7381)
);

INVx2_ASAP7_75t_L g7382 ( 
.A(n_7287),
.Y(n_7382)
);

NOR2xp33_ASAP7_75t_L g7383 ( 
.A(n_7292),
.B(n_7216),
.Y(n_7383)
);

INVx1_ASAP7_75t_L g7384 ( 
.A(n_7206),
.Y(n_7384)
);

INVx2_ASAP7_75t_SL g7385 ( 
.A(n_7335),
.Y(n_7385)
);

NAND2xp33_ASAP7_75t_SL g7386 ( 
.A(n_7274),
.B(n_3957),
.Y(n_7386)
);

INVx1_ASAP7_75t_L g7387 ( 
.A(n_7212),
.Y(n_7387)
);

AND2x2_ASAP7_75t_L g7388 ( 
.A(n_7215),
.B(n_3957),
.Y(n_7388)
);

INVx2_ASAP7_75t_L g7389 ( 
.A(n_7256),
.Y(n_7389)
);

NAND2xp5_ASAP7_75t_SL g7390 ( 
.A(n_7242),
.B(n_7207),
.Y(n_7390)
);

A2O1A1Ixp33_ASAP7_75t_L g7391 ( 
.A1(n_7293),
.A2(n_5281),
.B(n_5282),
.C(n_5280),
.Y(n_7391)
);

OAI32xp33_ASAP7_75t_L g7392 ( 
.A1(n_7259),
.A2(n_4179),
.A3(n_4176),
.B1(n_4186),
.B2(n_4102),
.Y(n_7392)
);

OAI21xp5_ASAP7_75t_L g7393 ( 
.A1(n_7198),
.A2(n_5063),
.B(n_5070),
.Y(n_7393)
);

NAND2xp5_ASAP7_75t_L g7394 ( 
.A(n_7324),
.B(n_5283),
.Y(n_7394)
);

INVx1_ASAP7_75t_L g7395 ( 
.A(n_7262),
.Y(n_7395)
);

AOI21xp5_ASAP7_75t_L g7396 ( 
.A1(n_7286),
.A2(n_5287),
.B(n_5292),
.Y(n_7396)
);

OAI221xp5_ASAP7_75t_L g7397 ( 
.A1(n_7321),
.A2(n_4186),
.B1(n_4179),
.B2(n_4102),
.C(n_5287),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_7263),
.Y(n_7398)
);

NAND2xp5_ASAP7_75t_SL g7399 ( 
.A(n_7290),
.B(n_3957),
.Y(n_7399)
);

AND2x2_ASAP7_75t_L g7400 ( 
.A(n_7278),
.B(n_3957),
.Y(n_7400)
);

O2A1O1Ixp33_ASAP7_75t_SL g7401 ( 
.A1(n_7252),
.A2(n_4586),
.B(n_4587),
.C(n_4584),
.Y(n_7401)
);

AOI221xp5_ASAP7_75t_L g7402 ( 
.A1(n_7275),
.A2(n_7299),
.B1(n_7306),
.B2(n_7318),
.C(n_7222),
.Y(n_7402)
);

INVx1_ASAP7_75t_L g7403 ( 
.A(n_7264),
.Y(n_7403)
);

AOI21xp33_ASAP7_75t_L g7404 ( 
.A1(n_7339),
.A2(n_4939),
.B(n_4937),
.Y(n_7404)
);

AOI22xp5_ASAP7_75t_L g7405 ( 
.A1(n_7224),
.A2(n_5185),
.B1(n_5176),
.B2(n_5292),
.Y(n_7405)
);

INVx1_ASAP7_75t_L g7406 ( 
.A(n_7256),
.Y(n_7406)
);

OAI22xp5_ASAP7_75t_SL g7407 ( 
.A1(n_7223),
.A2(n_3362),
.B1(n_3373),
.B2(n_3741),
.Y(n_7407)
);

NAND2xp5_ASAP7_75t_L g7408 ( 
.A(n_7336),
.B(n_5017),
.Y(n_7408)
);

OAI21xp33_ASAP7_75t_SL g7409 ( 
.A1(n_7294),
.A2(n_4585),
.B(n_4577),
.Y(n_7409)
);

OR2x2_ASAP7_75t_L g7410 ( 
.A(n_7229),
.B(n_5070),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_7272),
.Y(n_7411)
);

INVx2_ASAP7_75t_L g7412 ( 
.A(n_7272),
.Y(n_7412)
);

NOR2xp33_ASAP7_75t_L g7413 ( 
.A(n_7210),
.B(n_5295),
.Y(n_7413)
);

NAND3xp33_ASAP7_75t_SL g7414 ( 
.A(n_7289),
.B(n_5309),
.C(n_5301),
.Y(n_7414)
);

OAI21xp33_ASAP7_75t_SL g7415 ( 
.A1(n_7297),
.A2(n_4585),
.B(n_4577),
.Y(n_7415)
);

AND2x2_ASAP7_75t_L g7416 ( 
.A(n_7241),
.B(n_4015),
.Y(n_7416)
);

OR2x2_ASAP7_75t_L g7417 ( 
.A(n_7327),
.B(n_5103),
.Y(n_7417)
);

NAND2xp5_ASAP7_75t_L g7418 ( 
.A(n_7338),
.B(n_5017),
.Y(n_7418)
);

AOI22xp33_ASAP7_75t_L g7419 ( 
.A1(n_7251),
.A2(n_4939),
.B1(n_4937),
.B2(n_5295),
.Y(n_7419)
);

INVx1_ASAP7_75t_L g7420 ( 
.A(n_7302),
.Y(n_7420)
);

OAI221xp5_ASAP7_75t_L g7421 ( 
.A1(n_7244),
.A2(n_4186),
.B1(n_4102),
.B2(n_5309),
.C(n_5301),
.Y(n_7421)
);

OR2x2_ASAP7_75t_L g7422 ( 
.A(n_7280),
.B(n_5070),
.Y(n_7422)
);

INVx1_ASAP7_75t_L g7423 ( 
.A(n_7307),
.Y(n_7423)
);

INVx1_ASAP7_75t_L g7424 ( 
.A(n_7309),
.Y(n_7424)
);

AOI222xp33_ASAP7_75t_L g7425 ( 
.A1(n_7246),
.A2(n_5326),
.B1(n_5321),
.B2(n_5333),
.C1(n_5322),
.C2(n_5316),
.Y(n_7425)
);

AOI21xp33_ASAP7_75t_L g7426 ( 
.A1(n_7344),
.A2(n_4939),
.B(n_4937),
.Y(n_7426)
);

INVx2_ASAP7_75t_L g7427 ( 
.A(n_7340),
.Y(n_7427)
);

OAI22xp5_ASAP7_75t_L g7428 ( 
.A1(n_7248),
.A2(n_5316),
.B1(n_5322),
.B2(n_5321),
.Y(n_7428)
);

OAI221xp5_ASAP7_75t_L g7429 ( 
.A1(n_7235),
.A2(n_4186),
.B1(n_5333),
.B2(n_5337),
.C(n_5326),
.Y(n_7429)
);

INVx1_ASAP7_75t_L g7430 ( 
.A(n_7310),
.Y(n_7430)
);

INVx1_ASAP7_75t_L g7431 ( 
.A(n_7337),
.Y(n_7431)
);

NOR2xp33_ASAP7_75t_L g7432 ( 
.A(n_7249),
.B(n_5337),
.Y(n_7432)
);

NAND2xp5_ASAP7_75t_L g7433 ( 
.A(n_7326),
.B(n_5017),
.Y(n_7433)
);

A2O1A1Ixp33_ASAP7_75t_L g7434 ( 
.A1(n_7281),
.A2(n_5338),
.B(n_4505),
.C(n_4513),
.Y(n_7434)
);

AOI21xp5_ASAP7_75t_L g7435 ( 
.A1(n_7236),
.A2(n_5338),
.B(n_5063),
.Y(n_7435)
);

INVx1_ASAP7_75t_L g7436 ( 
.A(n_7337),
.Y(n_7436)
);

AND2x4_ASAP7_75t_L g7437 ( 
.A(n_7301),
.B(n_4123),
.Y(n_7437)
);

INVx1_ASAP7_75t_SL g7438 ( 
.A(n_7345),
.Y(n_7438)
);

INVx1_ASAP7_75t_L g7439 ( 
.A(n_7341),
.Y(n_7439)
);

AO22x1_ASAP7_75t_L g7440 ( 
.A1(n_7331),
.A2(n_4202),
.B1(n_4318),
.B2(n_4240),
.Y(n_7440)
);

NAND2xp5_ASAP7_75t_L g7441 ( 
.A(n_7316),
.B(n_5017),
.Y(n_7441)
);

AOI21xp5_ASAP7_75t_L g7442 ( 
.A1(n_7341),
.A2(n_5063),
.B(n_5070),
.Y(n_7442)
);

NOR2xp33_ASAP7_75t_L g7443 ( 
.A(n_7247),
.B(n_5020),
.Y(n_7443)
);

INVx1_ASAP7_75t_L g7444 ( 
.A(n_7342),
.Y(n_7444)
);

INVx1_ASAP7_75t_L g7445 ( 
.A(n_7342),
.Y(n_7445)
);

AOI221xp5_ASAP7_75t_L g7446 ( 
.A1(n_7315),
.A2(n_5185),
.B1(n_5176),
.B2(n_4526),
.C(n_4515),
.Y(n_7446)
);

NOR2xp33_ASAP7_75t_SL g7447 ( 
.A(n_7282),
.B(n_4096),
.Y(n_7447)
);

O2A1O1Ixp33_ASAP7_75t_L g7448 ( 
.A1(n_7204),
.A2(n_5185),
.B(n_5020),
.C(n_5063),
.Y(n_7448)
);

INVx1_ASAP7_75t_L g7449 ( 
.A(n_7209),
.Y(n_7449)
);

NAND2xp5_ASAP7_75t_L g7450 ( 
.A(n_7346),
.B(n_5020),
.Y(n_7450)
);

OAI22xp33_ASAP7_75t_L g7451 ( 
.A1(n_7269),
.A2(n_4515),
.B1(n_4526),
.B2(n_4508),
.Y(n_7451)
);

INVx1_ASAP7_75t_SL g7452 ( 
.A(n_7253),
.Y(n_7452)
);

AND2x2_ASAP7_75t_L g7453 ( 
.A(n_7322),
.B(n_7291),
.Y(n_7453)
);

INVx1_ASAP7_75t_L g7454 ( 
.A(n_7238),
.Y(n_7454)
);

NAND2xp5_ASAP7_75t_L g7455 ( 
.A(n_7346),
.B(n_5020),
.Y(n_7455)
);

INVx1_ASAP7_75t_SL g7456 ( 
.A(n_7314),
.Y(n_7456)
);

NAND2xp5_ASAP7_75t_L g7457 ( 
.A(n_7298),
.B(n_5103),
.Y(n_7457)
);

AOI222xp33_ASAP7_75t_L g7458 ( 
.A1(n_7332),
.A2(n_4804),
.B1(n_4652),
.B2(n_4645),
.C1(n_4653),
.C2(n_4647),
.Y(n_7458)
);

AOI22xp33_ASAP7_75t_L g7459 ( 
.A1(n_7319),
.A2(n_5103),
.B1(n_5336),
.B2(n_4804),
.Y(n_7459)
);

INVx1_ASAP7_75t_L g7460 ( 
.A(n_7261),
.Y(n_7460)
);

A2O1A1Ixp33_ASAP7_75t_L g7461 ( 
.A1(n_7303),
.A2(n_4645),
.B(n_4652),
.C(n_4630),
.Y(n_7461)
);

NAND4xp25_ASAP7_75t_L g7462 ( 
.A(n_7240),
.B(n_4181),
.C(n_4174),
.D(n_4157),
.Y(n_7462)
);

NAND2xp5_ASAP7_75t_SL g7463 ( 
.A(n_7298),
.B(n_7260),
.Y(n_7463)
);

AOI22xp33_ASAP7_75t_L g7464 ( 
.A1(n_7330),
.A2(n_5103),
.B1(n_5336),
.B2(n_4645),
.Y(n_7464)
);

INVx1_ASAP7_75t_SL g7465 ( 
.A(n_7296),
.Y(n_7465)
);

AND2x2_ASAP7_75t_L g7466 ( 
.A(n_7277),
.B(n_4015),
.Y(n_7466)
);

INVx1_ASAP7_75t_L g7467 ( 
.A(n_7273),
.Y(n_7467)
);

XNOR2x1_ASAP7_75t_L g7468 ( 
.A(n_7276),
.B(n_4574),
.Y(n_7468)
);

OAI32xp33_ASAP7_75t_L g7469 ( 
.A1(n_7284),
.A2(n_3991),
.A3(n_3760),
.B1(n_3741),
.B2(n_4181),
.Y(n_7469)
);

AOI22xp5_ASAP7_75t_L g7470 ( 
.A1(n_7329),
.A2(n_5342),
.B1(n_5241),
.B2(n_5320),
.Y(n_7470)
);

NAND2xp5_ASAP7_75t_SL g7471 ( 
.A(n_7260),
.B(n_4015),
.Y(n_7471)
);

NAND2xp5_ASAP7_75t_L g7472 ( 
.A(n_7317),
.B(n_5342),
.Y(n_7472)
);

AND2x2_ASAP7_75t_L g7473 ( 
.A(n_7239),
.B(n_4015),
.Y(n_7473)
);

NAND2xp5_ASAP7_75t_L g7474 ( 
.A(n_7325),
.B(n_5342),
.Y(n_7474)
);

OAI222xp33_ASAP7_75t_L g7475 ( 
.A1(n_7245),
.A2(n_4831),
.B1(n_4611),
.B2(n_4730),
.C1(n_4704),
.C2(n_4316),
.Y(n_7475)
);

OAI21xp33_ASAP7_75t_L g7476 ( 
.A1(n_7312),
.A2(n_4509),
.B(n_4044),
.Y(n_7476)
);

AOI221xp5_ASAP7_75t_L g7477 ( 
.A1(n_7283),
.A2(n_7334),
.B1(n_7333),
.B2(n_7257),
.C(n_7311),
.Y(n_7477)
);

NAND2xp5_ASAP7_75t_SL g7478 ( 
.A(n_7255),
.B(n_4015),
.Y(n_7478)
);

NOR2xp33_ASAP7_75t_L g7479 ( 
.A(n_7254),
.B(n_5342),
.Y(n_7479)
);

AOI221xp5_ASAP7_75t_L g7480 ( 
.A1(n_7266),
.A2(n_4652),
.B1(n_4653),
.B2(n_4647),
.C(n_4630),
.Y(n_7480)
);

NAND2xp5_ASAP7_75t_L g7481 ( 
.A(n_7288),
.B(n_4586),
.Y(n_7481)
);

NAND2xp5_ASAP7_75t_L g7482 ( 
.A(n_7354),
.B(n_7308),
.Y(n_7482)
);

AND2x2_ASAP7_75t_L g7483 ( 
.A(n_7362),
.B(n_7267),
.Y(n_7483)
);

NAND2xp5_ASAP7_75t_L g7484 ( 
.A(n_7352),
.B(n_7295),
.Y(n_7484)
);

OR2x2_ASAP7_75t_L g7485 ( 
.A(n_7374),
.B(n_7243),
.Y(n_7485)
);

NAND2xp5_ASAP7_75t_L g7486 ( 
.A(n_7356),
.B(n_7343),
.Y(n_7486)
);

AOI22xp5_ASAP7_75t_L g7487 ( 
.A1(n_7465),
.A2(n_7403),
.B1(n_7380),
.B2(n_7443),
.Y(n_7487)
);

INVx1_ASAP7_75t_L g7488 ( 
.A(n_7358),
.Y(n_7488)
);

BUFx3_ASAP7_75t_L g7489 ( 
.A(n_7347),
.Y(n_7489)
);

INVx1_ASAP7_75t_L g7490 ( 
.A(n_7363),
.Y(n_7490)
);

AOI221xp5_ASAP7_75t_L g7491 ( 
.A1(n_7349),
.A2(n_7435),
.B1(n_7419),
.B2(n_7409),
.C(n_7479),
.Y(n_7491)
);

AOI22xp5_ASAP7_75t_L g7492 ( 
.A1(n_7454),
.A2(n_7320),
.B1(n_7245),
.B2(n_7271),
.Y(n_7492)
);

OAI32xp33_ASAP7_75t_L g7493 ( 
.A1(n_7371),
.A2(n_7328),
.A3(n_3760),
.B1(n_3741),
.B2(n_4181),
.Y(n_7493)
);

AOI21xp33_ASAP7_75t_L g7494 ( 
.A1(n_7377),
.A2(n_5336),
.B(n_5320),
.Y(n_7494)
);

INVx2_ASAP7_75t_L g7495 ( 
.A(n_7355),
.Y(n_7495)
);

NAND2xp5_ASAP7_75t_L g7496 ( 
.A(n_7378),
.B(n_5241),
.Y(n_7496)
);

INVx1_ASAP7_75t_L g7497 ( 
.A(n_7355),
.Y(n_7497)
);

INVxp67_ASAP7_75t_L g7498 ( 
.A(n_7355),
.Y(n_7498)
);

AO21x1_ASAP7_75t_SL g7499 ( 
.A1(n_7350),
.A2(n_4590),
.B(n_4587),
.Y(n_7499)
);

INVx1_ASAP7_75t_SL g7500 ( 
.A(n_7375),
.Y(n_7500)
);

AOI221xp5_ASAP7_75t_L g7501 ( 
.A1(n_7409),
.A2(n_4653),
.B1(n_4655),
.B2(n_4647),
.C(n_4630),
.Y(n_7501)
);

OAI22xp33_ASAP7_75t_L g7502 ( 
.A1(n_7408),
.A2(n_5320),
.B1(n_5241),
.B2(n_4656),
.Y(n_7502)
);

OR2x2_ASAP7_75t_L g7503 ( 
.A(n_7389),
.B(n_5113),
.Y(n_7503)
);

AND2x2_ASAP7_75t_L g7504 ( 
.A(n_7364),
.B(n_4015),
.Y(n_7504)
);

AOI21xp5_ASAP7_75t_L g7505 ( 
.A1(n_7390),
.A2(n_7399),
.B(n_7386),
.Y(n_7505)
);

OAI22xp33_ASAP7_75t_L g7506 ( 
.A1(n_7365),
.A2(n_5320),
.B1(n_5241),
.B2(n_4656),
.Y(n_7506)
);

INVx1_ASAP7_75t_L g7507 ( 
.A(n_7412),
.Y(n_7507)
);

NAND2xp33_ASAP7_75t_SL g7508 ( 
.A(n_7385),
.B(n_4044),
.Y(n_7508)
);

INVx1_ASAP7_75t_L g7509 ( 
.A(n_7367),
.Y(n_7509)
);

AOI222xp33_ASAP7_75t_L g7510 ( 
.A1(n_7415),
.A2(n_4662),
.B1(n_4656),
.B2(n_4669),
.C1(n_4663),
.C2(n_4658),
.Y(n_7510)
);

INVx1_ASAP7_75t_L g7511 ( 
.A(n_7383),
.Y(n_7511)
);

OA22x2_ASAP7_75t_L g7512 ( 
.A1(n_7368),
.A2(n_4872),
.B1(n_4900),
.B2(n_4806),
.Y(n_7512)
);

INVx1_ASAP7_75t_L g7513 ( 
.A(n_7406),
.Y(n_7513)
);

AOI32xp33_ASAP7_75t_L g7514 ( 
.A1(n_7447),
.A2(n_4402),
.A3(n_4903),
.B1(n_4806),
.B2(n_4900),
.Y(n_7514)
);

NOR2xp33_ASAP7_75t_L g7515 ( 
.A(n_7360),
.B(n_4831),
.Y(n_7515)
);

INVx1_ASAP7_75t_L g7516 ( 
.A(n_7411),
.Y(n_7516)
);

NAND2x1_ASAP7_75t_SL g7517 ( 
.A(n_7373),
.B(n_4041),
.Y(n_7517)
);

INVx1_ASAP7_75t_L g7518 ( 
.A(n_7395),
.Y(n_7518)
);

NAND2xp5_ASAP7_75t_L g7519 ( 
.A(n_7400),
.B(n_4590),
.Y(n_7519)
);

NOR2xp33_ASAP7_75t_L g7520 ( 
.A(n_7438),
.B(n_4869),
.Y(n_7520)
);

INVxp67_ASAP7_75t_SL g7521 ( 
.A(n_7398),
.Y(n_7521)
);

AOI21xp33_ASAP7_75t_L g7522 ( 
.A1(n_7357),
.A2(n_4658),
.B(n_4655),
.Y(n_7522)
);

AND2x2_ASAP7_75t_L g7523 ( 
.A(n_7388),
.B(n_4044),
.Y(n_7523)
);

NAND2xp5_ASAP7_75t_L g7524 ( 
.A(n_7373),
.B(n_4591),
.Y(n_7524)
);

NOR2xp33_ASAP7_75t_L g7525 ( 
.A(n_7414),
.B(n_4869),
.Y(n_7525)
);

INVx1_ASAP7_75t_L g7526 ( 
.A(n_7353),
.Y(n_7526)
);

NAND2xp5_ASAP7_75t_L g7527 ( 
.A(n_7359),
.B(n_4591),
.Y(n_7527)
);

AOI322xp5_ASAP7_75t_L g7528 ( 
.A1(n_7361),
.A2(n_4663),
.A3(n_4658),
.B1(n_4667),
.B2(n_4669),
.C1(n_4662),
.C2(n_4655),
.Y(n_7528)
);

AND2x2_ASAP7_75t_L g7529 ( 
.A(n_7453),
.B(n_4044),
.Y(n_7529)
);

NAND2xp5_ASAP7_75t_L g7530 ( 
.A(n_7452),
.B(n_4594),
.Y(n_7530)
);

INVx1_ASAP7_75t_L g7531 ( 
.A(n_7431),
.Y(n_7531)
);

INVx1_ASAP7_75t_L g7532 ( 
.A(n_7436),
.Y(n_7532)
);

XNOR2xp5_ASAP7_75t_L g7533 ( 
.A(n_7402),
.B(n_4704),
.Y(n_7533)
);

AND2x4_ASAP7_75t_L g7534 ( 
.A(n_7460),
.B(n_4160),
.Y(n_7534)
);

INVx3_ASAP7_75t_L g7535 ( 
.A(n_7437),
.Y(n_7535)
);

NAND2xp5_ASAP7_75t_L g7536 ( 
.A(n_7467),
.B(n_4594),
.Y(n_7536)
);

INVxp67_ASAP7_75t_L g7537 ( 
.A(n_7413),
.Y(n_7537)
);

NAND2xp5_ASAP7_75t_L g7538 ( 
.A(n_7427),
.B(n_4595),
.Y(n_7538)
);

HB1xp67_ASAP7_75t_L g7539 ( 
.A(n_7439),
.Y(n_7539)
);

NOR2xp33_ASAP7_75t_L g7540 ( 
.A(n_7384),
.B(n_4889),
.Y(n_7540)
);

OR2x2_ASAP7_75t_L g7541 ( 
.A(n_7370),
.B(n_5113),
.Y(n_7541)
);

OAI22xp5_ASAP7_75t_L g7542 ( 
.A1(n_7382),
.A2(n_4595),
.B1(n_4608),
.B2(n_4606),
.Y(n_7542)
);

INVx1_ASAP7_75t_L g7543 ( 
.A(n_7444),
.Y(n_7543)
);

OAI22xp33_ASAP7_75t_L g7544 ( 
.A1(n_7418),
.A2(n_7422),
.B1(n_7397),
.B2(n_7441),
.Y(n_7544)
);

NOR2x1_ASAP7_75t_L g7545 ( 
.A(n_7445),
.B(n_7449),
.Y(n_7545)
);

INVx2_ASAP7_75t_L g7546 ( 
.A(n_7416),
.Y(n_7546)
);

INVx1_ASAP7_75t_L g7547 ( 
.A(n_7394),
.Y(n_7547)
);

INVx1_ASAP7_75t_L g7548 ( 
.A(n_7376),
.Y(n_7548)
);

NAND2xp5_ASAP7_75t_L g7549 ( 
.A(n_7432),
.B(n_4606),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7387),
.Y(n_7550)
);

NAND2xp5_ASAP7_75t_L g7551 ( 
.A(n_7420),
.B(n_4608),
.Y(n_7551)
);

INVx2_ASAP7_75t_L g7552 ( 
.A(n_7468),
.Y(n_7552)
);

NAND2xp5_ASAP7_75t_L g7553 ( 
.A(n_7423),
.B(n_7424),
.Y(n_7553)
);

AOI211xp5_ASAP7_75t_SL g7554 ( 
.A1(n_7430),
.A2(n_7477),
.B(n_7366),
.C(n_7379),
.Y(n_7554)
);

INVx1_ASAP7_75t_L g7555 ( 
.A(n_7410),
.Y(n_7555)
);

AOI21xp33_ASAP7_75t_L g7556 ( 
.A1(n_7472),
.A2(n_4663),
.B(n_4662),
.Y(n_7556)
);

XOR2xp5_ASAP7_75t_L g7557 ( 
.A(n_7456),
.B(n_4044),
.Y(n_7557)
);

NAND4xp25_ASAP7_75t_SL g7558 ( 
.A(n_7351),
.B(n_4402),
.C(n_4612),
.D(n_4609),
.Y(n_7558)
);

NAND3xp33_ASAP7_75t_L g7559 ( 
.A(n_7348),
.B(n_4415),
.C(n_4444),
.Y(n_7559)
);

INVx2_ASAP7_75t_L g7560 ( 
.A(n_7466),
.Y(n_7560)
);

NOR3xp33_ASAP7_75t_L g7561 ( 
.A(n_7404),
.B(n_3760),
.C(n_3741),
.Y(n_7561)
);

INVxp33_ASAP7_75t_L g7562 ( 
.A(n_7463),
.Y(n_7562)
);

NAND2xp5_ASAP7_75t_L g7563 ( 
.A(n_7396),
.B(n_4609),
.Y(n_7563)
);

NAND2xp5_ASAP7_75t_L g7564 ( 
.A(n_7474),
.B(n_4612),
.Y(n_7564)
);

OAI22xp5_ASAP7_75t_L g7565 ( 
.A1(n_7417),
.A2(n_4621),
.B1(n_4632),
.B2(n_4626),
.Y(n_7565)
);

OAI22xp5_ASAP7_75t_L g7566 ( 
.A1(n_7429),
.A2(n_4621),
.B1(n_4632),
.B2(n_4626),
.Y(n_7566)
);

OAI21xp5_ASAP7_75t_SL g7567 ( 
.A1(n_7433),
.A2(n_4045),
.B(n_4044),
.Y(n_7567)
);

NAND2xp5_ASAP7_75t_L g7568 ( 
.A(n_7473),
.B(n_4634),
.Y(n_7568)
);

INVx1_ASAP7_75t_L g7569 ( 
.A(n_7450),
.Y(n_7569)
);

NAND2xp5_ASAP7_75t_SL g7570 ( 
.A(n_7437),
.B(n_4045),
.Y(n_7570)
);

INVx1_ASAP7_75t_L g7571 ( 
.A(n_7455),
.Y(n_7571)
);

INVx1_ASAP7_75t_L g7572 ( 
.A(n_7401),
.Y(n_7572)
);

INVx1_ASAP7_75t_L g7573 ( 
.A(n_7481),
.Y(n_7573)
);

AND2x2_ASAP7_75t_L g7574 ( 
.A(n_7440),
.B(n_4045),
.Y(n_7574)
);

NAND2xp5_ASAP7_75t_L g7575 ( 
.A(n_7428),
.B(n_4634),
.Y(n_7575)
);

OAI22xp33_ASAP7_75t_L g7576 ( 
.A1(n_7457),
.A2(n_4669),
.B1(n_4667),
.B2(n_4817),
.Y(n_7576)
);

INVx1_ASAP7_75t_SL g7577 ( 
.A(n_7407),
.Y(n_7577)
);

AOI221xp5_ASAP7_75t_L g7578 ( 
.A1(n_7442),
.A2(n_4667),
.B1(n_4583),
.B2(n_4601),
.C(n_4600),
.Y(n_7578)
);

A2O1A1Ixp33_ASAP7_75t_L g7579 ( 
.A1(n_7415),
.A2(n_4583),
.B(n_4600),
.C(n_4589),
.Y(n_7579)
);

NAND2xp5_ASAP7_75t_L g7580 ( 
.A(n_7471),
.B(n_4635),
.Y(n_7580)
);

OAI22xp5_ASAP7_75t_L g7581 ( 
.A1(n_7421),
.A2(n_4635),
.B1(n_4648),
.B2(n_4638),
.Y(n_7581)
);

NAND2xp5_ASAP7_75t_L g7582 ( 
.A(n_7478),
.B(n_4638),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_7369),
.Y(n_7583)
);

OAI21xp33_ASAP7_75t_L g7584 ( 
.A1(n_7462),
.A2(n_4142),
.B(n_4045),
.Y(n_7584)
);

NAND2xp5_ASAP7_75t_L g7585 ( 
.A(n_7476),
.B(n_4648),
.Y(n_7585)
);

O2A1O1Ixp33_ASAP7_75t_SL g7586 ( 
.A1(n_7469),
.A2(n_4904),
.B(n_4902),
.C(n_4657),
.Y(n_7586)
);

AOI32xp33_ASAP7_75t_L g7587 ( 
.A1(n_7459),
.A2(n_4872),
.A3(n_4911),
.B1(n_4750),
.B2(n_3917),
.Y(n_7587)
);

NAND2xp5_ASAP7_75t_L g7588 ( 
.A(n_7372),
.B(n_4650),
.Y(n_7588)
);

OAI21xp5_ASAP7_75t_L g7589 ( 
.A1(n_7393),
.A2(n_4562),
.B(n_4750),
.Y(n_7589)
);

INVxp67_ASAP7_75t_L g7590 ( 
.A(n_7426),
.Y(n_7590)
);

NAND2xp5_ASAP7_75t_L g7591 ( 
.A(n_7391),
.B(n_7434),
.Y(n_7591)
);

OAI22xp5_ASAP7_75t_L g7592 ( 
.A1(n_7470),
.A2(n_4657),
.B1(n_4661),
.B2(n_4650),
.Y(n_7592)
);

OAI21xp33_ASAP7_75t_L g7593 ( 
.A1(n_7392),
.A2(n_4173),
.B(n_4142),
.Y(n_7593)
);

INVx1_ASAP7_75t_L g7594 ( 
.A(n_7381),
.Y(n_7594)
);

AND2x2_ASAP7_75t_L g7595 ( 
.A(n_7405),
.B(n_4142),
.Y(n_7595)
);

NAND2xp5_ASAP7_75t_L g7596 ( 
.A(n_7451),
.B(n_4661),
.Y(n_7596)
);

INVx2_ASAP7_75t_L g7597 ( 
.A(n_7517),
.Y(n_7597)
);

OAI22xp5_ASAP7_75t_L g7598 ( 
.A1(n_7500),
.A2(n_7464),
.B1(n_7446),
.B2(n_7448),
.Y(n_7598)
);

NOR2xp33_ASAP7_75t_L g7599 ( 
.A(n_7498),
.B(n_7475),
.Y(n_7599)
);

NOR2xp33_ASAP7_75t_L g7600 ( 
.A(n_7495),
.B(n_7461),
.Y(n_7600)
);

AND2x4_ASAP7_75t_L g7601 ( 
.A(n_7483),
.B(n_4123),
.Y(n_7601)
);

INVx2_ASAP7_75t_L g7602 ( 
.A(n_7485),
.Y(n_7602)
);

OR2x2_ASAP7_75t_L g7603 ( 
.A(n_7583),
.B(n_5113),
.Y(n_7603)
);

NAND2xp5_ASAP7_75t_L g7604 ( 
.A(n_7521),
.B(n_7425),
.Y(n_7604)
);

AND2x2_ASAP7_75t_L g7605 ( 
.A(n_7562),
.B(n_7458),
.Y(n_7605)
);

NOR2xp33_ASAP7_75t_L g7606 ( 
.A(n_7497),
.B(n_7480),
.Y(n_7606)
);

OR2x2_ASAP7_75t_L g7607 ( 
.A(n_7486),
.B(n_5113),
.Y(n_7607)
);

AND2x2_ASAP7_75t_L g7608 ( 
.A(n_7529),
.B(n_4142),
.Y(n_7608)
);

AND2x4_ASAP7_75t_L g7609 ( 
.A(n_7489),
.B(n_4160),
.Y(n_7609)
);

INVx1_ASAP7_75t_L g7610 ( 
.A(n_7539),
.Y(n_7610)
);

INVx1_ASAP7_75t_L g7611 ( 
.A(n_7488),
.Y(n_7611)
);

NOR2xp33_ASAP7_75t_L g7612 ( 
.A(n_7487),
.B(n_4871),
.Y(n_7612)
);

AOI222xp33_ASAP7_75t_L g7613 ( 
.A1(n_7559),
.A2(n_4605),
.B1(n_4589),
.B2(n_4616),
.C1(n_4607),
.C2(n_4601),
.Y(n_7613)
);

INVx1_ASAP7_75t_L g7614 ( 
.A(n_7490),
.Y(n_7614)
);

NAND2xp5_ASAP7_75t_L g7615 ( 
.A(n_7535),
.B(n_5113),
.Y(n_7615)
);

INVx1_ASAP7_75t_L g7616 ( 
.A(n_7507),
.Y(n_7616)
);

INVx2_ASAP7_75t_L g7617 ( 
.A(n_7535),
.Y(n_7617)
);

OR2x2_ASAP7_75t_L g7618 ( 
.A(n_7482),
.B(n_4666),
.Y(n_7618)
);

INVx1_ASAP7_75t_L g7619 ( 
.A(n_7545),
.Y(n_7619)
);

AND2x4_ASAP7_75t_L g7620 ( 
.A(n_7504),
.B(n_4160),
.Y(n_7620)
);

NAND2xp5_ASAP7_75t_L g7621 ( 
.A(n_7550),
.B(n_4666),
.Y(n_7621)
);

INVx2_ASAP7_75t_L g7622 ( 
.A(n_7523),
.Y(n_7622)
);

CKINVDCx16_ASAP7_75t_R g7623 ( 
.A(n_7487),
.Y(n_7623)
);

NAND2xp5_ASAP7_75t_L g7624 ( 
.A(n_7511),
.B(n_4670),
.Y(n_7624)
);

NAND2xp5_ASAP7_75t_L g7625 ( 
.A(n_7518),
.B(n_4670),
.Y(n_7625)
);

INVx1_ASAP7_75t_L g7626 ( 
.A(n_7553),
.Y(n_7626)
);

NOR2xp33_ASAP7_75t_L g7627 ( 
.A(n_7558),
.B(n_4871),
.Y(n_7627)
);

INVx1_ASAP7_75t_L g7628 ( 
.A(n_7509),
.Y(n_7628)
);

OR2x2_ASAP7_75t_L g7629 ( 
.A(n_7513),
.B(n_4673),
.Y(n_7629)
);

NAND2xp5_ASAP7_75t_L g7630 ( 
.A(n_7505),
.B(n_4673),
.Y(n_7630)
);

INVx1_ASAP7_75t_SL g7631 ( 
.A(n_7484),
.Y(n_7631)
);

AND2x2_ASAP7_75t_L g7632 ( 
.A(n_7534),
.B(n_4142),
.Y(n_7632)
);

HB1xp67_ASAP7_75t_L g7633 ( 
.A(n_7533),
.Y(n_7633)
);

NAND2xp5_ASAP7_75t_L g7634 ( 
.A(n_7554),
.B(n_4676),
.Y(n_7634)
);

INVx2_ASAP7_75t_L g7635 ( 
.A(n_7541),
.Y(n_7635)
);

NAND2x1_ASAP7_75t_SL g7636 ( 
.A(n_7492),
.B(n_4041),
.Y(n_7636)
);

INVx1_ASAP7_75t_L g7637 ( 
.A(n_7531),
.Y(n_7637)
);

NAND2xp5_ASAP7_75t_L g7638 ( 
.A(n_7532),
.B(n_4676),
.Y(n_7638)
);

INVx1_ASAP7_75t_L g7639 ( 
.A(n_7543),
.Y(n_7639)
);

OR2x2_ASAP7_75t_L g7640 ( 
.A(n_7516),
.B(n_4678),
.Y(n_7640)
);

OR2x2_ASAP7_75t_L g7641 ( 
.A(n_7546),
.B(n_4678),
.Y(n_7641)
);

INVx1_ASAP7_75t_SL g7642 ( 
.A(n_7526),
.Y(n_7642)
);

AND2x2_ASAP7_75t_L g7643 ( 
.A(n_7534),
.B(n_4268),
.Y(n_7643)
);

NOR2xp33_ASAP7_75t_L g7644 ( 
.A(n_7537),
.B(n_4880),
.Y(n_7644)
);

NAND2xp5_ASAP7_75t_L g7645 ( 
.A(n_7520),
.B(n_4680),
.Y(n_7645)
);

INVx2_ASAP7_75t_L g7646 ( 
.A(n_7560),
.Y(n_7646)
);

NAND2xp5_ASAP7_75t_L g7647 ( 
.A(n_7540),
.B(n_4680),
.Y(n_7647)
);

INVx1_ASAP7_75t_SL g7648 ( 
.A(n_7555),
.Y(n_7648)
);

INVx1_ASAP7_75t_L g7649 ( 
.A(n_7572),
.Y(n_7649)
);

INVx2_ASAP7_75t_SL g7650 ( 
.A(n_7574),
.Y(n_7650)
);

NOR2xp33_ASAP7_75t_L g7651 ( 
.A(n_7567),
.B(n_4880),
.Y(n_7651)
);

NAND2xp5_ASAP7_75t_L g7652 ( 
.A(n_7557),
.B(n_4681),
.Y(n_7652)
);

AOI22xp33_ASAP7_75t_L g7653 ( 
.A1(n_7594),
.A2(n_7569),
.B1(n_7571),
.B2(n_7552),
.Y(n_7653)
);

NAND2xp5_ASAP7_75t_L g7654 ( 
.A(n_7573),
.B(n_4681),
.Y(n_7654)
);

INVx1_ASAP7_75t_SL g7655 ( 
.A(n_7508),
.Y(n_7655)
);

INVx2_ASAP7_75t_L g7656 ( 
.A(n_7503),
.Y(n_7656)
);

AND2x2_ASAP7_75t_L g7657 ( 
.A(n_7548),
.B(n_4268),
.Y(n_7657)
);

AND2x2_ASAP7_75t_L g7658 ( 
.A(n_7492),
.B(n_4268),
.Y(n_7658)
);

INVx2_ASAP7_75t_SL g7659 ( 
.A(n_7570),
.Y(n_7659)
);

AND2x2_ASAP7_75t_L g7660 ( 
.A(n_7515),
.B(n_4268),
.Y(n_7660)
);

AND2x2_ASAP7_75t_L g7661 ( 
.A(n_7577),
.B(n_4268),
.Y(n_7661)
);

NAND2xp5_ASAP7_75t_L g7662 ( 
.A(n_7547),
.B(n_4682),
.Y(n_7662)
);

AOI22xp33_ASAP7_75t_L g7663 ( 
.A1(n_7590),
.A2(n_4607),
.B1(n_4616),
.B2(n_4605),
.Y(n_7663)
);

INVx1_ASAP7_75t_SL g7664 ( 
.A(n_7591),
.Y(n_7664)
);

INVxp67_ASAP7_75t_L g7665 ( 
.A(n_7496),
.Y(n_7665)
);

AND3x1_ASAP7_75t_L g7666 ( 
.A(n_7491),
.B(n_4684),
.C(n_4682),
.Y(n_7666)
);

NAND2xp33_ASAP7_75t_L g7667 ( 
.A(n_7527),
.B(n_4268),
.Y(n_7667)
);

INVx1_ASAP7_75t_L g7668 ( 
.A(n_7524),
.Y(n_7668)
);

INVx1_ASAP7_75t_L g7669 ( 
.A(n_7563),
.Y(n_7669)
);

AND2x2_ASAP7_75t_L g7670 ( 
.A(n_7512),
.B(n_4280),
.Y(n_7670)
);

AND2x2_ASAP7_75t_L g7671 ( 
.A(n_7584),
.B(n_4280),
.Y(n_7671)
);

INVx1_ASAP7_75t_L g7672 ( 
.A(n_7530),
.Y(n_7672)
);

INVxp67_ASAP7_75t_L g7673 ( 
.A(n_7551),
.Y(n_7673)
);

NAND2x1_ASAP7_75t_L g7674 ( 
.A(n_7595),
.B(n_4007),
.Y(n_7674)
);

NAND2xp5_ASAP7_75t_L g7675 ( 
.A(n_7525),
.B(n_4684),
.Y(n_7675)
);

AND2x2_ASAP7_75t_L g7676 ( 
.A(n_7499),
.B(n_4280),
.Y(n_7676)
);

AND2x2_ASAP7_75t_L g7677 ( 
.A(n_7561),
.B(n_7538),
.Y(n_7677)
);

NOR2xp33_ASAP7_75t_L g7678 ( 
.A(n_7544),
.B(n_7519),
.Y(n_7678)
);

NOR2xp33_ASAP7_75t_L g7679 ( 
.A(n_7549),
.B(n_4889),
.Y(n_7679)
);

NAND2xp5_ASAP7_75t_L g7680 ( 
.A(n_7568),
.B(n_7536),
.Y(n_7680)
);

INVx2_ASAP7_75t_L g7681 ( 
.A(n_7564),
.Y(n_7681)
);

AND2x2_ASAP7_75t_L g7682 ( 
.A(n_7493),
.B(n_7588),
.Y(n_7682)
);

INVx1_ASAP7_75t_L g7683 ( 
.A(n_7575),
.Y(n_7683)
);

INVxp67_ASAP7_75t_SL g7684 ( 
.A(n_7582),
.Y(n_7684)
);

OR2x2_ASAP7_75t_L g7685 ( 
.A(n_7585),
.B(n_4686),
.Y(n_7685)
);

AND2x2_ASAP7_75t_L g7686 ( 
.A(n_7580),
.B(n_4280),
.Y(n_7686)
);

AND2x2_ASAP7_75t_L g7687 ( 
.A(n_7593),
.B(n_4280),
.Y(n_7687)
);

AND2x4_ASAP7_75t_L g7688 ( 
.A(n_7596),
.B(n_4280),
.Y(n_7688)
);

NAND2x1_ASAP7_75t_SL g7689 ( 
.A(n_7586),
.B(n_4157),
.Y(n_7689)
);

NAND2xp5_ASAP7_75t_L g7690 ( 
.A(n_7528),
.B(n_4686),
.Y(n_7690)
);

NOR2xp33_ASAP7_75t_SL g7691 ( 
.A(n_7565),
.B(n_4096),
.Y(n_7691)
);

BUFx2_ASAP7_75t_L g7692 ( 
.A(n_7636),
.Y(n_7692)
);

NOR2xp33_ASAP7_75t_L g7693 ( 
.A(n_7623),
.B(n_7522),
.Y(n_7693)
);

INVx1_ASAP7_75t_L g7694 ( 
.A(n_7602),
.Y(n_7694)
);

OAI211xp5_ASAP7_75t_L g7695 ( 
.A1(n_7631),
.A2(n_7587),
.B(n_7514),
.C(n_7494),
.Y(n_7695)
);

INVx2_ASAP7_75t_L g7696 ( 
.A(n_7631),
.Y(n_7696)
);

INVx1_ASAP7_75t_L g7697 ( 
.A(n_7617),
.Y(n_7697)
);

NAND4xp25_ASAP7_75t_SL g7698 ( 
.A(n_7642),
.B(n_7589),
.C(n_7556),
.D(n_7510),
.Y(n_7698)
);

AOI221xp5_ASAP7_75t_L g7699 ( 
.A1(n_7598),
.A2(n_7648),
.B1(n_7599),
.B2(n_7665),
.C(n_7610),
.Y(n_7699)
);

NAND3xp33_ASAP7_75t_L g7700 ( 
.A(n_7619),
.B(n_7592),
.C(n_7566),
.Y(n_7700)
);

NOR2xp33_ASAP7_75t_L g7701 ( 
.A(n_7642),
.B(n_7576),
.Y(n_7701)
);

NAND3xp33_ASAP7_75t_L g7702 ( 
.A(n_7653),
.B(n_7581),
.C(n_7502),
.Y(n_7702)
);

OAI322xp33_ASAP7_75t_L g7703 ( 
.A1(n_7648),
.A2(n_7691),
.A3(n_7603),
.B1(n_7604),
.B2(n_7628),
.C1(n_7655),
.C2(n_7678),
.Y(n_7703)
);

OAI22xp33_ASAP7_75t_L g7704 ( 
.A1(n_7611),
.A2(n_7506),
.B1(n_7542),
.B2(n_7501),
.Y(n_7704)
);

NAND4xp25_ASAP7_75t_L g7705 ( 
.A(n_7664),
.B(n_7579),
.C(n_7578),
.D(n_4157),
.Y(n_7705)
);

INVx1_ASAP7_75t_L g7706 ( 
.A(n_7646),
.Y(n_7706)
);

INVx1_ASAP7_75t_L g7707 ( 
.A(n_7605),
.Y(n_7707)
);

NAND2xp5_ASAP7_75t_L g7708 ( 
.A(n_7676),
.B(n_4893),
.Y(n_7708)
);

AOI21xp5_ASAP7_75t_L g7709 ( 
.A1(n_7634),
.A2(n_4444),
.B(n_4690),
.Y(n_7709)
);

NAND2xp5_ASAP7_75t_L g7710 ( 
.A(n_7664),
.B(n_4893),
.Y(n_7710)
);

NAND4xp25_ASAP7_75t_L g7711 ( 
.A(n_7612),
.B(n_4157),
.C(n_3760),
.D(n_4401),
.Y(n_7711)
);

INVx1_ASAP7_75t_L g7712 ( 
.A(n_7616),
.Y(n_7712)
);

NOR2xp33_ASAP7_75t_L g7713 ( 
.A(n_7650),
.B(n_4892),
.Y(n_7713)
);

NOR3x1_ASAP7_75t_L g7714 ( 
.A(n_7659),
.B(n_4911),
.C(n_4620),
.Y(n_7714)
);

NOR3xp33_ASAP7_75t_L g7715 ( 
.A(n_7614),
.B(n_4625),
.C(n_4619),
.Y(n_7715)
);

NAND2xp5_ASAP7_75t_L g7716 ( 
.A(n_7658),
.B(n_4892),
.Y(n_7716)
);

NAND3xp33_ASAP7_75t_SL g7717 ( 
.A(n_7649),
.B(n_4203),
.C(n_4183),
.Y(n_7717)
);

NAND2xp5_ASAP7_75t_L g7718 ( 
.A(n_7670),
.B(n_4896),
.Y(n_7718)
);

OAI22xp5_ASAP7_75t_L g7719 ( 
.A1(n_7626),
.A2(n_4689),
.B1(n_4691),
.B2(n_4690),
.Y(n_7719)
);

INVx1_ASAP7_75t_L g7720 ( 
.A(n_7657),
.Y(n_7720)
);

NOR3x1_ASAP7_75t_L g7721 ( 
.A(n_7684),
.B(n_4620),
.C(n_3894),
.Y(n_7721)
);

NAND4xp25_ASAP7_75t_SL g7722 ( 
.A(n_7637),
.B(n_4691),
.C(n_4700),
.D(n_4689),
.Y(n_7722)
);

AND2x2_ASAP7_75t_L g7723 ( 
.A(n_7609),
.B(n_4142),
.Y(n_7723)
);

NAND2xp5_ASAP7_75t_SL g7724 ( 
.A(n_7601),
.B(n_4173),
.Y(n_7724)
);

INVx2_ASAP7_75t_SL g7725 ( 
.A(n_7609),
.Y(n_7725)
);

NOR2x1_ASAP7_75t_SL g7726 ( 
.A(n_7597),
.B(n_3242),
.Y(n_7726)
);

NAND3xp33_ASAP7_75t_L g7727 ( 
.A(n_7633),
.B(n_4415),
.C(n_4493),
.Y(n_7727)
);

AOI221x1_ASAP7_75t_L g7728 ( 
.A1(n_7639),
.A2(n_4700),
.B1(n_4715),
.B2(n_4712),
.C(n_4710),
.Y(n_7728)
);

AOI211xp5_ASAP7_75t_L g7729 ( 
.A1(n_7669),
.A2(n_3894),
.B(n_4241),
.C(n_4173),
.Y(n_7729)
);

AOI22xp5_ASAP7_75t_L g7730 ( 
.A1(n_7660),
.A2(n_4096),
.B1(n_4625),
.B2(n_4619),
.Y(n_7730)
);

OAI21xp5_ASAP7_75t_L g7731 ( 
.A1(n_7673),
.A2(n_7680),
.B(n_7681),
.Y(n_7731)
);

NOR2xp33_ASAP7_75t_SL g7732 ( 
.A(n_7622),
.B(n_4096),
.Y(n_7732)
);

NAND4xp25_ASAP7_75t_SL g7733 ( 
.A(n_7661),
.B(n_4712),
.C(n_4715),
.D(n_4710),
.Y(n_7733)
);

AOI221xp5_ASAP7_75t_SL g7734 ( 
.A1(n_7667),
.A2(n_4724),
.B1(n_4725),
.B2(n_4723),
.C(n_4719),
.Y(n_7734)
);

OR2x2_ASAP7_75t_L g7735 ( 
.A(n_7641),
.B(n_4415),
.Y(n_7735)
);

INVx1_ASAP7_75t_L g7736 ( 
.A(n_7615),
.Y(n_7736)
);

OAI22xp5_ASAP7_75t_L g7737 ( 
.A1(n_7666),
.A2(n_4723),
.B1(n_4724),
.B2(n_4719),
.Y(n_7737)
);

NAND3xp33_ASAP7_75t_SL g7738 ( 
.A(n_7600),
.B(n_4203),
.C(n_4693),
.Y(n_7738)
);

NAND3xp33_ASAP7_75t_L g7739 ( 
.A(n_7606),
.B(n_4415),
.C(n_4493),
.Y(n_7739)
);

AO22x2_ASAP7_75t_L g7740 ( 
.A1(n_7635),
.A2(n_4693),
.B1(n_4722),
.B2(n_4702),
.Y(n_7740)
);

NOR3xp33_ASAP7_75t_L g7741 ( 
.A(n_7656),
.B(n_4722),
.C(n_4702),
.Y(n_7741)
);

NAND3xp33_ASAP7_75t_SL g7742 ( 
.A(n_7682),
.B(n_4780),
.C(n_4778),
.Y(n_7742)
);

NOR2xp33_ASAP7_75t_SL g7743 ( 
.A(n_7672),
.B(n_4202),
.Y(n_7743)
);

NOR3xp33_ASAP7_75t_L g7744 ( 
.A(n_7668),
.B(n_4780),
.C(n_4778),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_7666),
.Y(n_7745)
);

NOR2xp67_ASAP7_75t_L g7746 ( 
.A(n_7601),
.B(n_4173),
.Y(n_7746)
);

INVx1_ASAP7_75t_L g7747 ( 
.A(n_7607),
.Y(n_7747)
);

NAND4xp25_ASAP7_75t_L g7748 ( 
.A(n_7683),
.B(n_3898),
.C(n_4012),
.D(n_4182),
.Y(n_7748)
);

NOR2xp67_ASAP7_75t_L g7749 ( 
.A(n_7629),
.B(n_4173),
.Y(n_7749)
);

OAI322xp33_ASAP7_75t_L g7750 ( 
.A1(n_7691),
.A2(n_4824),
.A3(n_4821),
.B1(n_4825),
.B2(n_4836),
.C1(n_4823),
.C2(n_4817),
.Y(n_7750)
);

NOR3xp33_ASAP7_75t_L g7751 ( 
.A(n_7677),
.B(n_4786),
.C(n_4782),
.Y(n_7751)
);

NOR3xp33_ASAP7_75t_SL g7752 ( 
.A(n_7630),
.B(n_7624),
.C(n_7621),
.Y(n_7752)
);

NAND4xp25_ASAP7_75t_L g7753 ( 
.A(n_7644),
.B(n_4012),
.C(n_4213),
.D(n_4182),
.Y(n_7753)
);

INVx2_ASAP7_75t_L g7754 ( 
.A(n_7689),
.Y(n_7754)
);

INVx1_ASAP7_75t_L g7755 ( 
.A(n_7640),
.Y(n_7755)
);

NAND2xp5_ASAP7_75t_SL g7756 ( 
.A(n_7688),
.B(n_4173),
.Y(n_7756)
);

NAND2xp5_ASAP7_75t_L g7757 ( 
.A(n_7686),
.B(n_4896),
.Y(n_7757)
);

AOI222xp33_ASAP7_75t_L g7758 ( 
.A1(n_7627),
.A2(n_4816),
.B1(n_4786),
.B2(n_4808),
.C1(n_4782),
.C2(n_4746),
.Y(n_7758)
);

INVx1_ASAP7_75t_L g7759 ( 
.A(n_7618),
.Y(n_7759)
);

INVx1_ASAP7_75t_L g7760 ( 
.A(n_7647),
.Y(n_7760)
);

NAND3xp33_ASAP7_75t_L g7761 ( 
.A(n_7674),
.B(n_4493),
.C(n_4808),
.Y(n_7761)
);

NAND2xp5_ASAP7_75t_L g7762 ( 
.A(n_7688),
.B(n_4897),
.Y(n_7762)
);

NOR3xp33_ASAP7_75t_L g7763 ( 
.A(n_7662),
.B(n_4816),
.C(n_4393),
.Y(n_7763)
);

NAND3xp33_ASAP7_75t_SL g7764 ( 
.A(n_7625),
.B(n_4737),
.C(n_4733),
.Y(n_7764)
);

INVx1_ASAP7_75t_L g7765 ( 
.A(n_7638),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_7654),
.Y(n_7766)
);

NOR2xp33_ASAP7_75t_L g7767 ( 
.A(n_7652),
.B(n_7679),
.Y(n_7767)
);

HB1xp67_ASAP7_75t_L g7768 ( 
.A(n_7632),
.Y(n_7768)
);

XNOR2xp5_ASAP7_75t_L g7769 ( 
.A(n_7620),
.B(n_4611),
.Y(n_7769)
);

NAND2xp5_ASAP7_75t_L g7770 ( 
.A(n_7608),
.B(n_4897),
.Y(n_7770)
);

INVx1_ASAP7_75t_L g7771 ( 
.A(n_7645),
.Y(n_7771)
);

NAND2xp5_ASAP7_75t_L g7772 ( 
.A(n_7643),
.B(n_4906),
.Y(n_7772)
);

INVx1_ASAP7_75t_L g7773 ( 
.A(n_7685),
.Y(n_7773)
);

NAND2xp5_ASAP7_75t_L g7774 ( 
.A(n_7746),
.B(n_7671),
.Y(n_7774)
);

NAND2xp5_ASAP7_75t_L g7775 ( 
.A(n_7696),
.B(n_7651),
.Y(n_7775)
);

NAND4xp25_ASAP7_75t_L g7776 ( 
.A(n_7699),
.B(n_7620),
.C(n_7687),
.D(n_7690),
.Y(n_7776)
);

NAND2xp5_ASAP7_75t_L g7777 ( 
.A(n_7749),
.B(n_7675),
.Y(n_7777)
);

NOR2xp33_ASAP7_75t_L g7778 ( 
.A(n_7707),
.B(n_7663),
.Y(n_7778)
);

NAND2xp5_ASAP7_75t_SL g7779 ( 
.A(n_7694),
.B(n_7613),
.Y(n_7779)
);

NAND2x1_ASAP7_75t_L g7780 ( 
.A(n_7692),
.B(n_4241),
.Y(n_7780)
);

AO21x1_ASAP7_75t_L g7781 ( 
.A1(n_7745),
.A2(n_4851),
.B(n_4847),
.Y(n_7781)
);

NOR2xp67_ASAP7_75t_SL g7782 ( 
.A(n_7706),
.B(n_3362),
.Y(n_7782)
);

NAND2xp5_ASAP7_75t_L g7783 ( 
.A(n_7693),
.B(n_4906),
.Y(n_7783)
);

NAND3xp33_ASAP7_75t_L g7784 ( 
.A(n_7701),
.B(n_4737),
.C(n_4733),
.Y(n_7784)
);

OAI321xp33_ASAP7_75t_L g7785 ( 
.A1(n_7695),
.A2(n_4393),
.A3(n_4385),
.B1(n_4372),
.B2(n_4316),
.C(n_3926),
.Y(n_7785)
);

NOR2x1_ASAP7_75t_SL g7786 ( 
.A(n_7754),
.B(n_3242),
.Y(n_7786)
);

AOI21xp33_ASAP7_75t_SL g7787 ( 
.A1(n_7702),
.A2(n_4444),
.B(n_4562),
.Y(n_7787)
);

AOI211xp5_ASAP7_75t_L g7788 ( 
.A1(n_7703),
.A2(n_4241),
.B(n_3820),
.C(n_4611),
.Y(n_7788)
);

AOI222xp33_ASAP7_75t_L g7789 ( 
.A1(n_7742),
.A2(n_4769),
.B1(n_4748),
.B2(n_4746),
.C1(n_4752),
.C2(n_4747),
.Y(n_7789)
);

NAND2xp5_ASAP7_75t_SL g7790 ( 
.A(n_7697),
.B(n_4241),
.Y(n_7790)
);

INVx1_ASAP7_75t_L g7791 ( 
.A(n_7768),
.Y(n_7791)
);

INVx2_ASAP7_75t_L g7792 ( 
.A(n_7725),
.Y(n_7792)
);

AOI22xp5_ASAP7_75t_L g7793 ( 
.A1(n_7698),
.A2(n_4742),
.B1(n_4748),
.B2(n_4747),
.Y(n_7793)
);

NAND2xp5_ASAP7_75t_L g7794 ( 
.A(n_7759),
.B(n_4493),
.Y(n_7794)
);

INVx1_ASAP7_75t_L g7795 ( 
.A(n_7712),
.Y(n_7795)
);

NAND3xp33_ASAP7_75t_L g7796 ( 
.A(n_7731),
.B(n_4752),
.C(n_4742),
.Y(n_7796)
);

NAND2xp5_ASAP7_75t_SL g7797 ( 
.A(n_7732),
.B(n_7743),
.Y(n_7797)
);

OR2x2_ASAP7_75t_L g7798 ( 
.A(n_7753),
.B(n_4444),
.Y(n_7798)
);

NAND4xp25_ASAP7_75t_L g7799 ( 
.A(n_7767),
.B(n_4730),
.C(n_4704),
.D(n_3956),
.Y(n_7799)
);

OAI22xp5_ASAP7_75t_L g7800 ( 
.A1(n_7720),
.A2(n_7700),
.B1(n_7766),
.B2(n_7765),
.Y(n_7800)
);

NAND4xp25_ASAP7_75t_L g7801 ( 
.A(n_7710),
.B(n_4730),
.C(n_4704),
.D(n_4048),
.Y(n_7801)
);

OAI21xp33_ASAP7_75t_L g7802 ( 
.A1(n_7752),
.A2(n_4241),
.B(n_4725),
.Y(n_7802)
);

NAND2xp5_ASAP7_75t_L g7803 ( 
.A(n_7755),
.B(n_4821),
.Y(n_7803)
);

AOI21xp5_ASAP7_75t_L g7804 ( 
.A1(n_7704),
.A2(n_4732),
.B(n_4727),
.Y(n_7804)
);

NOR2xp33_ASAP7_75t_SL g7805 ( 
.A(n_7773),
.B(n_4202),
.Y(n_7805)
);

AOI21xp33_ASAP7_75t_SL g7806 ( 
.A1(n_7747),
.A2(n_4177),
.B(n_4013),
.Y(n_7806)
);

INVx2_ASAP7_75t_SL g7807 ( 
.A(n_7723),
.Y(n_7807)
);

XNOR2xp5_ASAP7_75t_L g7808 ( 
.A(n_7769),
.B(n_4730),
.Y(n_7808)
);

HB1xp67_ASAP7_75t_L g7809 ( 
.A(n_7713),
.Y(n_7809)
);

AOI221xp5_ASAP7_75t_L g7810 ( 
.A1(n_7705),
.A2(n_4768),
.B1(n_4769),
.B2(n_4767),
.C(n_4759),
.Y(n_7810)
);

AOI22xp5_ASAP7_75t_L g7811 ( 
.A1(n_7718),
.A2(n_4767),
.B1(n_4768),
.B2(n_4759),
.Y(n_7811)
);

NAND2xp5_ASAP7_75t_L g7812 ( 
.A(n_7708),
.B(n_7771),
.Y(n_7812)
);

AOI211xp5_ASAP7_75t_L g7813 ( 
.A1(n_7760),
.A2(n_4241),
.B(n_4884),
.C(n_4882),
.Y(n_7813)
);

INVx1_ASAP7_75t_L g7814 ( 
.A(n_7757),
.Y(n_7814)
);

NAND2xp5_ASAP7_75t_SL g7815 ( 
.A(n_7736),
.B(n_4240),
.Y(n_7815)
);

NAND4xp25_ASAP7_75t_SL g7816 ( 
.A(n_7734),
.B(n_4732),
.C(n_4734),
.D(n_4727),
.Y(n_7816)
);

NAND2xp5_ASAP7_75t_L g7817 ( 
.A(n_7721),
.B(n_7756),
.Y(n_7817)
);

NAND2xp5_ASAP7_75t_L g7818 ( 
.A(n_7714),
.B(n_4823),
.Y(n_7818)
);

INVx1_ASAP7_75t_L g7819 ( 
.A(n_7762),
.Y(n_7819)
);

INVxp67_ASAP7_75t_SL g7820 ( 
.A(n_7726),
.Y(n_7820)
);

NAND4xp25_ASAP7_75t_L g7821 ( 
.A(n_7724),
.B(n_4074),
.C(n_4213),
.D(n_4182),
.Y(n_7821)
);

INVx1_ASAP7_75t_L g7822 ( 
.A(n_7716),
.Y(n_7822)
);

NAND3xp33_ASAP7_75t_L g7823 ( 
.A(n_7751),
.B(n_4774),
.C(n_4824),
.Y(n_7823)
);

NAND3xp33_ASAP7_75t_SL g7824 ( 
.A(n_7763),
.B(n_4774),
.C(n_4825),
.Y(n_7824)
);

OAI211xp5_ASAP7_75t_SL g7825 ( 
.A1(n_7709),
.A2(n_4740),
.B(n_4741),
.C(n_4734),
.Y(n_7825)
);

NOR2xp67_ASAP7_75t_L g7826 ( 
.A(n_7733),
.B(n_3242),
.Y(n_7826)
);

NAND2xp5_ASAP7_75t_L g7827 ( 
.A(n_7770),
.B(n_4836),
.Y(n_7827)
);

INVx1_ASAP7_75t_L g7828 ( 
.A(n_7772),
.Y(n_7828)
);

OAI211xp5_ASAP7_75t_L g7829 ( 
.A1(n_7711),
.A2(n_4014),
.B(n_3889),
.C(n_4740),
.Y(n_7829)
);

NAND3xp33_ASAP7_75t_L g7830 ( 
.A(n_7715),
.B(n_4854),
.C(n_4849),
.Y(n_7830)
);

NOR3xp33_ASAP7_75t_L g7831 ( 
.A(n_7738),
.B(n_4854),
.C(n_4849),
.Y(n_7831)
);

AOI211xp5_ASAP7_75t_L g7832 ( 
.A1(n_7737),
.A2(n_4109),
.B(n_4753),
.C(n_4741),
.Y(n_7832)
);

INVx2_ASAP7_75t_L g7833 ( 
.A(n_7735),
.Y(n_7833)
);

AOI22xp5_ASAP7_75t_L g7834 ( 
.A1(n_7727),
.A2(n_4318),
.B1(n_4343),
.B2(n_4240),
.Y(n_7834)
);

NOR2xp33_ASAP7_75t_L g7835 ( 
.A(n_7717),
.B(n_4240),
.Y(n_7835)
);

NAND2xp5_ASAP7_75t_L g7836 ( 
.A(n_7728),
.B(n_4753),
.Y(n_7836)
);

NAND2x1_ASAP7_75t_L g7837 ( 
.A(n_7730),
.B(n_4007),
.Y(n_7837)
);

NAND4xp25_ASAP7_75t_L g7838 ( 
.A(n_7748),
.B(n_4213),
.C(n_4361),
.D(n_3873),
.Y(n_7838)
);

NOR2xp33_ASAP7_75t_L g7839 ( 
.A(n_7739),
.B(n_4318),
.Y(n_7839)
);

NAND2xp5_ASAP7_75t_SL g7840 ( 
.A(n_7729),
.B(n_7761),
.Y(n_7840)
);

A2O1A1Ixp33_ASAP7_75t_L g7841 ( 
.A1(n_7741),
.A2(n_4761),
.B(n_4764),
.C(n_4756),
.Y(n_7841)
);

NAND4xp25_ASAP7_75t_L g7842 ( 
.A(n_7744),
.B(n_4213),
.C(n_3916),
.D(n_4178),
.Y(n_7842)
);

NOR3xp33_ASAP7_75t_L g7843 ( 
.A(n_7764),
.B(n_4083),
.C(n_4059),
.Y(n_7843)
);

OR2x2_ASAP7_75t_L g7844 ( 
.A(n_7722),
.B(n_4756),
.Y(n_7844)
);

NOR2xp33_ASAP7_75t_L g7845 ( 
.A(n_7750),
.B(n_4318),
.Y(n_7845)
);

INVx3_ASAP7_75t_L g7846 ( 
.A(n_7740),
.Y(n_7846)
);

BUFx12f_ASAP7_75t_L g7847 ( 
.A(n_7729),
.Y(n_7847)
);

NAND3xp33_ASAP7_75t_SL g7848 ( 
.A(n_7758),
.B(n_4405),
.C(n_4117),
.Y(n_7848)
);

AOI21xp5_ASAP7_75t_L g7849 ( 
.A1(n_7740),
.A2(n_4764),
.B(n_4761),
.Y(n_7849)
);

NAND2xp5_ASAP7_75t_L g7850 ( 
.A(n_7719),
.B(n_4766),
.Y(n_7850)
);

NAND3xp33_ASAP7_75t_L g7851 ( 
.A(n_7699),
.B(n_4343),
.C(n_3080),
.Y(n_7851)
);

INVx1_ASAP7_75t_SL g7852 ( 
.A(n_7696),
.Y(n_7852)
);

AND2x2_ASAP7_75t_L g7853 ( 
.A(n_7696),
.B(n_4766),
.Y(n_7853)
);

OAI21xp33_ASAP7_75t_L g7854 ( 
.A1(n_7694),
.A2(n_4771),
.B(n_4770),
.Y(n_7854)
);

AOI22xp33_ASAP7_75t_L g7855 ( 
.A1(n_7791),
.A2(n_4343),
.B1(n_4771),
.B2(n_4770),
.Y(n_7855)
);

AOI21xp5_ASAP7_75t_L g7856 ( 
.A1(n_7779),
.A2(n_4775),
.B(n_4773),
.Y(n_7856)
);

OAI22xp5_ASAP7_75t_L g7857 ( 
.A1(n_7852),
.A2(n_4775),
.B1(n_4781),
.B2(n_4773),
.Y(n_7857)
);

NAND2xp5_ASAP7_75t_SL g7858 ( 
.A(n_7792),
.B(n_4343),
.Y(n_7858)
);

XNOR2xp5_ASAP7_75t_L g7859 ( 
.A(n_7851),
.B(n_4372),
.Y(n_7859)
);

INVxp67_ASAP7_75t_L g7860 ( 
.A(n_7809),
.Y(n_7860)
);

BUFx2_ASAP7_75t_L g7861 ( 
.A(n_7847),
.Y(n_7861)
);

OAI21xp5_ASAP7_75t_SL g7862 ( 
.A1(n_7795),
.A2(n_4185),
.B(n_4013),
.Y(n_7862)
);

OAI22xp5_ASAP7_75t_L g7863 ( 
.A1(n_7820),
.A2(n_4783),
.B1(n_4790),
.B2(n_4781),
.Y(n_7863)
);

OAI221xp5_ASAP7_75t_L g7864 ( 
.A1(n_7780),
.A2(n_4088),
.B1(n_4007),
.B2(n_4790),
.C(n_4783),
.Y(n_7864)
);

NOR2x1_ASAP7_75t_L g7865 ( 
.A(n_7776),
.B(n_4791),
.Y(n_7865)
);

INVx1_ASAP7_75t_SL g7866 ( 
.A(n_7812),
.Y(n_7866)
);

AOI31xp33_ASAP7_75t_L g7867 ( 
.A1(n_7800),
.A2(n_3947),
.A3(n_3968),
.B(n_3900),
.Y(n_7867)
);

NAND4xp75_ASAP7_75t_L g7868 ( 
.A(n_7778),
.B(n_4258),
.C(n_4332),
.D(n_4177),
.Y(n_7868)
);

INVx1_ASAP7_75t_L g7869 ( 
.A(n_7846),
.Y(n_7869)
);

AOI22xp33_ASAP7_75t_L g7870 ( 
.A1(n_7833),
.A2(n_4792),
.B1(n_4797),
.B2(n_4791),
.Y(n_7870)
);

OAI21xp5_ASAP7_75t_L g7871 ( 
.A1(n_7817),
.A2(n_4797),
.B(n_4792),
.Y(n_7871)
);

INVx1_ASAP7_75t_L g7872 ( 
.A(n_7846),
.Y(n_7872)
);

INVx1_ASAP7_75t_L g7873 ( 
.A(n_7836),
.Y(n_7873)
);

XNOR2x1_ASAP7_75t_L g7874 ( 
.A(n_7775),
.B(n_4400),
.Y(n_7874)
);

INVx1_ASAP7_75t_L g7875 ( 
.A(n_7790),
.Y(n_7875)
);

INVx1_ASAP7_75t_L g7876 ( 
.A(n_7781),
.Y(n_7876)
);

INVx1_ASAP7_75t_L g7877 ( 
.A(n_7777),
.Y(n_7877)
);

NAND2xp5_ASAP7_75t_L g7878 ( 
.A(n_7808),
.B(n_4801),
.Y(n_7878)
);

XNOR2xp5_ASAP7_75t_L g7879 ( 
.A(n_7797),
.B(n_4400),
.Y(n_7879)
);

AOI211xp5_ASAP7_75t_L g7880 ( 
.A1(n_7807),
.A2(n_4904),
.B(n_4801),
.C(n_4815),
.Y(n_7880)
);

INVx1_ASAP7_75t_L g7881 ( 
.A(n_7774),
.Y(n_7881)
);

OAI22xp5_ASAP7_75t_SL g7882 ( 
.A1(n_7835),
.A2(n_3373),
.B1(n_3362),
.B2(n_4007),
.Y(n_7882)
);

INVx2_ASAP7_75t_L g7883 ( 
.A(n_7786),
.Y(n_7883)
);

NAND2xp5_ASAP7_75t_L g7884 ( 
.A(n_7845),
.B(n_7787),
.Y(n_7884)
);

AOI22xp5_ASAP7_75t_L g7885 ( 
.A1(n_7839),
.A2(n_4308),
.B1(n_4331),
.B2(n_4261),
.Y(n_7885)
);

XOR2xp5_ASAP7_75t_L g7886 ( 
.A(n_7815),
.B(n_3808),
.Y(n_7886)
);

INVx2_ASAP7_75t_SL g7887 ( 
.A(n_7853),
.Y(n_7887)
);

NOR2x1_ASAP7_75t_L g7888 ( 
.A(n_7819),
.B(n_4811),
.Y(n_7888)
);

HB1xp67_ASAP7_75t_L g7889 ( 
.A(n_7814),
.Y(n_7889)
);

INVx1_ASAP7_75t_L g7890 ( 
.A(n_7803),
.Y(n_7890)
);

INVx1_ASAP7_75t_L g7891 ( 
.A(n_7818),
.Y(n_7891)
);

NOR2x1_ASAP7_75t_L g7892 ( 
.A(n_7828),
.B(n_4811),
.Y(n_7892)
);

AOI21xp5_ASAP7_75t_L g7893 ( 
.A1(n_7840),
.A2(n_7805),
.B(n_7822),
.Y(n_7893)
);

AOI221xp5_ASAP7_75t_L g7894 ( 
.A1(n_7782),
.A2(n_7794),
.B1(n_7825),
.B2(n_7783),
.C(n_7804),
.Y(n_7894)
);

NAND2xp5_ASAP7_75t_L g7895 ( 
.A(n_7788),
.B(n_4815),
.Y(n_7895)
);

OAI21xp5_ASAP7_75t_SL g7896 ( 
.A1(n_7829),
.A2(n_7834),
.B(n_7802),
.Y(n_7896)
);

NAND2xp5_ASAP7_75t_L g7897 ( 
.A(n_7826),
.B(n_4818),
.Y(n_7897)
);

NAND2xp5_ASAP7_75t_SL g7898 ( 
.A(n_7785),
.B(n_4818),
.Y(n_7898)
);

AOI221xp5_ASAP7_75t_L g7899 ( 
.A1(n_7824),
.A2(n_4827),
.B1(n_4829),
.B2(n_4826),
.C(n_4820),
.Y(n_7899)
);

OAI21xp5_ASAP7_75t_L g7900 ( 
.A1(n_7798),
.A2(n_7796),
.B(n_7784),
.Y(n_7900)
);

AOI22xp5_ASAP7_75t_L g7901 ( 
.A1(n_7837),
.A2(n_4308),
.B1(n_4331),
.B2(n_4261),
.Y(n_7901)
);

INVx1_ASAP7_75t_L g7902 ( 
.A(n_7844),
.Y(n_7902)
);

INVx1_ASAP7_75t_SL g7903 ( 
.A(n_7827),
.Y(n_7903)
);

AOI222xp33_ASAP7_75t_L g7904 ( 
.A1(n_7848),
.A2(n_4829),
.B1(n_4820),
.B2(n_4830),
.C1(n_4827),
.C2(n_4826),
.Y(n_7904)
);

INVx1_ASAP7_75t_L g7905 ( 
.A(n_7850),
.Y(n_7905)
);

AOI22xp5_ASAP7_75t_L g7906 ( 
.A1(n_7854),
.A2(n_4308),
.B1(n_4331),
.B2(n_4261),
.Y(n_7906)
);

AOI32xp33_ASAP7_75t_L g7907 ( 
.A1(n_7813),
.A2(n_4832),
.A3(n_4834),
.B1(n_4833),
.B2(n_4830),
.Y(n_7907)
);

INVx1_ASAP7_75t_SL g7908 ( 
.A(n_7793),
.Y(n_7908)
);

INVx1_ASAP7_75t_L g7909 ( 
.A(n_7816),
.Y(n_7909)
);

AOI21xp5_ASAP7_75t_L g7910 ( 
.A1(n_7849),
.A2(n_4833),
.B(n_4832),
.Y(n_7910)
);

NAND2xp5_ASAP7_75t_SL g7911 ( 
.A(n_7813),
.B(n_4834),
.Y(n_7911)
);

OAI211xp5_ASAP7_75t_L g7912 ( 
.A1(n_7832),
.A2(n_4014),
.B(n_3889),
.C(n_4837),
.Y(n_7912)
);

NAND2xp5_ASAP7_75t_L g7913 ( 
.A(n_7841),
.B(n_4837),
.Y(n_7913)
);

XNOR2xp5_ASAP7_75t_L g7914 ( 
.A(n_7799),
.B(n_3926),
.Y(n_7914)
);

NOR3x1_ASAP7_75t_L g7915 ( 
.A(n_7821),
.B(n_3616),
.C(n_4838),
.Y(n_7915)
);

INVx1_ASAP7_75t_L g7916 ( 
.A(n_7831),
.Y(n_7916)
);

OAI221xp5_ASAP7_75t_L g7917 ( 
.A1(n_7838),
.A2(n_4088),
.B1(n_4843),
.B2(n_4847),
.C(n_4838),
.Y(n_7917)
);

INVx1_ASAP7_75t_L g7918 ( 
.A(n_7830),
.Y(n_7918)
);

OAI22xp33_ASAP7_75t_SL g7919 ( 
.A1(n_7866),
.A2(n_7811),
.B1(n_7823),
.B2(n_7801),
.Y(n_7919)
);

INVx1_ASAP7_75t_L g7920 ( 
.A(n_7889),
.Y(n_7920)
);

AO22x2_ASAP7_75t_L g7921 ( 
.A1(n_7876),
.A2(n_7843),
.B1(n_7806),
.B2(n_7842),
.Y(n_7921)
);

AOI22xp5_ASAP7_75t_L g7922 ( 
.A1(n_7881),
.A2(n_7810),
.B1(n_7789),
.B2(n_3117),
.Y(n_7922)
);

AOI211xp5_ASAP7_75t_SL g7923 ( 
.A1(n_7893),
.A2(n_3879),
.B(n_4851),
.C(n_4843),
.Y(n_7923)
);

INVx1_ASAP7_75t_L g7924 ( 
.A(n_7860),
.Y(n_7924)
);

INVx1_ASAP7_75t_L g7925 ( 
.A(n_7861),
.Y(n_7925)
);

OAI22xp5_ASAP7_75t_SL g7926 ( 
.A1(n_7883),
.A2(n_3373),
.B1(n_4088),
.B2(n_4261),
.Y(n_7926)
);

INVx1_ASAP7_75t_L g7927 ( 
.A(n_7873),
.Y(n_7927)
);

AOI22xp5_ASAP7_75t_L g7928 ( 
.A1(n_7877),
.A2(n_3117),
.B1(n_3118),
.B2(n_4308),
.Y(n_7928)
);

NOR2x1_ASAP7_75t_L g7929 ( 
.A(n_7875),
.B(n_4852),
.Y(n_7929)
);

INVx1_ASAP7_75t_L g7930 ( 
.A(n_7869),
.Y(n_7930)
);

NAND2xp5_ASAP7_75t_L g7931 ( 
.A(n_7872),
.B(n_4852),
.Y(n_7931)
);

INVx1_ASAP7_75t_L g7932 ( 
.A(n_7865),
.Y(n_7932)
);

AO22x2_ASAP7_75t_L g7933 ( 
.A1(n_7903),
.A2(n_7887),
.B1(n_7902),
.B2(n_7908),
.Y(n_7933)
);

NOR4xp25_ASAP7_75t_L g7934 ( 
.A(n_7891),
.B(n_7918),
.C(n_7916),
.D(n_7890),
.Y(n_7934)
);

NOR2xp33_ASAP7_75t_L g7935 ( 
.A(n_7884),
.B(n_4088),
.Y(n_7935)
);

NAND2xp5_ASAP7_75t_L g7936 ( 
.A(n_7914),
.B(n_4858),
.Y(n_7936)
);

INVx1_ASAP7_75t_L g7937 ( 
.A(n_7892),
.Y(n_7937)
);

INVx1_ASAP7_75t_L g7938 ( 
.A(n_7888),
.Y(n_7938)
);

INVx1_ASAP7_75t_L g7939 ( 
.A(n_7915),
.Y(n_7939)
);

AOI22xp5_ASAP7_75t_L g7940 ( 
.A1(n_7894),
.A2(n_3117),
.B1(n_3118),
.B2(n_4331),
.Y(n_7940)
);

INVx1_ASAP7_75t_L g7941 ( 
.A(n_7895),
.Y(n_7941)
);

AOI22xp5_ASAP7_75t_L g7942 ( 
.A1(n_7905),
.A2(n_3118),
.B1(n_4866),
.B2(n_4858),
.Y(n_7942)
);

NAND2xp5_ASAP7_75t_L g7943 ( 
.A(n_7879),
.B(n_4866),
.Y(n_7943)
);

NAND2xp5_ASAP7_75t_SL g7944 ( 
.A(n_7909),
.B(n_4867),
.Y(n_7944)
);

NOR4xp25_ASAP7_75t_L g7945 ( 
.A(n_7896),
.B(n_4873),
.C(n_4882),
.D(n_4867),
.Y(n_7945)
);

NAND2xp5_ASAP7_75t_L g7946 ( 
.A(n_7856),
.B(n_4873),
.Y(n_7946)
);

INVx1_ASAP7_75t_L g7947 ( 
.A(n_7897),
.Y(n_7947)
);

NOR2x1_ASAP7_75t_L g7948 ( 
.A(n_7858),
.B(n_4884),
.Y(n_7948)
);

AO22x2_ASAP7_75t_L g7949 ( 
.A1(n_7896),
.A2(n_4890),
.B1(n_4888),
.B2(n_3520),
.Y(n_7949)
);

AND2x2_ASAP7_75t_L g7950 ( 
.A(n_7874),
.B(n_4369),
.Y(n_7950)
);

AOI221xp5_ASAP7_75t_L g7951 ( 
.A1(n_7900),
.A2(n_4888),
.B1(n_4890),
.B2(n_4279),
.C(n_4266),
.Y(n_7951)
);

AND2x2_ASAP7_75t_L g7952 ( 
.A(n_7855),
.B(n_4369),
.Y(n_7952)
);

OAI22xp5_ASAP7_75t_L g7953 ( 
.A1(n_7886),
.A2(n_4014),
.B1(n_3889),
.B2(n_4212),
.Y(n_7953)
);

AOI22xp5_ASAP7_75t_L g7954 ( 
.A1(n_7898),
.A2(n_4307),
.B1(n_4369),
.B2(n_4177),
.Y(n_7954)
);

NOR4xp25_ASAP7_75t_L g7955 ( 
.A(n_7912),
.B(n_4335),
.C(n_4383),
.D(n_4354),
.Y(n_7955)
);

INVx1_ASAP7_75t_L g7956 ( 
.A(n_7878),
.Y(n_7956)
);

NAND2xp5_ASAP7_75t_L g7957 ( 
.A(n_7859),
.B(n_3992),
.Y(n_7957)
);

INVx1_ASAP7_75t_L g7958 ( 
.A(n_7911),
.Y(n_7958)
);

INVx2_ASAP7_75t_L g7959 ( 
.A(n_7913),
.Y(n_7959)
);

NAND2xp5_ASAP7_75t_L g7960 ( 
.A(n_7904),
.B(n_3992),
.Y(n_7960)
);

INVx1_ASAP7_75t_L g7961 ( 
.A(n_7871),
.Y(n_7961)
);

NAND2xp5_ASAP7_75t_SL g7962 ( 
.A(n_7882),
.B(n_4369),
.Y(n_7962)
);

OAI22xp5_ASAP7_75t_SL g7963 ( 
.A1(n_7901),
.A2(n_3857),
.B1(n_3625),
.B2(n_4377),
.Y(n_7963)
);

INVx1_ASAP7_75t_L g7964 ( 
.A(n_7910),
.Y(n_7964)
);

INVx1_ASAP7_75t_L g7965 ( 
.A(n_7857),
.Y(n_7965)
);

AOI22xp5_ASAP7_75t_L g7966 ( 
.A1(n_7885),
.A2(n_4307),
.B1(n_4177),
.B2(n_3992),
.Y(n_7966)
);

NAND2xp5_ASAP7_75t_L g7967 ( 
.A(n_7907),
.B(n_7870),
.Y(n_7967)
);

OA22x2_ASAP7_75t_L g7968 ( 
.A1(n_7906),
.A2(n_7862),
.B1(n_7863),
.B2(n_7917),
.Y(n_7968)
);

NAND2xp5_ASAP7_75t_L g7969 ( 
.A(n_7899),
.B(n_4258),
.Y(n_7969)
);

NAND2xp5_ASAP7_75t_L g7970 ( 
.A(n_7920),
.B(n_7880),
.Y(n_7970)
);

AOI21xp5_ASAP7_75t_L g7971 ( 
.A1(n_7925),
.A2(n_7864),
.B(n_7880),
.Y(n_7971)
);

AOI31xp33_ASAP7_75t_L g7972 ( 
.A1(n_7924),
.A2(n_7867),
.A3(n_7868),
.B(n_4185),
.Y(n_7972)
);

NAND2xp33_ASAP7_75t_SL g7973 ( 
.A(n_7932),
.B(n_3616),
.Y(n_7973)
);

NAND3xp33_ASAP7_75t_L g7974 ( 
.A(n_7930),
.B(n_4332),
.C(n_4258),
.Y(n_7974)
);

AND2x2_ASAP7_75t_L g7975 ( 
.A(n_7933),
.B(n_7950),
.Y(n_7975)
);

INVx1_ASAP7_75t_L g7976 ( 
.A(n_7933),
.Y(n_7976)
);

INVxp67_ASAP7_75t_L g7977 ( 
.A(n_7927),
.Y(n_7977)
);

INVx1_ASAP7_75t_L g7978 ( 
.A(n_7937),
.Y(n_7978)
);

NOR2xp67_ASAP7_75t_L g7979 ( 
.A(n_7938),
.B(n_3856),
.Y(n_7979)
);

AOI21xp5_ASAP7_75t_L g7980 ( 
.A1(n_7919),
.A2(n_4014),
.B(n_3889),
.Y(n_7980)
);

NAND2xp5_ASAP7_75t_L g7981 ( 
.A(n_7934),
.B(n_4258),
.Y(n_7981)
);

AND2x4_ASAP7_75t_L g7982 ( 
.A(n_7929),
.B(n_4307),
.Y(n_7982)
);

NAND2xp5_ASAP7_75t_L g7983 ( 
.A(n_7947),
.B(n_4332),
.Y(n_7983)
);

INVx1_ASAP7_75t_L g7984 ( 
.A(n_7921),
.Y(n_7984)
);

INVx1_ASAP7_75t_L g7985 ( 
.A(n_7921),
.Y(n_7985)
);

NAND2x1_ASAP7_75t_SL g7986 ( 
.A(n_7958),
.B(n_4352),
.Y(n_7986)
);

NOR2x1_ASAP7_75t_L g7987 ( 
.A(n_7964),
.B(n_4377),
.Y(n_7987)
);

NOR3xp33_ASAP7_75t_L g7988 ( 
.A(n_7956),
.B(n_3945),
.C(n_4366),
.Y(n_7988)
);

NAND2xp5_ASAP7_75t_L g7989 ( 
.A(n_7939),
.B(n_4332),
.Y(n_7989)
);

NOR3xp33_ASAP7_75t_L g7990 ( 
.A(n_7941),
.B(n_3845),
.C(n_3858),
.Y(n_7990)
);

AOI221xp5_ASAP7_75t_L g7991 ( 
.A1(n_7935),
.A2(n_4307),
.B1(n_3836),
.B2(n_3825),
.C(n_4354),
.Y(n_7991)
);

INVx2_ASAP7_75t_L g7992 ( 
.A(n_7959),
.Y(n_7992)
);

NOR2xp67_ASAP7_75t_L g7993 ( 
.A(n_7961),
.B(n_7965),
.Y(n_7993)
);

OR2x2_ASAP7_75t_L g7994 ( 
.A(n_7957),
.B(n_7960),
.Y(n_7994)
);

NAND2xp5_ASAP7_75t_L g7995 ( 
.A(n_7922),
.B(n_7952),
.Y(n_7995)
);

NAND2xp5_ASAP7_75t_L g7996 ( 
.A(n_7948),
.B(n_4357),
.Y(n_7996)
);

AOI21xp5_ASAP7_75t_L g7997 ( 
.A1(n_7967),
.A2(n_7944),
.B(n_7931),
.Y(n_7997)
);

NAND2xp5_ASAP7_75t_L g7998 ( 
.A(n_7936),
.B(n_4357),
.Y(n_7998)
);

OR2x2_ASAP7_75t_L g7999 ( 
.A(n_7955),
.B(n_3520),
.Y(n_7999)
);

NAND2xp5_ASAP7_75t_L g8000 ( 
.A(n_7946),
.B(n_4357),
.Y(n_8000)
);

NOR2x1_ASAP7_75t_L g8001 ( 
.A(n_7962),
.B(n_4377),
.Y(n_8001)
);

NAND2xp5_ASAP7_75t_L g8002 ( 
.A(n_7943),
.B(n_4357),
.Y(n_8002)
);

AOI22xp33_ASAP7_75t_SL g8003 ( 
.A1(n_7968),
.A2(n_3889),
.B1(n_4014),
.B2(n_3881),
.Y(n_8003)
);

NOR2x1_ASAP7_75t_L g8004 ( 
.A(n_7969),
.B(n_4377),
.Y(n_8004)
);

NAND3xp33_ASAP7_75t_L g8005 ( 
.A(n_7940),
.B(n_3926),
.C(n_4242),
.Y(n_8005)
);

INVx1_ASAP7_75t_L g8006 ( 
.A(n_7949),
.Y(n_8006)
);

INVx1_ASAP7_75t_L g8007 ( 
.A(n_7949),
.Y(n_8007)
);

NAND2xp5_ASAP7_75t_L g8008 ( 
.A(n_7945),
.B(n_4368),
.Y(n_8008)
);

OAI22xp5_ASAP7_75t_L g8009 ( 
.A1(n_7984),
.A2(n_7954),
.B1(n_7928),
.B2(n_7926),
.Y(n_8009)
);

OR2x6_ASAP7_75t_L g8010 ( 
.A(n_7976),
.B(n_7953),
.Y(n_8010)
);

NAND4xp25_ASAP7_75t_L g8011 ( 
.A(n_7993),
.B(n_7923),
.C(n_7942),
.D(n_7951),
.Y(n_8011)
);

NOR3xp33_ASAP7_75t_L g8012 ( 
.A(n_7985),
.B(n_7963),
.C(n_7966),
.Y(n_8012)
);

HB1xp67_ASAP7_75t_L g8013 ( 
.A(n_7975),
.Y(n_8013)
);

NOR2x1_ASAP7_75t_L g8014 ( 
.A(n_7978),
.B(n_4316),
.Y(n_8014)
);

NAND3x1_ASAP7_75t_L g8015 ( 
.A(n_7970),
.B(n_3853),
.C(n_4355),
.Y(n_8015)
);

NOR3xp33_ASAP7_75t_L g8016 ( 
.A(n_7977),
.B(n_3798),
.C(n_3785),
.Y(n_8016)
);

NOR2x1_ASAP7_75t_L g8017 ( 
.A(n_8006),
.B(n_3881),
.Y(n_8017)
);

INVx2_ASAP7_75t_L g8018 ( 
.A(n_7986),
.Y(n_8018)
);

NAND3xp33_ASAP7_75t_L g8019 ( 
.A(n_7992),
.B(n_4269),
.C(n_4256),
.Y(n_8019)
);

INVx2_ASAP7_75t_L g8020 ( 
.A(n_8007),
.Y(n_8020)
);

NAND4xp75_ASAP7_75t_L g8021 ( 
.A(n_7997),
.B(n_4387),
.C(n_4368),
.D(n_3862),
.Y(n_8021)
);

INVx1_ASAP7_75t_L g8022 ( 
.A(n_7981),
.Y(n_8022)
);

AND4x1_ASAP7_75t_L g8023 ( 
.A(n_7971),
.B(n_3850),
.C(n_3843),
.D(n_3775),
.Y(n_8023)
);

INVxp33_ASAP7_75t_L g8024 ( 
.A(n_7995),
.Y(n_8024)
);

OR3x1_ASAP7_75t_L g8025 ( 
.A(n_7973),
.B(n_8003),
.C(n_7980),
.Y(n_8025)
);

HB1xp67_ASAP7_75t_L g8026 ( 
.A(n_7994),
.Y(n_8026)
);

NAND4xp25_ASAP7_75t_L g8027 ( 
.A(n_8001),
.B(n_4210),
.C(n_4219),
.D(n_4200),
.Y(n_8027)
);

NOR3xp33_ASAP7_75t_L g8028 ( 
.A(n_7972),
.B(n_3891),
.C(n_3868),
.Y(n_8028)
);

HB1xp67_ASAP7_75t_L g8029 ( 
.A(n_7982),
.Y(n_8029)
);

OAI21xp5_ASAP7_75t_L g8030 ( 
.A1(n_7989),
.A2(n_3610),
.B(n_3499),
.Y(n_8030)
);

NOR3xp33_ASAP7_75t_L g8031 ( 
.A(n_8004),
.B(n_7983),
.C(n_7987),
.Y(n_8031)
);

INVx1_ASAP7_75t_SL g8032 ( 
.A(n_7982),
.Y(n_8032)
);

NOR2x1_ASAP7_75t_L g8033 ( 
.A(n_7999),
.B(n_3639),
.Y(n_8033)
);

OAI211xp5_ASAP7_75t_SL g8034 ( 
.A1(n_7998),
.A2(n_4079),
.B(n_4113),
.C(n_4228),
.Y(n_8034)
);

NAND3xp33_ASAP7_75t_SL g8035 ( 
.A(n_8000),
.B(n_4405),
.C(n_4185),
.Y(n_8035)
);

NOR2xp33_ASAP7_75t_L g8036 ( 
.A(n_8008),
.B(n_3527),
.Y(n_8036)
);

NAND4xp25_ASAP7_75t_SL g8037 ( 
.A(n_7996),
.B(n_3853),
.C(n_4356),
.D(n_4355),
.Y(n_8037)
);

AND2x2_ASAP7_75t_L g8038 ( 
.A(n_7979),
.B(n_3918),
.Y(n_8038)
);

NOR3xp33_ASAP7_75t_L g8039 ( 
.A(n_8002),
.B(n_3610),
.C(n_3838),
.Y(n_8039)
);

AND2x4_ASAP7_75t_L g8040 ( 
.A(n_8005),
.B(n_3574),
.Y(n_8040)
);

NAND3xp33_ASAP7_75t_SL g8041 ( 
.A(n_7988),
.B(n_7990),
.C(n_7974),
.Y(n_8041)
);

NOR4xp25_ASAP7_75t_L g8042 ( 
.A(n_7991),
.B(n_4356),
.C(n_4365),
.D(n_4358),
.Y(n_8042)
);

OR2x2_ASAP7_75t_L g8043 ( 
.A(n_7976),
.B(n_4845),
.Y(n_8043)
);

NOR3xp33_ASAP7_75t_L g8044 ( 
.A(n_7976),
.B(n_3895),
.C(n_3838),
.Y(n_8044)
);

NOR3xp33_ASAP7_75t_L g8045 ( 
.A(n_8013),
.B(n_3260),
.C(n_3245),
.Y(n_8045)
);

INVx1_ASAP7_75t_L g8046 ( 
.A(n_8026),
.Y(n_8046)
);

NOR2x1_ASAP7_75t_L g8047 ( 
.A(n_8020),
.B(n_3639),
.Y(n_8047)
);

NAND4xp75_ASAP7_75t_L g8048 ( 
.A(n_8022),
.B(n_4387),
.C(n_4368),
.D(n_3834),
.Y(n_8048)
);

AND2x4_ASAP7_75t_L g8049 ( 
.A(n_8029),
.B(n_8032),
.Y(n_8049)
);

OAI22xp5_ASAP7_75t_L g8050 ( 
.A1(n_8024),
.A2(n_4365),
.B1(n_4376),
.B2(n_4358),
.Y(n_8050)
);

NOR2xp33_ASAP7_75t_L g8051 ( 
.A(n_8018),
.B(n_3527),
.Y(n_8051)
);

AND2x2_ASAP7_75t_L g8052 ( 
.A(n_8033),
.B(n_3918),
.Y(n_8052)
);

INVx1_ASAP7_75t_L g8053 ( 
.A(n_8017),
.Y(n_8053)
);

AOI22xp33_ASAP7_75t_L g8054 ( 
.A1(n_8031),
.A2(n_4387),
.B1(n_4368),
.B2(n_3634),
.Y(n_8054)
);

OR2x2_ASAP7_75t_L g8055 ( 
.A(n_8011),
.B(n_4845),
.Y(n_8055)
);

INVx1_ASAP7_75t_L g8056 ( 
.A(n_8043),
.Y(n_8056)
);

NAND2xp5_ASAP7_75t_L g8057 ( 
.A(n_8038),
.B(n_4387),
.Y(n_8057)
);

AOI221xp5_ASAP7_75t_L g8058 ( 
.A1(n_8009),
.A2(n_4380),
.B1(n_4384),
.B2(n_4378),
.C(n_4376),
.Y(n_8058)
);

AOI21xp5_ASAP7_75t_L g8059 ( 
.A1(n_8010),
.A2(n_4133),
.B(n_3743),
.Y(n_8059)
);

NOR3xp33_ASAP7_75t_L g8060 ( 
.A(n_8012),
.B(n_3260),
.C(n_3245),
.Y(n_8060)
);

INVx1_ASAP7_75t_L g8061 ( 
.A(n_8025),
.Y(n_8061)
);

NAND2xp5_ASAP7_75t_L g8062 ( 
.A(n_8036),
.B(n_4845),
.Y(n_8062)
);

NOR2x1_ASAP7_75t_L g8063 ( 
.A(n_8010),
.B(n_3786),
.Y(n_8063)
);

NAND4xp75_ASAP7_75t_L g8064 ( 
.A(n_8014),
.B(n_4380),
.C(n_4384),
.D(n_4378),
.Y(n_8064)
);

NAND3xp33_ASAP7_75t_SL g8065 ( 
.A(n_8044),
.B(n_8016),
.C(n_8028),
.Y(n_8065)
);

AND2x2_ASAP7_75t_L g8066 ( 
.A(n_8040),
.B(n_3918),
.Y(n_8066)
);

INVx1_ASAP7_75t_L g8067 ( 
.A(n_8041),
.Y(n_8067)
);

AOI22xp5_ASAP7_75t_L g8068 ( 
.A1(n_8037),
.A2(n_4322),
.B1(n_4340),
.B2(n_4281),
.Y(n_8068)
);

NOR4xp25_ASAP7_75t_L g8069 ( 
.A(n_8046),
.B(n_8015),
.C(n_8019),
.D(n_8035),
.Y(n_8069)
);

NAND3xp33_ASAP7_75t_SL g8070 ( 
.A(n_8061),
.B(n_8039),
.C(n_8042),
.Y(n_8070)
);

AND2x4_ASAP7_75t_SL g8071 ( 
.A(n_8049),
.B(n_8023),
.Y(n_8071)
);

AOI22xp5_ASAP7_75t_L g8072 ( 
.A1(n_8049),
.A2(n_8021),
.B1(n_8034),
.B2(n_8027),
.Y(n_8072)
);

HB1xp67_ASAP7_75t_L g8073 ( 
.A(n_8067),
.Y(n_8073)
);

NOR3x1_ASAP7_75t_L g8074 ( 
.A(n_8053),
.B(n_8030),
.C(n_3863),
.Y(n_8074)
);

INVx2_ASAP7_75t_L g8075 ( 
.A(n_8063),
.Y(n_8075)
);

OR2x6_ASAP7_75t_L g8076 ( 
.A(n_8056),
.B(n_3153),
.Y(n_8076)
);

NOR3x2_ASAP7_75t_L g8077 ( 
.A(n_8055),
.B(n_3649),
.C(n_3625),
.Y(n_8077)
);

AND4x1_ASAP7_75t_L g8078 ( 
.A(n_8047),
.B(n_4353),
.C(n_4327),
.D(n_4165),
.Y(n_8078)
);

AND3x4_ASAP7_75t_L g8079 ( 
.A(n_8060),
.B(n_3510),
.C(n_3556),
.Y(n_8079)
);

NAND3xp33_ASAP7_75t_SL g8080 ( 
.A(n_8052),
.B(n_4238),
.C(n_4013),
.Y(n_8080)
);

INVx1_ASAP7_75t_L g8081 ( 
.A(n_8065),
.Y(n_8081)
);

OR2x2_ASAP7_75t_L g8082 ( 
.A(n_8062),
.B(n_4845),
.Y(n_8082)
);

NAND2xp5_ASAP7_75t_L g8083 ( 
.A(n_8051),
.B(n_4845),
.Y(n_8083)
);

OR2x2_ASAP7_75t_L g8084 ( 
.A(n_8057),
.B(n_4845),
.Y(n_8084)
);

OR4x1_ASAP7_75t_L g8085 ( 
.A(n_8045),
.B(n_3742),
.C(n_3688),
.D(n_3724),
.Y(n_8085)
);

INVx1_ASAP7_75t_L g8086 ( 
.A(n_8066),
.Y(n_8086)
);

NOR2xp33_ASAP7_75t_L g8087 ( 
.A(n_8073),
.B(n_8064),
.Y(n_8087)
);

NAND2xp5_ASAP7_75t_L g8088 ( 
.A(n_8081),
.B(n_8071),
.Y(n_8088)
);

INVx2_ASAP7_75t_L g8089 ( 
.A(n_8075),
.Y(n_8089)
);

INVxp67_ASAP7_75t_L g8090 ( 
.A(n_8070),
.Y(n_8090)
);

NOR2xp33_ASAP7_75t_L g8091 ( 
.A(n_8086),
.B(n_8059),
.Y(n_8091)
);

OAI21xp33_ASAP7_75t_L g8092 ( 
.A1(n_8072),
.A2(n_8068),
.B(n_8058),
.Y(n_8092)
);

XNOR2xp5_ASAP7_75t_L g8093 ( 
.A(n_8069),
.B(n_8048),
.Y(n_8093)
);

NAND2xp5_ASAP7_75t_L g8094 ( 
.A(n_8082),
.B(n_8054),
.Y(n_8094)
);

AOI22xp5_ASAP7_75t_L g8095 ( 
.A1(n_8076),
.A2(n_8050),
.B1(n_3625),
.B2(n_4322),
.Y(n_8095)
);

NAND2xp33_ASAP7_75t_L g8096 ( 
.A(n_8083),
.B(n_3503),
.Y(n_8096)
);

INVx1_ASAP7_75t_L g8097 ( 
.A(n_8077),
.Y(n_8097)
);

INVx1_ASAP7_75t_L g8098 ( 
.A(n_8074),
.Y(n_8098)
);

OAI22xp5_ASAP7_75t_L g8099 ( 
.A1(n_8076),
.A2(n_8084),
.B1(n_8079),
.B2(n_8085),
.Y(n_8099)
);

NOR2xp67_ASAP7_75t_L g8100 ( 
.A(n_8080),
.B(n_3649),
.Y(n_8100)
);

INVx1_ASAP7_75t_L g8101 ( 
.A(n_8078),
.Y(n_8101)
);

XOR2xp5_ASAP7_75t_L g8102 ( 
.A(n_8088),
.B(n_3786),
.Y(n_8102)
);

INVx1_ASAP7_75t_L g8103 ( 
.A(n_8089),
.Y(n_8103)
);

INVx1_ASAP7_75t_L g8104 ( 
.A(n_8090),
.Y(n_8104)
);

INVx2_ASAP7_75t_L g8105 ( 
.A(n_8098),
.Y(n_8105)
);

INVx1_ASAP7_75t_L g8106 ( 
.A(n_8093),
.Y(n_8106)
);

XNOR2x1_ASAP7_75t_L g8107 ( 
.A(n_8097),
.B(n_4238),
.Y(n_8107)
);

AOI22xp5_ASAP7_75t_L g8108 ( 
.A1(n_8087),
.A2(n_3625),
.B1(n_4322),
.B2(n_4281),
.Y(n_8108)
);

OAI22xp5_ASAP7_75t_L g8109 ( 
.A1(n_8101),
.A2(n_3625),
.B1(n_4238),
.B2(n_4405),
.Y(n_8109)
);

INVx1_ASAP7_75t_L g8110 ( 
.A(n_8099),
.Y(n_8110)
);

INVx2_ASAP7_75t_L g8111 ( 
.A(n_8094),
.Y(n_8111)
);

XOR2xp5_ASAP7_75t_L g8112 ( 
.A(n_8091),
.B(n_3900),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_8096),
.Y(n_8113)
);

INVx1_ASAP7_75t_L g8114 ( 
.A(n_8092),
.Y(n_8114)
);

INVx1_ASAP7_75t_L g8115 ( 
.A(n_8100),
.Y(n_8115)
);

INVx2_ASAP7_75t_L g8116 ( 
.A(n_8104),
.Y(n_8116)
);

INVx1_ASAP7_75t_L g8117 ( 
.A(n_8103),
.Y(n_8117)
);

INVx1_ASAP7_75t_L g8118 ( 
.A(n_8111),
.Y(n_8118)
);

XOR2x1_ASAP7_75t_L g8119 ( 
.A(n_8115),
.B(n_8095),
.Y(n_8119)
);

AOI22xp5_ASAP7_75t_L g8120 ( 
.A1(n_8114),
.A2(n_4281),
.B1(n_4340),
.B2(n_4322),
.Y(n_8120)
);

INVxp67_ASAP7_75t_L g8121 ( 
.A(n_8106),
.Y(n_8121)
);

AOI22xp5_ASAP7_75t_L g8122 ( 
.A1(n_8110),
.A2(n_4281),
.B1(n_4340),
.B2(n_3514),
.Y(n_8122)
);

OAI21xp5_ASAP7_75t_L g8123 ( 
.A1(n_8105),
.A2(n_3602),
.B(n_4144),
.Y(n_8123)
);

AOI221xp5_ASAP7_75t_SL g8124 ( 
.A1(n_8113),
.A2(n_3815),
.B1(n_4391),
.B2(n_4394),
.C(n_4388),
.Y(n_8124)
);

INVxp67_ASAP7_75t_L g8125 ( 
.A(n_8102),
.Y(n_8125)
);

AOI22xp5_ASAP7_75t_L g8126 ( 
.A1(n_8107),
.A2(n_4340),
.B1(n_3088),
.B2(n_3090),
.Y(n_8126)
);

HB1xp67_ASAP7_75t_L g8127 ( 
.A(n_8118),
.Y(n_8127)
);

INVx1_ASAP7_75t_L g8128 ( 
.A(n_8116),
.Y(n_8128)
);

INVx1_ASAP7_75t_L g8129 ( 
.A(n_8121),
.Y(n_8129)
);

INVxp67_ASAP7_75t_SL g8130 ( 
.A(n_8117),
.Y(n_8130)
);

INVx1_ASAP7_75t_L g8131 ( 
.A(n_8119),
.Y(n_8131)
);

INVx1_ASAP7_75t_L g8132 ( 
.A(n_8125),
.Y(n_8132)
);

INVx1_ASAP7_75t_L g8133 ( 
.A(n_8126),
.Y(n_8133)
);

OA21x2_ASAP7_75t_L g8134 ( 
.A1(n_8130),
.A2(n_8108),
.B(n_8123),
.Y(n_8134)
);

INVx1_ASAP7_75t_L g8135 ( 
.A(n_8127),
.Y(n_8135)
);

OAI21x1_ASAP7_75t_L g8136 ( 
.A1(n_8128),
.A2(n_8112),
.B(n_8122),
.Y(n_8136)
);

INVx1_ASAP7_75t_L g8137 ( 
.A(n_8135),
.Y(n_8137)
);

INVx1_ASAP7_75t_L g8138 ( 
.A(n_8134),
.Y(n_8138)
);

AOI21xp5_ASAP7_75t_L g8139 ( 
.A1(n_8136),
.A2(n_8131),
.B(n_8129),
.Y(n_8139)
);

XNOR2xp5_ASAP7_75t_L g8140 ( 
.A(n_8139),
.B(n_8132),
.Y(n_8140)
);

AOI222xp33_ASAP7_75t_L g8141 ( 
.A1(n_8138),
.A2(n_8133),
.B1(n_8109),
.B2(n_8124),
.C1(n_8120),
.C2(n_3088),
.Y(n_8141)
);

OAI22xp5_ASAP7_75t_L g8142 ( 
.A1(n_8137),
.A2(n_3047),
.B1(n_4230),
.B2(n_3075),
.Y(n_8142)
);

OAI221xp5_ASAP7_75t_R g8143 ( 
.A1(n_8140),
.A2(n_3153),
.B1(n_3681),
.B2(n_4398),
.C(n_4397),
.Y(n_8143)
);

AOI22xp5_ASAP7_75t_L g8144 ( 
.A1(n_8143),
.A2(n_8141),
.B1(n_8142),
.B2(n_3088),
.Y(n_8144)
);

AOI21xp5_ASAP7_75t_L g8145 ( 
.A1(n_8144),
.A2(n_4133),
.B(n_3153),
.Y(n_8145)
);

AOI22x1_ASAP7_75t_L g8146 ( 
.A1(n_8145),
.A2(n_3075),
.B1(n_3142),
.B2(n_3063),
.Y(n_8146)
);

OAI221xp5_ASAP7_75t_R g8147 ( 
.A1(n_8146),
.A2(n_4404),
.B1(n_3153),
.B2(n_3882),
.C(n_3200),
.Y(n_8147)
);

AOI22xp5_ASAP7_75t_L g8148 ( 
.A1(n_8147),
.A2(n_3047),
.B1(n_3090),
.B2(n_3063),
.Y(n_8148)
);

AOI211xp5_ASAP7_75t_L g8149 ( 
.A1(n_8148),
.A2(n_3142),
.B(n_3181),
.C(n_3063),
.Y(n_8149)
);


endmodule