module fake_netlist_1_6020_n_32 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2xp33_ASAP7_75t_L g9 ( .A(n_3), .B(n_1), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_8), .B(n_3), .Y(n_10) );
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_4), .B(n_0), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
AND3x2_ASAP7_75t_L g13 ( .A(n_1), .B(n_5), .C(n_0), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_15), .Y(n_17) );
INVx8_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
AO21x2_ASAP7_75t_L g20 ( .A1(n_10), .A2(n_2), .B(n_11), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
INVxp67_ASAP7_75t_SL g22 ( .A(n_19), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_16), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_17), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
NAND4xp25_ASAP7_75t_L g26 ( .A(n_24), .B(n_9), .C(n_17), .D(n_13), .Y(n_26) );
AOI21xp5_ASAP7_75t_SL g27 ( .A1(n_24), .A2(n_21), .B(n_20), .Y(n_27) );
INVx2_ASAP7_75t_SL g28 ( .A(n_27), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_25), .B1(n_18), .B2(n_16), .Y(n_29) );
NAND4xp25_ASAP7_75t_L g30 ( .A(n_29), .B(n_25), .C(n_23), .D(n_18), .Y(n_30) );
OAI22xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_16), .B1(n_23), .B2(n_20), .Y(n_31) );
OAI21x1_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_16), .B(n_30), .Y(n_32) );
endmodule