module fake_jpeg_13753_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_24),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_37),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_50),
.Y(n_70)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_19),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_1),
.Y(n_74)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_55),
.B1(n_54),
.B2(n_52),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_81),
.B1(n_58),
.B2(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_78),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_49),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_57),
.B(n_53),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_54),
.B1(n_56),
.B2(n_43),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_40),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_71),
.B1(n_63),
.B2(n_59),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_85),
.B1(n_89),
.B2(n_7),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_69),
.B1(n_42),
.B2(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_73),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_71),
.B1(n_79),
.B2(n_68),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_47),
.B1(n_4),
.B2(n_7),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

BUFx24_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_94),
.C(n_12),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g93 ( 
.A(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_98),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_2),
.B(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_8),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_9),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_108),
.B(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_9),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_10),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_11),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_16),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_13),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_15),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_118),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_20),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_21),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_22),
.C(n_25),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_128),
.C(n_30),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_27),
.C(n_29),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_132),
.C(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_102),
.B(n_123),
.Y(n_134)
);

AOI21x1_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_136),
.B(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_138),
.B(n_106),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_106),
.B(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_112),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_125),
.B(n_120),
.Y(n_142)
);

AO21x1_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_137),
.B(n_127),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_143),
.Y(n_144)
);


endmodule