module fake_jpeg_20982_n_144 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_14),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_25),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_15),
.B1(n_16),
.B2(n_14),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_37),
.B1(n_12),
.B2(n_17),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_23),
.A2(n_15),
.B1(n_13),
.B2(n_16),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_43),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_21),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_41),
.B1(n_30),
.B2(n_10),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_33),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_22),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_47),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_66),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_10),
.B(n_46),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_10),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_82),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_56),
.C(n_59),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_42),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_50),
.B1(n_30),
.B2(n_38),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_71),
.B1(n_69),
.B2(n_68),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_50),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_10),
.B(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_42),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_31),
.B1(n_28),
.B2(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_86),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_76),
.C(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_93),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_84),
.B1(n_93),
.B2(n_18),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_114),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_13),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_112),
.B1(n_31),
.B2(n_28),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_120),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_99),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_105),
.C(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_122),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_98),
.C(n_18),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_18),
.C(n_6),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_117),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_112),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_126),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_117),
.A2(n_0),
.B(n_1),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_1),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_6),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_133),
.Y(n_136)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_5),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_129),
.B(n_7),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_8),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_137),
.A2(n_135),
.B(n_131),
.C(n_136),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_2),
.B(n_3),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_28),
.Y(n_144)
);


endmodule