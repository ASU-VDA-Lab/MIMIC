module fake_jpeg_28855_n_325 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_325);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx2_ASAP7_75t_SL g104 ( 
.A(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_45),
.Y(n_58)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_0),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_71),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_0),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_30),
.B(n_0),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_20),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_1),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_81),
.B1(n_22),
.B2(n_42),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_20),
.Y(n_78)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_17),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_29),
.B1(n_20),
.B2(n_37),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_88),
.A2(n_113),
.B1(n_58),
.B2(n_55),
.Y(n_123)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_SL g95 ( 
.A(n_56),
.Y(n_95)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_33),
.Y(n_135)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_117),
.B1(n_27),
.B2(n_26),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_60),
.A2(n_37),
.B1(n_22),
.B2(n_23),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_33),
.B1(n_24),
.B2(n_26),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_61),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_125),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_136),
.B1(n_151),
.B2(n_88),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_23),
.C(n_24),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_86),
.A2(n_62),
.B1(n_64),
.B2(n_49),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_127),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_57),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_75),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_130),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_95),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_129),
.B(n_131),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_65),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_35),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_72),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_138),
.A3(n_147),
.B1(n_99),
.B2(n_38),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_113),
.A2(n_74),
.B(n_78),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_140),
.B(n_149),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_150),
.B1(n_44),
.B2(n_38),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_27),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_58),
.B(n_78),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_51),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_148),
.B1(n_98),
.B2(n_84),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_35),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_83),
.B(n_28),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_34),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_67),
.B1(n_79),
.B2(n_59),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_166),
.B1(n_141),
.B2(n_134),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_167),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_135),
.B1(n_130),
.B2(n_136),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_164),
.B1(n_140),
.B2(n_116),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_54),
.B1(n_82),
.B2(n_87),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_82),
.B1(n_109),
.B2(n_89),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_127),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_119),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_178),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_130),
.B1(n_126),
.B2(n_109),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_180),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_99),
.B1(n_110),
.B2(n_116),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_186),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_138),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_167),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_126),
.B1(n_89),
.B2(n_124),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_131),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_153),
.B(n_168),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_159),
.C(n_154),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_198),
.C(n_175),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_192),
.B(n_141),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_162),
.B(n_159),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_159),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_177),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_204),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_158),
.C(n_164),
.Y(n_198)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_200),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_157),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_179),
.B1(n_183),
.B2(n_177),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_205),
.A2(n_210),
.B1(n_211),
.B2(n_217),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_191),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_206),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_194),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_199),
.B(n_187),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_183),
.B1(n_174),
.B2(n_178),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_178),
.B1(n_186),
.B2(n_181),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_190),
.B(n_203),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_189),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_195),
.A2(n_186),
.B1(n_182),
.B2(n_184),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_215),
.A2(n_219),
.B1(n_202),
.B2(n_204),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_172),
.B1(n_171),
.B2(n_158),
.Y(n_217)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_201),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_126),
.B1(n_171),
.B2(n_120),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_220),
.A2(n_225),
.B1(n_205),
.B2(n_210),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_226),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_224),
.C(n_228),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_198),
.C(n_190),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_202),
.B1(n_196),
.B2(n_201),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_203),
.C(n_169),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_169),
.C(n_149),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_139),
.B(n_148),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_216),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_219),
.B1(n_211),
.B2(n_212),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_153),
.B1(n_155),
.B2(n_124),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_241),
.B(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_244),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_234),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_250),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_165),
.B(n_208),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_217),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_247),
.C(n_223),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_165),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_137),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_161),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_249),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_220),
.A2(n_34),
.B1(n_44),
.B2(n_46),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_225),
.B(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_265),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_235),
.B(n_230),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_259),
.C(n_264),
.Y(n_274)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

INVx13_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_99),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_129),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_231),
.B1(n_171),
.B2(n_120),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_263),
.B1(n_245),
.B2(n_247),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_155),
.C(n_146),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_143),
.C(n_144),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_267),
.B(n_265),
.Y(n_281)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_276),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_246),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_277),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_235),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_260),
.A2(n_142),
.B1(n_110),
.B2(n_145),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_133),
.B1(n_115),
.B2(n_47),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_254),
.Y(n_285)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_257),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_286),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_122),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_251),
.B1(n_261),
.B2(n_266),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_290),
.B1(n_283),
.B2(n_289),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_264),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_291),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_273),
.C(n_259),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_255),
.C(n_266),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_292),
.A2(n_114),
.B(n_50),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_278),
.C(n_279),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_300),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_133),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_299),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_1),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_287),
.C(n_48),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_1),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_302),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_80),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_303),
.B(n_305),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_2),
.B(n_3),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_2),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_310),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_2),
.B(n_4),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_311),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_4),
.C(n_5),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_313),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_4),
.C(n_6),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_9),
.C(n_10),
.Y(n_316)
);

OAI31xp33_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_308),
.A3(n_304),
.B(n_12),
.Y(n_318)
);

AOI321xp33_ASAP7_75t_SL g322 ( 
.A1(n_318),
.A2(n_122),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.C(n_9),
.Y(n_322)
);

AOI21x1_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_314),
.B(n_308),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_321),
.A2(n_322),
.B(n_319),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_14),
.B(n_16),
.Y(n_324)
);

OAI311xp33_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_14),
.A3(n_80),
.B1(n_122),
.C1(n_322),
.Y(n_325)
);


endmodule