module fake_netlist_6_2396_n_1760 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1760);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1760;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_6),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_52),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_99),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_159),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_65),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_32),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_75),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_106),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_40),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_0),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_28),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_78),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_120),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_23),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_12),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_112),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_117),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_67),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_3),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_175),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_22),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_101),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_53),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_81),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_46),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_68),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_16),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_41),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_57),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_138),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_25),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_46),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_114),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_5),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_94),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_61),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_77),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_17),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_9),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_148),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_149),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_146),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_22),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_163),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_172),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_26),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_52),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_104),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_118),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_25),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_16),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_3),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_105),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_131),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_32),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_74),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_35),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_1),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_43),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_51),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_70),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_85),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_28),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_136),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_39),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_36),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_2),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_89),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_102),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_40),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_59),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_41),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_145),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_147),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_142),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_95),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_8),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_100),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_69),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_57),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_71),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_107),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_123),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_13),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_126),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_50),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_150),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_4),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_56),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_24),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_18),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_7),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_130),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_37),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_38),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_48),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_110),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_173),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_19),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_33),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_9),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_11),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_82),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_63),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_34),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_1),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_51),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_141),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_36),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_53),
.Y(n_298)
);

BUFx2_ASAP7_75t_SL g299 ( 
.A(n_113),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_93),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_35),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_124),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_168),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_116),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_155),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_14),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_72),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_8),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_21),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_33),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_29),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_54),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_11),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_47),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_171),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_24),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_26),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_44),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_161),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_19),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_87),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_88),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_103),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_56),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_154),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_14),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_121),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_12),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_49),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_37),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_132),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_153),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_6),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_83),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_45),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_50),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_137),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_48),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_49),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_10),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_91),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_96),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_31),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_30),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_119),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_79),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_162),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_15),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_31),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_23),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_0),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_140),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_160),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_191),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_219),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_199),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_219),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_210),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_213),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_196),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_196),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_177),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_298),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_196),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_276),
.B(n_2),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_263),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_196),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_276),
.B(n_4),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_296),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_331),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_196),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_177),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_196),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_196),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_196),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_305),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_320),
.B(n_7),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_251),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_320),
.B(n_10),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_251),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_251),
.Y(n_382)
);

INVxp33_ASAP7_75t_L g383 ( 
.A(n_179),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_352),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_251),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_211),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_212),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_316),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_316),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_216),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_214),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_223),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_224),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_231),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_232),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_219),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_239),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_241),
.B(n_15),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_348),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_348),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_251),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_283),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_240),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_220),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_185),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_272),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_238),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_283),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_283),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_283),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_180),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_221),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_243),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_339),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_188),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_262),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_225),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_185),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_190),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_192),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_193),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_201),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_245),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_246),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_247),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_209),
.B(n_217),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_184),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_226),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_229),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_262),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_235),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_248),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_258),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_277),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_282),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_253),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_262),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_287),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_215),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_197),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_186),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_289),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_230),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_393),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_359),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_368),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_406),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_361),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_354),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_373),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_359),
.B(n_267),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_414),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_420),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_407),
.B(n_257),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_421),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_431),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_432),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_379),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_R g464 ( 
.A(n_446),
.B(n_233),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_362),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_356),
.Y(n_466)
);

BUFx8_ASAP7_75t_L g467 ( 
.A(n_443),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_358),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_381),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_381),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_418),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_367),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_365),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_370),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_440),
.B(n_267),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_387),
.B(n_267),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_386),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_368),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_400),
.B(n_257),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_371),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_384),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_385),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_386),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_385),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_389),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_377),
.B(n_337),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_411),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_389),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_411),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_409),
.A2(n_324),
.B1(n_340),
.B2(n_350),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_360),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_360),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_372),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_392),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_392),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_412),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_412),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_372),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_403),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_R g502 ( 
.A(n_394),
.B(n_234),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_388),
.B(n_309),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_374),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_394),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_408),
.B(n_301),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_R g507 ( 
.A(n_395),
.B(n_244),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_404),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_419),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_364),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_395),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_374),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_419),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_364),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_396),
.B(n_337),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_413),
.B(n_178),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_375),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_375),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_376),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_430),
.B(n_215),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_396),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_376),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_481),
.B(n_250),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_481),
.B(n_521),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_444),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_523),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_523),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_480),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_508),
.B(n_397),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_521),
.B(n_250),
.Y(n_531)
);

AO22x2_ASAP7_75t_L g532 ( 
.A1(n_476),
.A2(n_295),
.B1(n_297),
.B2(n_228),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_479),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_480),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_493),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_501),
.Y(n_536)
);

CKINVDCx8_ASAP7_75t_R g537 ( 
.A(n_471),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_519),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_521),
.B(n_250),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_519),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_521),
.B(n_250),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_503),
.B(n_438),
.Y(n_542)
);

OR2x2_ASAP7_75t_SL g543 ( 
.A(n_471),
.B(n_429),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_519),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_480),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_493),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_495),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_519),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_506),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_449),
.B(n_250),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_453),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_458),
.B(n_399),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_495),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_494),
.B(n_443),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_516),
.B(n_405),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_495),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_500),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_449),
.B(n_405),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_449),
.B(n_415),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_494),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_449),
.B(n_415),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_511),
.B(n_355),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_488),
.B(n_426),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_513),
.B(n_426),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_486),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_517),
.B(n_275),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_486),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_503),
.A2(n_369),
.B1(n_366),
.B2(n_380),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_513),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_517),
.B(n_275),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_513),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_502),
.B(n_275),
.Y(n_572)
);

BUFx4f_ASAP7_75t_L g573 ( 
.A(n_486),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_513),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_486),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_486),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_455),
.B(n_427),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_500),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_485),
.B(n_427),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_509),
.B(n_438),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_L g581 ( 
.A1(n_492),
.A2(n_344),
.B1(n_288),
.B2(n_268),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_518),
.Y(n_582)
);

BUFx8_ASAP7_75t_SL g583 ( 
.A(n_466),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_452),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_511),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_500),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_504),
.B(n_428),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_504),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_504),
.B(n_428),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_520),
.B(n_435),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_464),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_468),
.Y(n_592)
);

OAI21xp33_ASAP7_75t_SL g593 ( 
.A1(n_478),
.A2(n_378),
.B(n_335),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_452),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_515),
.B(n_433),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_520),
.B(n_435),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_520),
.B(n_439),
.Y(n_597)
);

AND2x2_ASAP7_75t_SL g598 ( 
.A(n_522),
.B(n_275),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_515),
.A2(n_439),
.B1(n_433),
.B2(n_357),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_465),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_507),
.B(n_275),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_465),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_450),
.A2(n_398),
.B1(n_183),
.B2(n_182),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_465),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_474),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_478),
.B(n_317),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_474),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_461),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_461),
.B(n_442),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_463),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_463),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_469),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_509),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_450),
.B(n_390),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_454),
.A2(n_442),
.B1(n_336),
.B2(n_318),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_470),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_487),
.B(n_194),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_470),
.B(n_204),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_473),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_473),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_477),
.B(n_442),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_510),
.B(n_417),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_477),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_484),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_484),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_489),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_489),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_490),
.B(n_383),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_491),
.B(n_498),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_491),
.B(n_205),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_510),
.B(n_391),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_514),
.B(n_401),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_498),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_499),
.B(n_514),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_499),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_522),
.B(n_424),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_454),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_496),
.B(n_402),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_459),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_459),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_448),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_497),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_505),
.B(n_218),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_448),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_467),
.B(n_273),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_492),
.B(n_222),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_467),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_467),
.A2(n_299),
.B1(n_441),
.B2(n_437),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_467),
.B(n_281),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_512),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_447),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_451),
.B(n_423),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_456),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_457),
.B(n_429),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_460),
.B(n_434),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_462),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_472),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_475),
.B(n_256),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_482),
.B(n_227),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_483),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_611),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_598),
.A2(n_286),
.B1(n_261),
.B2(n_264),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_525),
.A2(n_436),
.B(n_445),
.C(n_425),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_525),
.B(n_527),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_611),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_528),
.B(n_626),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_631),
.Y(n_667)
);

BUFx12f_ASAP7_75t_L g668 ( 
.A(n_533),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_612),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_626),
.B(n_608),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_598),
.B(n_178),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_530),
.B(n_181),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_580),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_626),
.B(n_236),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_558),
.B(n_237),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_631),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_608),
.B(n_242),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_632),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_612),
.Y(n_679)
);

INVx8_ASAP7_75t_L g680 ( 
.A(n_654),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_552),
.B(n_183),
.Y(n_681)
);

A2O1A1Ixp33_ASAP7_75t_L g682 ( 
.A1(n_593),
.A2(n_252),
.B(n_300),
.C(n_292),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_628),
.B(n_187),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_632),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_536),
.B(n_559),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_561),
.B(n_249),
.Y(n_686)
);

NOR2xp67_ASAP7_75t_L g687 ( 
.A(n_591),
.B(n_266),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_564),
.B(n_259),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_600),
.B(n_285),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_577),
.A2(n_307),
.B1(n_269),
.B2(n_270),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_636),
.B(n_187),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_550),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_546),
.B(n_422),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_636),
.B(n_291),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_587),
.B(n_189),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_591),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_646),
.A2(n_342),
.B1(n_346),
.B2(n_353),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_622),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_622),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_636),
.B(n_189),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_555),
.B(n_195),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_589),
.B(n_195),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_563),
.A2(n_206),
.B1(n_202),
.B2(n_200),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_638),
.B(n_198),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_653),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_600),
.B(n_271),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_622),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_582),
.B(n_302),
.Y(n_708)
);

AND2x2_ASAP7_75t_SL g709 ( 
.A(n_648),
.B(n_422),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_590),
.A2(n_321),
.B1(n_303),
.B2(n_304),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_595),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_596),
.B(n_198),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_597),
.A2(n_322),
.B1(n_319),
.B2(n_315),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_594),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_613),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_524),
.A2(n_445),
.B(n_425),
.C(n_416),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_652),
.B(n_200),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_620),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_610),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_646),
.A2(n_197),
.B1(n_351),
.B2(n_349),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_526),
.B(n_202),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_610),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_614),
.B(n_206),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_610),
.B(n_208),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_623),
.B(n_208),
.Y(n_725)
);

AND2x2_ASAP7_75t_SL g726 ( 
.A(n_659),
.B(n_416),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_617),
.B(n_323),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_646),
.A2(n_327),
.B1(n_323),
.B2(n_347),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_542),
.B(n_325),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_623),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_580),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_624),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_623),
.B(n_325),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_616),
.B(n_327),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_542),
.B(n_332),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_624),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_646),
.A2(n_332),
.B1(n_334),
.B2(n_347),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_619),
.B(n_334),
.Y(n_738)
);

INVxp33_ASAP7_75t_L g739 ( 
.A(n_535),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_633),
.B(n_341),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_635),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_654),
.B(n_17),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_625),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_542),
.B(n_345),
.Y(n_744)
);

NOR2x1p5_ASAP7_75t_L g745 ( 
.A(n_647),
.B(n_203),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_546),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_615),
.B(n_306),
.C(n_254),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_524),
.B(n_345),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_560),
.B(n_255),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_560),
.B(n_260),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_L g751 ( 
.A(n_618),
.B(n_265),
.Y(n_751)
);

HB1xp67_ASAP7_75t_SL g752 ( 
.A(n_537),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_646),
.A2(n_351),
.B1(n_349),
.B2(n_343),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_554),
.B(n_203),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_585),
.B(n_274),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_617),
.B(n_278),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_581),
.B(n_310),
.C(n_279),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_580),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_585),
.B(n_599),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_569),
.B(n_280),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_531),
.A2(n_343),
.B(n_338),
.C(n_333),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_655),
.B(n_284),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_625),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_655),
.B(n_290),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_627),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_643),
.B(n_313),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_571),
.B(n_314),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_574),
.B(n_312),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_562),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_634),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_643),
.B(n_293),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_658),
.B(n_294),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_531),
.A2(n_338),
.B(n_333),
.C(n_330),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_642),
.B(n_308),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_642),
.B(n_647),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_629),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_637),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_644),
.B(n_90),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_529),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_573),
.A2(n_329),
.B(n_328),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_566),
.B(n_330),
.Y(n_781)
);

NOR3xp33_ASAP7_75t_L g782 ( 
.A(n_549),
.B(n_329),
.C(n_328),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_618),
.B(n_326),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_529),
.Y(n_784)
);

NOR2x1p5_ASAP7_75t_L g785 ( 
.A(n_647),
.B(n_326),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_583),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_562),
.B(n_637),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_534),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_644),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_566),
.A2(n_207),
.B(n_20),
.C(n_21),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_539),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_639),
.B(n_207),
.Y(n_792)
);

OAI221xp5_ASAP7_75t_L g793 ( 
.A1(n_568),
.A2(n_18),
.B1(n_20),
.B2(n_27),
.C(n_29),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_646),
.A2(n_86),
.B1(n_166),
.B2(n_165),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_639),
.B(n_27),
.Y(n_795)
);

INVx8_ASAP7_75t_L g796 ( 
.A(n_654),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_654),
.B(n_642),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_539),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_582),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_541),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_641),
.B(n_30),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_640),
.B(n_34),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_534),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_645),
.B(n_38),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_570),
.B(n_97),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_541),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_545),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_SL g808 ( 
.A(n_649),
.B(n_42),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_570),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_603),
.B(n_45),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_776),
.B(n_770),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_787),
.B(n_579),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_721),
.B(n_572),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_721),
.B(n_572),
.Y(n_814)
);

OAI321xp33_ASAP7_75t_L g815 ( 
.A1(n_793),
.A2(n_601),
.A3(n_651),
.B1(n_656),
.B2(n_532),
.C(n_657),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_681),
.A2(n_606),
.B1(n_532),
.B2(n_659),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_681),
.B(n_601),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_756),
.A2(n_606),
.B(n_630),
.C(n_607),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_672),
.A2(n_532),
.B1(n_618),
.B2(n_657),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_726),
.B(n_533),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_673),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_746),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_673),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_685),
.A2(n_548),
.B(n_575),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_666),
.A2(n_548),
.B(n_575),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_758),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_791),
.A2(n_800),
.B(n_798),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_731),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_706),
.A2(n_575),
.B(n_567),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_726),
.B(n_533),
.Y(n_830)
);

AO21x2_ASAP7_75t_L g831 ( 
.A1(n_708),
.A2(n_630),
.B(n_584),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_787),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_693),
.B(n_650),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_731),
.Y(n_834)
);

NOR3xp33_ASAP7_75t_L g835 ( 
.A(n_756),
.B(n_660),
.C(n_543),
.Y(n_835)
);

AOI21x1_ASAP7_75t_L g836 ( 
.A1(n_689),
.A2(n_588),
.B(n_557),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_695),
.B(n_544),
.Y(n_837)
);

NAND3xp33_ASAP7_75t_L g838 ( 
.A(n_727),
.B(n_650),
.C(n_660),
.Y(n_838)
);

NOR3xp33_ASAP7_75t_L g839 ( 
.A(n_766),
.B(n_621),
.C(n_609),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_766),
.A2(n_544),
.B(n_538),
.C(n_540),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_695),
.B(n_540),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_771),
.A2(n_544),
.B(n_538),
.C(n_540),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_806),
.A2(n_586),
.B(n_556),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_705),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_702),
.B(n_538),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_698),
.B(n_551),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_661),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_772),
.A2(n_618),
.B1(n_594),
.B2(n_602),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_789),
.B(n_537),
.Y(n_849)
);

BUFx12f_ASAP7_75t_L g850 ( 
.A(n_668),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_719),
.A2(n_545),
.B(n_557),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_697),
.A2(n_720),
.B1(n_753),
.B2(n_809),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_697),
.A2(n_588),
.B1(n_553),
.B2(n_556),
.Y(n_853)
);

NOR2x1p5_ASAP7_75t_SL g854 ( 
.A(n_779),
.B(n_578),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_702),
.B(n_578),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_686),
.A2(n_688),
.B(n_708),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_771),
.A2(n_605),
.B(n_604),
.C(n_547),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_739),
.B(n_592),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_665),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_724),
.A2(n_576),
.B(n_565),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_725),
.A2(n_586),
.B(n_553),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_733),
.A2(n_605),
.B(n_604),
.Y(n_862)
);

AOI21x1_ASAP7_75t_L g863 ( 
.A1(n_674),
.A2(n_618),
.B(n_550),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_711),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_769),
.B(n_592),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_705),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_741),
.B(n_550),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_720),
.A2(n_551),
.B1(n_54),
.B2(n_55),
.Y(n_868)
);

NOR2x1_ASAP7_75t_L g869 ( 
.A(n_687),
.B(n_583),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_805),
.A2(n_550),
.B(n_111),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_727),
.A2(n_550),
.B1(n_115),
.B2(n_122),
.Y(n_871)
);

OAI321xp33_ASAP7_75t_L g872 ( 
.A1(n_753),
.A2(n_47),
.A3(n_55),
.B1(n_58),
.B2(n_60),
.C(n_62),
.Y(n_872)
);

AOI21xp33_ASAP7_75t_L g873 ( 
.A1(n_701),
.A2(n_58),
.B(n_64),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_759),
.B(n_66),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_715),
.B(n_73),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_667),
.B(n_76),
.Y(n_876)
);

INVx11_ASAP7_75t_L g877 ( 
.A(n_752),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_809),
.A2(n_80),
.B1(n_84),
.B2(n_92),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_799),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_723),
.B(n_98),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_777),
.B(n_108),
.Y(n_881)
);

AO21x1_ASAP7_75t_L g882 ( 
.A1(n_671),
.A2(n_125),
.B(n_127),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_799),
.A2(n_133),
.B(n_135),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_676),
.B(n_139),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_722),
.A2(n_144),
.B(n_156),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_730),
.A2(n_157),
.B(n_158),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_669),
.A2(n_164),
.B(n_176),
.Y(n_887)
);

AOI22x1_ASAP7_75t_L g888 ( 
.A1(n_679),
.A2(n_736),
.B1(n_732),
.B2(n_743),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_678),
.B(n_684),
.Y(n_889)
);

AND2x2_ASAP7_75t_SL g890 ( 
.A(n_810),
.B(n_709),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_797),
.B(n_709),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_728),
.A2(n_737),
.B1(n_662),
.B2(n_790),
.Y(n_892)
);

BUFx8_ASAP7_75t_L g893 ( 
.A(n_801),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_795),
.A2(n_707),
.B1(n_699),
.B2(n_781),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_723),
.B(n_675),
.Y(n_895)
);

OAI22x1_ASAP7_75t_L g896 ( 
.A1(n_696),
.A2(n_786),
.B1(n_762),
.B2(n_764),
.Y(n_896)
);

AOI21x1_ASAP7_75t_L g897 ( 
.A1(n_763),
.A2(n_765),
.B(n_718),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_775),
.A2(n_712),
.B1(n_694),
.B2(n_677),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_710),
.B(n_713),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_680),
.Y(n_900)
);

BUFx8_ASAP7_75t_SL g901 ( 
.A(n_742),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_736),
.A2(n_784),
.B(n_807),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_680),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_760),
.A2(n_767),
.B(n_768),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_694),
.A2(n_748),
.B1(n_683),
.B2(n_704),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_680),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_795),
.A2(n_794),
.B1(n_802),
.B2(n_804),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_761),
.A2(n_773),
.B(n_792),
.C(n_663),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_788),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_803),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_716),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_734),
.A2(n_740),
.B(n_738),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_692),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_717),
.B(n_780),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_682),
.A2(n_783),
.B(n_751),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_690),
.B(n_703),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_802),
.B(n_729),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_691),
.A2(n_700),
.B(n_757),
.C(n_735),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_744),
.A2(n_755),
.B(n_750),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_749),
.A2(n_754),
.B(n_774),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_742),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_782),
.B(n_785),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_692),
.A2(n_808),
.B(n_747),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_692),
.A2(n_796),
.B(n_742),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_692),
.A2(n_796),
.B(n_745),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_796),
.A2(n_697),
.B1(n_753),
.B2(n_720),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_776),
.B(n_770),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_L g928 ( 
.A(n_727),
.B(n_766),
.C(n_756),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_739),
.B(n_408),
.Y(n_929)
);

OR2x6_ASAP7_75t_L g930 ( 
.A(n_680),
.B(n_796),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_776),
.A2(n_525),
.B1(n_770),
.B2(n_681),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_697),
.A2(n_753),
.B1(n_720),
.B2(n_809),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_776),
.B(n_770),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_776),
.B(n_770),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_673),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_776),
.B(n_770),
.Y(n_939)
);

NOR3xp33_ASAP7_75t_L g940 ( 
.A(n_756),
.B(n_628),
.C(n_577),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_673),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_L g942 ( 
.A(n_727),
.B(n_766),
.C(n_756),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_787),
.B(n_693),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_756),
.A2(n_771),
.B(n_766),
.C(n_727),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_776),
.B(n_770),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_776),
.B(n_770),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_697),
.A2(n_753),
.B1(n_720),
.B2(n_809),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_776),
.B(n_770),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_756),
.A2(n_771),
.B(n_766),
.C(n_727),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_758),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_714),
.A2(n_664),
.B(n_670),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_661),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_778),
.Y(n_960)
);

AOI33xp33_ASAP7_75t_L g961 ( 
.A1(n_720),
.A2(n_492),
.A3(n_581),
.B1(n_408),
.B2(n_753),
.B3(n_640),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_756),
.A2(n_771),
.B(n_766),
.C(n_727),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_726),
.B(n_598),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_776),
.B(n_770),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_664),
.A2(n_525),
.B(n_776),
.Y(n_965)
);

INVx5_ASAP7_75t_L g966 ( 
.A(n_692),
.Y(n_966)
);

NOR2xp67_ASAP7_75t_L g967 ( 
.A(n_696),
.B(n_650),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_673),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_946),
.A2(n_962),
.B(n_954),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_865),
.B(n_812),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_943),
.B(n_811),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_823),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_900),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_927),
.B(n_933),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_847),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_832),
.B(n_928),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_888),
.A2(n_902),
.B(n_836),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_826),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_861),
.A2(n_862),
.B(n_860),
.Y(n_979)
);

AOI21x1_ASAP7_75t_SL g980 ( 
.A1(n_916),
.A2(n_880),
.B(n_914),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_955),
.Y(n_981)
);

OAI22x1_ASAP7_75t_L g982 ( 
.A1(n_816),
.A2(n_942),
.B1(n_819),
.B2(n_921),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_890),
.B(n_849),
.Y(n_983)
);

BUFx12f_ASAP7_75t_L g984 ( 
.A(n_850),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_935),
.B(n_939),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_929),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_947),
.B(n_949),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_966),
.A2(n_936),
.B(n_934),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_940),
.A2(n_874),
.B(n_931),
.C(n_895),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_844),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_951),
.B(n_964),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_960),
.B(n_917),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_852),
.A2(n_950),
.B(n_932),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_960),
.B(n_817),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_822),
.Y(n_995)
);

AO31x2_ASAP7_75t_L g996 ( 
.A1(n_840),
.A2(n_842),
.A3(n_907),
.B(n_950),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_859),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_966),
.A2(n_944),
.B(n_937),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_900),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_900),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_966),
.A2(n_948),
.B(n_945),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_960),
.B(n_813),
.Y(n_1002)
);

AO21x1_ASAP7_75t_L g1003 ( 
.A1(n_907),
.A2(n_932),
.B(n_852),
.Y(n_1003)
);

AO21x1_ASAP7_75t_L g1004 ( 
.A1(n_814),
.A2(n_878),
.B(n_926),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_926),
.A2(n_891),
.B1(n_963),
.B2(n_878),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_966),
.A2(n_952),
.B(n_953),
.Y(n_1006)
);

CKINVDCx11_ASAP7_75t_R g1007 ( 
.A(n_846),
.Y(n_1007)
);

AOI21x1_ASAP7_75t_L g1008 ( 
.A1(n_837),
.A2(n_845),
.B(n_841),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_930),
.B(n_903),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_956),
.A2(n_958),
.B(n_957),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_829),
.A2(n_904),
.B(n_856),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_903),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_866),
.Y(n_1013)
);

AOI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_892),
.A2(n_815),
.B(n_899),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_825),
.A2(n_915),
.B(n_965),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_915),
.A2(n_965),
.B(n_824),
.Y(n_1016)
);

O2A1O1Ixp5_ASAP7_75t_L g1017 ( 
.A1(n_818),
.A2(n_912),
.B(n_894),
.C(n_908),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_820),
.B(n_830),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_851),
.A2(n_863),
.B(n_843),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_846),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_SL g1021 ( 
.A(n_868),
.B(n_967),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_833),
.B(n_905),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_855),
.A2(n_848),
.B(n_827),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_959),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_858),
.B(n_864),
.Y(n_1025)
);

INVx5_ASAP7_75t_L g1026 ( 
.A(n_930),
.Y(n_1026)
);

BUFx4f_ASAP7_75t_L g1027 ( 
.A(n_903),
.Y(n_1027)
);

BUFx12f_ASAP7_75t_L g1028 ( 
.A(n_893),
.Y(n_1028)
);

NAND2x1_ASAP7_75t_L g1029 ( 
.A(n_823),
.B(n_968),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_827),
.A2(n_913),
.B(n_968),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_889),
.B(n_918),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_961),
.A2(n_919),
.B(n_920),
.C(n_898),
.Y(n_1032)
);

AOI21x1_ASAP7_75t_L g1033 ( 
.A1(n_876),
.A2(n_884),
.B(n_875),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_892),
.A2(n_868),
.B1(n_894),
.B2(n_835),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_930),
.B(n_906),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_887),
.A2(n_821),
.B1(n_938),
.B2(n_941),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_SL g1037 ( 
.A1(n_881),
.A2(n_873),
.B(n_887),
.C(n_857),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_839),
.B(n_941),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_834),
.A2(n_919),
.B(n_867),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_909),
.B(n_828),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_879),
.B(n_911),
.Y(n_1041)
);

OA21x2_ASAP7_75t_L g1042 ( 
.A1(n_853),
.A2(n_920),
.B(n_882),
.Y(n_1042)
);

AO31x2_ASAP7_75t_L g1043 ( 
.A1(n_923),
.A2(n_870),
.A3(n_886),
.B(n_885),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_SL g1044 ( 
.A1(n_922),
.A2(n_872),
.B(n_854),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_871),
.A2(n_838),
.B(n_925),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_924),
.A2(n_883),
.B(n_869),
.C(n_906),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_831),
.A2(n_896),
.B(n_877),
.Y(n_1047)
);

OAI22x1_ASAP7_75t_L g1048 ( 
.A1(n_901),
.A2(n_816),
.B1(n_942),
.B2(n_928),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_943),
.B(n_811),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_943),
.B(n_946),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_897),
.A2(n_902),
.B(n_836),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_900),
.Y(n_1052)
);

AO31x2_ASAP7_75t_L g1053 ( 
.A1(n_946),
.A2(n_962),
.A3(n_954),
.B(n_842),
.Y(n_1053)
);

OAI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_946),
.A2(n_954),
.B(n_962),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_888),
.A2(n_902),
.B(n_836),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_844),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_966),
.A2(n_936),
.B(n_934),
.Y(n_1057)
);

INVx3_ASAP7_75t_SL g1058 ( 
.A(n_846),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_946),
.A2(n_962),
.B(n_954),
.Y(n_1059)
);

BUFx12f_ASAP7_75t_L g1060 ( 
.A(n_850),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_946),
.A2(n_962),
.B(n_954),
.C(n_942),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_812),
.B(n_832),
.Y(n_1062)
);

AO31x2_ASAP7_75t_L g1063 ( 
.A1(n_946),
.A2(n_962),
.A3(n_954),
.B(n_842),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_L g1064 ( 
.A1(n_897),
.A2(n_902),
.B(n_836),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_943),
.B(n_811),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_910),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_L g1067 ( 
.A(n_946),
.B(n_954),
.Y(n_1067)
);

BUFx4f_ASAP7_75t_L g1068 ( 
.A(n_900),
.Y(n_1068)
);

AO31x2_ASAP7_75t_L g1069 ( 
.A1(n_946),
.A2(n_962),
.A3(n_954),
.B(n_842),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_823),
.Y(n_1070)
);

INVx3_ASAP7_75t_SL g1071 ( 
.A(n_846),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_823),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_966),
.A2(n_936),
.B(n_934),
.Y(n_1073)
);

OA21x2_ASAP7_75t_L g1074 ( 
.A1(n_840),
.A2(n_842),
.B(n_851),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_946),
.A2(n_962),
.B(n_954),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_844),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_946),
.A2(n_962),
.B(n_954),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_930),
.B(n_680),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_844),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_910),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_865),
.B(n_549),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_966),
.A2(n_936),
.B(n_934),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_844),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_946),
.A2(n_962),
.A3(n_954),
.B(n_842),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_943),
.B(n_811),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_844),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_823),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_910),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_943),
.B(n_946),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_812),
.B(n_943),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_966),
.A2(n_936),
.B(n_934),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_900),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_943),
.B(n_811),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_900),
.Y(n_1094)
);

AO21x1_ASAP7_75t_L g1095 ( 
.A1(n_907),
.A2(n_932),
.B(n_852),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_SL g1096 ( 
.A1(n_928),
.A2(n_942),
.B(n_946),
.Y(n_1096)
);

AO31x2_ASAP7_75t_L g1097 ( 
.A1(n_946),
.A2(n_962),
.A3(n_954),
.B(n_842),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_966),
.A2(n_936),
.B(n_934),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_946),
.A2(n_962),
.B(n_954),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_865),
.B(n_549),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_984),
.Y(n_1101)
);

BUFx2_ASAP7_75t_R g1102 ( 
.A(n_1058),
.Y(n_1102)
);

OAI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_985),
.A2(n_987),
.B(n_974),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_970),
.B(n_1081),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_1026),
.B(n_1009),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1010),
.A2(n_1011),
.B(n_1067),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_988),
.A2(n_1001),
.B(n_998),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_978),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_1100),
.B(n_1090),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_995),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_985),
.A2(n_987),
.B1(n_991),
.B2(n_1005),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_1026),
.B(n_1027),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_971),
.B(n_1049),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_981),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_975),
.Y(n_1115)
);

INVx5_ASAP7_75t_L g1116 ( 
.A(n_973),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_1056),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_986),
.B(n_1062),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1026),
.B(n_1009),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_1079),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_SL g1121 ( 
.A1(n_1021),
.A2(n_983),
.B1(n_1099),
.B2(n_969),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_L g1122 ( 
.A1(n_969),
.A2(n_1099),
.B(n_1077),
.C(n_1075),
.Y(n_1122)
);

AND2x2_ASAP7_75t_SL g1123 ( 
.A(n_1021),
.B(n_1034),
.Y(n_1123)
);

AO21x2_ASAP7_75t_L g1124 ( 
.A1(n_1059),
.A2(n_1077),
.B(n_1075),
.Y(n_1124)
);

OR2x6_ASAP7_75t_L g1125 ( 
.A(n_1078),
.B(n_1035),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1034),
.A2(n_1054),
.B1(n_1003),
.B2(n_1095),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1006),
.A2(n_1098),
.B(n_1057),
.Y(n_1127)
);

INVx4_ASAP7_75t_SL g1128 ( 
.A(n_1071),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_976),
.B(n_1065),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1073),
.A2(n_1091),
.B(n_1082),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1027),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_SL g1132 ( 
.A1(n_1047),
.A2(n_1031),
.B(n_1038),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_997),
.Y(n_1133)
);

AO21x2_ASAP7_75t_L g1134 ( 
.A1(n_1059),
.A2(n_1015),
.B(n_1016),
.Y(n_1134)
);

O2A1O1Ixp5_ASAP7_75t_SL g1135 ( 
.A1(n_1014),
.A2(n_993),
.B(n_1045),
.C(n_1038),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1085),
.B(n_1093),
.Y(n_1136)
);

INVx4_ASAP7_75t_L g1137 ( 
.A(n_1068),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_1007),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1083),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_1061),
.A2(n_1004),
.A3(n_1032),
.B(n_982),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1035),
.B(n_1078),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_1086),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_1060),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1054),
.A2(n_1096),
.B1(n_1005),
.B2(n_993),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1024),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_992),
.B(n_989),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1066),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1078),
.B(n_1012),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1041),
.Y(n_1149)
);

AOI222xp33_ASAP7_75t_L g1150 ( 
.A1(n_1048),
.A2(n_1096),
.B1(n_1020),
.B2(n_1089),
.C1(n_1050),
.C2(n_1025),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1079),
.B(n_1013),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1022),
.B(n_1018),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1068),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1080),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_994),
.B(n_1002),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1088),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1050),
.B(n_1089),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1040),
.Y(n_1158)
);

INVx3_ASAP7_75t_SL g1159 ( 
.A(n_973),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1014),
.A2(n_1042),
.B1(n_1036),
.B2(n_1039),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1023),
.B(n_1084),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_973),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1053),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_999),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_L g1165 ( 
.A(n_1052),
.B(n_1046),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1052),
.B(n_1000),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1037),
.A2(n_1017),
.B(n_1030),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_999),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_999),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1000),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1053),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1042),
.A2(n_1094),
.B1(n_1092),
.B2(n_1000),
.Y(n_1172)
);

INVx3_ASAP7_75t_SL g1173 ( 
.A(n_1092),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1063),
.B(n_1084),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1092),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_972),
.Y(n_1176)
);

NOR2x1_ASAP7_75t_SL g1177 ( 
.A(n_1033),
.B(n_1094),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1094),
.Y(n_1178)
);

NAND2x1p5_ASAP7_75t_L g1179 ( 
.A(n_1070),
.B(n_1072),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1063),
.B(n_1097),
.Y(n_1180)
);

BUFx4_ASAP7_75t_SL g1181 ( 
.A(n_1028),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1072),
.B(n_1087),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1063),
.B(n_1097),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1069),
.B(n_1084),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_996),
.B(n_1008),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1029),
.Y(n_1186)
);

NOR2xp67_ASAP7_75t_L g1187 ( 
.A(n_1051),
.B(n_1064),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1043),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1074),
.A2(n_1044),
.B1(n_980),
.B2(n_1019),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1074),
.B(n_1043),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_979),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1043),
.B(n_986),
.Y(n_1192)
);

NOR2x1_ASAP7_75t_SL g1193 ( 
.A(n_1078),
.B(n_960),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_985),
.B(n_987),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_978),
.Y(n_1195)
);

CKINVDCx16_ASAP7_75t_R g1196 ( 
.A(n_1076),
.Y(n_1196)
);

INVx3_ASAP7_75t_SL g1197 ( 
.A(n_1076),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_986),
.B(n_642),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_989),
.A2(n_946),
.B(n_962),
.C(n_954),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1026),
.B(n_1009),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_978),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_985),
.B(n_987),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1034),
.A2(n_928),
.B1(n_942),
.B2(n_940),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_970),
.B(n_1081),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1061),
.A2(n_954),
.B(n_946),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_985),
.B(n_987),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_984),
.Y(n_1207)
);

OA21x2_ASAP7_75t_L g1208 ( 
.A1(n_1017),
.A2(n_1055),
.B(n_977),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1010),
.A2(n_1011),
.B(n_1067),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_972),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_978),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_970),
.B(n_1081),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1090),
.B(n_983),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_SL g1214 ( 
.A1(n_969),
.A2(n_1059),
.B(n_1077),
.C(n_1075),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1026),
.B(n_1009),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1090),
.B(n_983),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_986),
.B(n_812),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_975),
.Y(n_1218)
);

INVx4_ASAP7_75t_L g1219 ( 
.A(n_1027),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_990),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1003),
.A2(n_928),
.B1(n_942),
.B2(n_940),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_1076),
.Y(n_1222)
);

OAI21xp33_ASAP7_75t_L g1223 ( 
.A1(n_985),
.A2(n_954),
.B(n_946),
.Y(n_1223)
);

O2A1O1Ixp5_ASAP7_75t_L g1224 ( 
.A1(n_969),
.A2(n_954),
.B(n_962),
.C(n_946),
.Y(n_1224)
);

AO21x1_ASAP7_75t_L g1225 ( 
.A1(n_1014),
.A2(n_1067),
.B(n_1059),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1026),
.B(n_1009),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_972),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1026),
.B(n_1009),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_SL g1229 ( 
.A1(n_969),
.A2(n_1059),
.B(n_1077),
.C(n_1075),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_970),
.B(n_1081),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1010),
.A2(n_1011),
.B(n_1067),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1026),
.B(n_1009),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_985),
.A2(n_932),
.B1(n_950),
.B2(n_852),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1108),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1120),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_1104),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1114),
.Y(n_1237)
);

BUFx2_ASAP7_75t_SL g1238 ( 
.A(n_1116),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1131),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1171),
.Y(n_1240)
);

NAND2x1p5_ASAP7_75t_L g1241 ( 
.A(n_1165),
.B(n_1123),
.Y(n_1241)
);

AO21x2_ASAP7_75t_L g1242 ( 
.A1(n_1107),
.A2(n_1130),
.B(n_1127),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1129),
.A2(n_1136),
.B1(n_1233),
.B2(n_1124),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1199),
.A2(n_1233),
.B(n_1167),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1151),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1116),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1113),
.B(n_1194),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1203),
.A2(n_1150),
.B1(n_1121),
.B2(n_1221),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1155),
.B(n_1203),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1140),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1110),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1150),
.A2(n_1144),
.B1(n_1124),
.B2(n_1223),
.Y(n_1252)
);

BUFx10_ASAP7_75t_L g1253 ( 
.A(n_1131),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1144),
.A2(n_1223),
.B1(n_1152),
.B2(n_1225),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1210),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1195),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1217),
.A2(n_1113),
.B1(n_1118),
.B2(n_1216),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1174),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1116),
.Y(n_1259)
);

BUFx10_ASAP7_75t_L g1260 ( 
.A(n_1131),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1194),
.B(n_1202),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1213),
.A2(n_1111),
.B1(n_1103),
.B2(n_1198),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1139),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1183),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1184),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1143),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1184),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1180),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1161),
.Y(n_1269)
);

INVx4_ASAP7_75t_SL g1270 ( 
.A(n_1140),
.Y(n_1270)
);

INVx5_ASAP7_75t_SL g1271 ( 
.A(n_1125),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1188),
.B(n_1192),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1103),
.A2(n_1111),
.B1(n_1126),
.B2(n_1146),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1126),
.A2(n_1230),
.B1(n_1204),
.B2(n_1212),
.Y(n_1274)
);

INVxp33_ASAP7_75t_L g1275 ( 
.A(n_1109),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1218),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1201),
.Y(n_1277)
);

AO21x1_ASAP7_75t_SL g1278 ( 
.A1(n_1185),
.A2(n_1160),
.B(n_1190),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1202),
.B(n_1206),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1211),
.Y(n_1280)
);

BUFx8_ASAP7_75t_L g1281 ( 
.A(n_1153),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1159),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1206),
.B(n_1149),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1141),
.B(n_1193),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1140),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1117),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1157),
.A2(n_1125),
.B1(n_1196),
.B2(n_1197),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1106),
.A2(n_1209),
.B(n_1231),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1141),
.A2(n_1134),
.B1(n_1132),
.B2(n_1138),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1133),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1157),
.B(n_1158),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1227),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1222),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1142),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1214),
.B(n_1229),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1227),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1145),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1147),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1154),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1105),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1178),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1156),
.Y(n_1302)
);

AOI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1189),
.A2(n_1185),
.B(n_1187),
.Y(n_1303)
);

BUFx4f_ASAP7_75t_SL g1304 ( 
.A(n_1173),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1105),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1119),
.A2(n_1200),
.B1(n_1232),
.B2(n_1215),
.Y(n_1306)
);

CKINVDCx6p67_ASAP7_75t_R g1307 ( 
.A(n_1137),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1179),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1208),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1205),
.A2(n_1112),
.B1(n_1219),
.B2(n_1137),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1224),
.B(n_1122),
.Y(n_1311)
);

BUFx12f_ASAP7_75t_L g1312 ( 
.A(n_1101),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1119),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1169),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1102),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1189),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1181),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1135),
.B(n_1176),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1182),
.Y(n_1319)
);

AOI222xp33_ASAP7_75t_L g1320 ( 
.A1(n_1128),
.A2(n_1200),
.B1(n_1228),
.B2(n_1215),
.C1(n_1226),
.C2(n_1220),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1182),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1177),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1191),
.B(n_1186),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1112),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1226),
.A2(n_1228),
.B1(n_1148),
.B2(n_1219),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1128),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1170),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1172),
.B(n_1148),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1169),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1169),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1166),
.A2(n_1162),
.B(n_1175),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1164),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1207),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1164),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1168),
.A2(n_1123),
.B1(n_942),
.B2(n_928),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1168),
.A2(n_940),
.B(n_506),
.Y(n_1336)
);

BUFx5_ASAP7_75t_L g1337 ( 
.A(n_1163),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1123),
.A2(n_942),
.B1(n_928),
.B2(n_940),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1120),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1115),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1108),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1108),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1116),
.Y(n_1343)
);

BUFx8_ASAP7_75t_L g1344 ( 
.A(n_1131),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1210),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1108),
.Y(n_1346)
);

BUFx4f_ASAP7_75t_SL g1347 ( 
.A(n_1222),
.Y(n_1347)
);

AOI222xp33_ASAP7_75t_L g1348 ( 
.A1(n_1123),
.A2(n_868),
.B1(n_646),
.B2(n_950),
.C1(n_932),
.C2(n_852),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1108),
.Y(n_1349)
);

BUFx2_ASAP7_75t_R g1350 ( 
.A(n_1101),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1123),
.A2(n_942),
.B1(n_928),
.B2(n_940),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1115),
.Y(n_1352)
);

AO21x2_ASAP7_75t_L g1353 ( 
.A1(n_1107),
.A2(n_1059),
.B(n_969),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1108),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1323),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1343),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1240),
.Y(n_1357)
);

BUFx2_ASAP7_75t_SL g1358 ( 
.A(n_1343),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1288),
.A2(n_1303),
.B(n_1316),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1288),
.A2(n_1316),
.B(n_1309),
.Y(n_1360)
);

INVxp67_ASAP7_75t_SL g1361 ( 
.A(n_1339),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1249),
.B(n_1261),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1235),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1328),
.B(n_1284),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1249),
.B(n_1261),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1240),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1337),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1337),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1328),
.B(n_1284),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1311),
.B(n_1250),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1337),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1337),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1338),
.A2(n_1351),
.B(n_1243),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1235),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1245),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1269),
.B(n_1268),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1311),
.B(n_1250),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1331),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1331),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1285),
.B(n_1318),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1258),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1284),
.B(n_1270),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1343),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1270),
.B(n_1322),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1295),
.B(n_1285),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1318),
.B(n_1283),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1248),
.A2(n_1348),
.B1(n_1252),
.B2(n_1335),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1273),
.A2(n_1254),
.B(n_1336),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1272),
.B(n_1244),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1295),
.B(n_1264),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1347),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1236),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1283),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1280),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1242),
.A2(n_1353),
.B(n_1262),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1265),
.B(n_1267),
.Y(n_1396)
);

AO21x2_ASAP7_75t_L g1397 ( 
.A1(n_1353),
.A2(n_1265),
.B(n_1267),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1247),
.B(n_1279),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1287),
.A2(n_1354),
.B(n_1234),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1293),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1272),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1308),
.B(n_1319),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1257),
.B(n_1291),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1241),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1274),
.B(n_1275),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1271),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1278),
.B(n_1241),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1301),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1237),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1256),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1277),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1294),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1341),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1342),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1294),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1346),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1278),
.B(n_1241),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1349),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1297),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1319),
.B(n_1321),
.Y(n_1420)
);

BUFx4f_ASAP7_75t_SL g1421 ( 
.A(n_1312),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1310),
.A2(n_1289),
.B(n_1290),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1386),
.B(n_1275),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1370),
.B(n_1352),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1382),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1385),
.B(n_1271),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1385),
.B(n_1340),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1370),
.B(n_1377),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1377),
.B(n_1340),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_SL g1430 ( 
.A(n_1389),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1378),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1380),
.B(n_1276),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1395),
.B(n_1298),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1397),
.B(n_1302),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1379),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1397),
.B(n_1299),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1382),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1355),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1395),
.B(n_1251),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1395),
.B(n_1292),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1390),
.B(n_1330),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1387),
.A2(n_1320),
.B1(n_1325),
.B2(n_1306),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1363),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1357),
.Y(n_1444)
);

OAI33xp33_ASAP7_75t_L g1445 ( 
.A1(n_1375),
.A2(n_1403),
.A3(n_1398),
.B1(n_1390),
.B2(n_1405),
.B3(n_1409),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1389),
.B(n_1360),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1384),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1389),
.B(n_1255),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1389),
.B(n_1296),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1389),
.B(n_1296),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1357),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1399),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1359),
.B(n_1345),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1366),
.B(n_1329),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1428),
.B(n_1364),
.Y(n_1455)
);

NOR3xp33_ASAP7_75t_L g1456 ( 
.A(n_1445),
.B(n_1388),
.C(n_1373),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1428),
.B(n_1364),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1423),
.B(n_1361),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1442),
.A2(n_1404),
.B1(n_1400),
.B2(n_1407),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1452),
.B(n_1392),
.C(n_1422),
.Y(n_1460)
);

AOI21xp33_ASAP7_75t_L g1461 ( 
.A1(n_1439),
.A2(n_1399),
.B(n_1404),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1423),
.B(n_1374),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1443),
.B(n_1391),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1443),
.B(n_1393),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1424),
.B(n_1429),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1424),
.B(n_1362),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1442),
.A2(n_1407),
.B1(n_1417),
.B2(n_1415),
.Y(n_1467)
);

OAI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1452),
.A2(n_1333),
.B1(n_1326),
.B2(n_1315),
.C(n_1412),
.Y(n_1468)
);

AOI21xp33_ASAP7_75t_L g1469 ( 
.A1(n_1439),
.A2(n_1399),
.B(n_1417),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_SL g1470 ( 
.A(n_1445),
.B(n_1350),
.Y(n_1470)
);

OAI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1439),
.A2(n_1362),
.B(n_1365),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1430),
.A2(n_1369),
.B1(n_1401),
.B2(n_1420),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1424),
.B(n_1365),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1433),
.B(n_1408),
.C(n_1414),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1432),
.B(n_1369),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1429),
.B(n_1394),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1448),
.B(n_1367),
.Y(n_1477)
);

NAND2xp33_ASAP7_75t_SL g1478 ( 
.A(n_1430),
.B(n_1317),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1430),
.A2(n_1401),
.B1(n_1420),
.B2(n_1402),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1448),
.B(n_1368),
.Y(n_1480)
);

OAI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1426),
.A2(n_1313),
.B1(n_1305),
.B2(n_1263),
.C(n_1324),
.Y(n_1481)
);

AOI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1430),
.A2(n_1419),
.B1(n_1409),
.B2(n_1410),
.C(n_1411),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1449),
.B(n_1368),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1447),
.A2(n_1383),
.B(n_1356),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1441),
.B(n_1416),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1426),
.A2(n_1402),
.B1(n_1420),
.B2(n_1421),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1441),
.A2(n_1396),
.B1(n_1376),
.B2(n_1381),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1444),
.B(n_1418),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1426),
.A2(n_1420),
.B1(n_1402),
.B2(n_1406),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1449),
.B(n_1371),
.Y(n_1490)
);

AND2x2_ASAP7_75t_SL g1491 ( 
.A(n_1446),
.B(n_1355),
.Y(n_1491)
);

OAI221xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1446),
.A2(n_1433),
.B1(n_1440),
.B2(n_1307),
.C(n_1427),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_L g1493 ( 
.A(n_1433),
.B(n_1410),
.C(n_1411),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1434),
.B(n_1413),
.C(n_1414),
.Y(n_1494)
);

OA211x2_ASAP7_75t_L g1495 ( 
.A1(n_1447),
.A2(n_1358),
.B(n_1383),
.C(n_1356),
.Y(n_1495)
);

OAI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1438),
.A2(n_1305),
.B1(n_1313),
.B2(n_1263),
.C(n_1282),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1444),
.B(n_1418),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1450),
.B(n_1372),
.Y(n_1498)
);

NAND3xp33_ASAP7_75t_L g1499 ( 
.A(n_1434),
.B(n_1419),
.C(n_1413),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1450),
.B(n_1372),
.Y(n_1500)
);

OAI221xp5_ASAP7_75t_L g1501 ( 
.A1(n_1438),
.A2(n_1282),
.B1(n_1286),
.B2(n_1239),
.C(n_1300),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1450),
.B(n_1440),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1502),
.B(n_1446),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1502),
.B(n_1425),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1491),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1477),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1488),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1491),
.B(n_1440),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1468),
.B(n_1454),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1477),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1480),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1497),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1491),
.B(n_1453),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1480),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1455),
.B(n_1453),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1457),
.B(n_1453),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1494),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1460),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1493),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1494),
.B(n_1451),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1456),
.B(n_1454),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1483),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1493),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1499),
.Y(n_1524)
);

NAND2x1p5_ASAP7_75t_SL g1525 ( 
.A(n_1470),
.B(n_1438),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1485),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1499),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1471),
.B(n_1436),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1476),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1471),
.B(n_1436),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1474),
.B(n_1431),
.Y(n_1531)
);

AND2x2_ASAP7_75t_SL g1532 ( 
.A(n_1470),
.B(n_1482),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1487),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1464),
.B(n_1451),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1474),
.B(n_1431),
.Y(n_1535)
);

NOR2x1_ASAP7_75t_L g1536 ( 
.A(n_1521),
.B(n_1460),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1532),
.A2(n_1467),
.B1(n_1459),
.B2(n_1486),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1521),
.B(n_1466),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1527),
.B(n_1465),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1520),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1511),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1518),
.B(n_1509),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1527),
.B(n_1473),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1520),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1513),
.B(n_1490),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1520),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1534),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1533),
.B(n_1519),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1517),
.Y(n_1549)
);

INVx3_ASAP7_75t_SL g1550 ( 
.A(n_1532),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1509),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1517),
.Y(n_1552)
);

NOR3xp33_ASAP7_75t_L g1553 ( 
.A(n_1518),
.B(n_1501),
.C(n_1496),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1529),
.B(n_1462),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1505),
.B(n_1425),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1513),
.B(n_1490),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1511),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_L g1558 ( 
.A(n_1519),
.B(n_1484),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1534),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1511),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1533),
.B(n_1458),
.Y(n_1561)
);

INVx3_ASAP7_75t_R g1562 ( 
.A(n_1534),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1529),
.B(n_1475),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1523),
.B(n_1492),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1524),
.Y(n_1565)
);

NOR2x1p5_ASAP7_75t_L g1566 ( 
.A(n_1505),
.B(n_1528),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1513),
.B(n_1498),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1524),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1503),
.B(n_1508),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1505),
.B(n_1437),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1523),
.B(n_1435),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1503),
.B(n_1498),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1526),
.B(n_1500),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1535),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1503),
.B(n_1500),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1562),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1547),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1551),
.B(n_1515),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1548),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1542),
.B(n_1266),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1550),
.A2(n_1532),
.B1(n_1505),
.B2(n_1525),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1540),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1569),
.B(n_1505),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1555),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1540),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_SL g1586 ( 
.A(n_1550),
.B(n_1532),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1569),
.B(n_1566),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1548),
.B(n_1528),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1555),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1546),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1537),
.A2(n_1472),
.B1(n_1479),
.B2(n_1530),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1559),
.B(n_1530),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1545),
.B(n_1504),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1546),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1541),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1545),
.B(n_1504),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1556),
.B(n_1504),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1541),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1561),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1561),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1536),
.A2(n_1478),
.B1(n_1469),
.B2(n_1481),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1553),
.B(n_1515),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1549),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1538),
.B(n_1515),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1549),
.B(n_1535),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1564),
.B(n_1543),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1571),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1557),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1564),
.A2(n_1506),
.B1(n_1510),
.B2(n_1514),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1552),
.B(n_1461),
.C(n_1531),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1571),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1555),
.Y(n_1612)
);

INVxp67_ASAP7_75t_SL g1613 ( 
.A(n_1558),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1556),
.B(n_1504),
.Y(n_1614)
);

AOI21xp33_ASAP7_75t_L g1615 ( 
.A1(n_1552),
.A2(n_1531),
.B(n_1535),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1565),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1565),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1554),
.B(n_1266),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1543),
.B(n_1516),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1576),
.B(n_1570),
.Y(n_1620)
);

CKINVDCx16_ASAP7_75t_R g1621 ( 
.A(n_1586),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1581),
.A2(n_1568),
.B1(n_1574),
.B2(n_1544),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1606),
.B(n_1568),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1595),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1582),
.Y(n_1625)
);

INVxp33_ASAP7_75t_L g1626 ( 
.A(n_1580),
.Y(n_1626)
);

NOR2x1p5_ASAP7_75t_L g1627 ( 
.A(n_1613),
.B(n_1317),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1584),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1582),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1587),
.B(n_1570),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1595),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1601),
.A2(n_1525),
.B1(n_1562),
.B2(n_1539),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1587),
.B(n_1570),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1579),
.B(n_1539),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1598),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1602),
.A2(n_1591),
.B1(n_1610),
.B2(n_1600),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1618),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1585),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1593),
.B(n_1567),
.Y(n_1639)
);

NOR2x1_ASAP7_75t_L g1640 ( 
.A(n_1603),
.B(n_1616),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1584),
.B(n_1567),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1593),
.B(n_1572),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1596),
.B(n_1572),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1598),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1608),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1578),
.B(n_1312),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1605),
.B(n_1557),
.Y(n_1647)
);

CKINVDCx16_ASAP7_75t_R g1648 ( 
.A(n_1609),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1605),
.B(n_1560),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1608),
.A2(n_1560),
.B(n_1522),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1596),
.B(n_1575),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1589),
.B(n_1575),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1599),
.B(n_1516),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1585),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1590),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_L g1656 ( 
.A(n_1622),
.B(n_1615),
.C(n_1617),
.Y(n_1656)
);

AOI222xp33_ASAP7_75t_L g1657 ( 
.A1(n_1636),
.A2(n_1611),
.B1(n_1607),
.B2(n_1577),
.C1(n_1583),
.C2(n_1590),
.Y(n_1657)
);

INVxp67_ASAP7_75t_SL g1658 ( 
.A(n_1627),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1625),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1625),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1629),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1636),
.A2(n_1607),
.B1(n_1611),
.B2(n_1594),
.C(n_1577),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1629),
.Y(n_1663)
);

AOI31xp33_ASAP7_75t_L g1664 ( 
.A1(n_1626),
.A2(n_1589),
.A3(n_1612),
.B(n_1592),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1648),
.A2(n_1594),
.B(n_1588),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1623),
.B(n_1604),
.Y(n_1666)
);

AOI211xp5_ASAP7_75t_L g1667 ( 
.A1(n_1622),
.A2(n_1632),
.B(n_1623),
.C(n_1648),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1620),
.B(n_1597),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1637),
.B(n_1583),
.Y(n_1669)
);

AOI211x1_ASAP7_75t_L g1670 ( 
.A1(n_1632),
.A2(n_1619),
.B(n_1614),
.C(n_1597),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1620),
.Y(n_1671)
);

AOI21xp33_ASAP7_75t_SL g1672 ( 
.A1(n_1621),
.A2(n_1525),
.B(n_1592),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1640),
.A2(n_1646),
.B(n_1634),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1630),
.B(n_1614),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1628),
.Y(n_1675)
);

AOI321xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1621),
.A2(n_1514),
.A3(n_1506),
.B1(n_1510),
.B2(n_1463),
.C(n_1588),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1628),
.B(n_1627),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1640),
.A2(n_1612),
.B(n_1484),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1639),
.B(n_1516),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1641),
.A2(n_1508),
.B1(n_1504),
.B2(n_1522),
.Y(n_1680)
);

OAI21xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1630),
.A2(n_1633),
.B(n_1639),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1658),
.B(n_1668),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1659),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1671),
.B(n_1642),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1677),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1667),
.A2(n_1641),
.B1(n_1652),
.B2(n_1653),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1660),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1661),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1677),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1663),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1675),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1665),
.B(n_1642),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1665),
.B(n_1643),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1662),
.B(n_1641),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1669),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1681),
.Y(n_1696)
);

NOR2x1_ASAP7_75t_L g1697 ( 
.A(n_1656),
.B(n_1638),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1666),
.B(n_1634),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1657),
.B(n_1643),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1674),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1662),
.B(n_1651),
.Y(n_1701)
);

AOI21xp33_ASAP7_75t_SL g1702 ( 
.A1(n_1686),
.A2(n_1664),
.B(n_1673),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1682),
.B(n_1670),
.Y(n_1703)
);

OAI21xp33_ASAP7_75t_L g1704 ( 
.A1(n_1699),
.A2(n_1672),
.B(n_1633),
.Y(n_1704)
);

OAI211xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1697),
.A2(n_1678),
.B(n_1676),
.C(n_1638),
.Y(n_1705)
);

OAI21xp33_ASAP7_75t_L g1706 ( 
.A1(n_1701),
.A2(n_1678),
.B(n_1641),
.Y(n_1706)
);

OAI221xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1692),
.A2(n_1679),
.B1(n_1647),
.B2(n_1649),
.C(n_1654),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1682),
.B(n_1651),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1685),
.B(n_1293),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1689),
.Y(n_1710)
);

AOI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1694),
.A2(n_1654),
.B1(n_1680),
.B2(n_1655),
.C(n_1652),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1689),
.B(n_1652),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1694),
.A2(n_1655),
.B(n_1631),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1710),
.Y(n_1714)
);

OA22x2_ASAP7_75t_L g1715 ( 
.A1(n_1706),
.A2(n_1685),
.B1(n_1696),
.B2(n_1693),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1708),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1709),
.B(n_1695),
.Y(n_1717)
);

NOR3xp33_ASAP7_75t_L g1718 ( 
.A(n_1702),
.B(n_1691),
.C(n_1684),
.Y(n_1718)
);

NOR3xp33_ASAP7_75t_L g1719 ( 
.A(n_1704),
.B(n_1687),
.C(n_1683),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1712),
.B(n_1700),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_SL g1721 ( 
.A(n_1711),
.B(n_1703),
.C(n_1713),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1707),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1705),
.A2(n_1700),
.B(n_1698),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1710),
.B(n_1698),
.Y(n_1724)
);

CKINVDCx6p67_ASAP7_75t_R g1725 ( 
.A(n_1710),
.Y(n_1725)
);

OAI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1718),
.A2(n_1690),
.B1(n_1688),
.B2(n_1655),
.C(n_1645),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1725),
.B(n_1724),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1720),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1723),
.B(n_1652),
.Y(n_1729)
);

AOI211x1_ASAP7_75t_SL g1730 ( 
.A1(n_1721),
.A2(n_1645),
.B(n_1644),
.C(n_1635),
.Y(n_1730)
);

AOI33xp33_ASAP7_75t_L g1731 ( 
.A1(n_1722),
.A2(n_1635),
.A3(n_1624),
.B1(n_1631),
.B2(n_1644),
.B3(n_1645),
.Y(n_1731)
);

NAND4xp25_ASAP7_75t_L g1732 ( 
.A(n_1717),
.B(n_1624),
.C(n_1631),
.D(n_1635),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1727),
.B(n_1715),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1731),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1729),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1728),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_SL g1737 ( 
.A1(n_1726),
.A2(n_1714),
.B1(n_1716),
.B2(n_1304),
.Y(n_1737)
);

AOI31xp33_ASAP7_75t_L g1738 ( 
.A1(n_1730),
.A2(n_1719),
.A3(n_1649),
.B(n_1647),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1732),
.A2(n_1624),
.B1(n_1644),
.B2(n_1650),
.Y(n_1739)
);

NOR2xp67_ASAP7_75t_SL g1740 ( 
.A(n_1733),
.B(n_1736),
.Y(n_1740)
);

NAND4xp75_ASAP7_75t_L g1741 ( 
.A(n_1734),
.B(n_1495),
.C(n_1246),
.D(n_1259),
.Y(n_1741)
);

NOR3xp33_ASAP7_75t_L g1742 ( 
.A(n_1737),
.B(n_1282),
.C(n_1650),
.Y(n_1742)
);

OAI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1735),
.A2(n_1239),
.B1(n_1238),
.B2(n_1512),
.C(n_1507),
.Y(n_1743)
);

NOR4xp75_ASAP7_75t_SL g1744 ( 
.A(n_1738),
.B(n_1344),
.C(n_1307),
.D(n_1573),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1739),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1741),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1742),
.B(n_1745),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1743),
.B(n_1563),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1747),
.Y(n_1749)
);

NAND4xp25_ASAP7_75t_L g1750 ( 
.A(n_1749),
.B(n_1746),
.C(n_1748),
.D(n_1740),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1750),
.Y(n_1751)
);

AOI22x1_ASAP7_75t_L g1752 ( 
.A1(n_1750),
.A2(n_1748),
.B1(n_1744),
.B2(n_1238),
.Y(n_1752)
);

AOI21xp33_ASAP7_75t_L g1753 ( 
.A1(n_1751),
.A2(n_1344),
.B(n_1281),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1752),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1753),
.A2(n_1327),
.B(n_1259),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1754),
.A2(n_1344),
.B1(n_1281),
.B2(n_1327),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1756),
.A2(n_1246),
.B(n_1281),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1757),
.A2(n_1755),
.B1(n_1260),
.B2(n_1253),
.Y(n_1758)
);

OAI221xp5_ASAP7_75t_R g1759 ( 
.A1(n_1758),
.A2(n_1253),
.B1(n_1260),
.B2(n_1489),
.C(n_1495),
.Y(n_1759)
);

AOI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1759),
.A2(n_1314),
.B(n_1334),
.C(n_1332),
.Y(n_1760)
);


endmodule