module fake_jpeg_16783_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_54),
.Y(n_67)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_43),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_49),
.B1(n_46),
.B2(n_51),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_73),
.B1(n_74),
.B2(n_2),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_78),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_47),
.B1(n_56),
.B2(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_58),
.B1(n_50),
.B2(n_42),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_48),
.B1(n_1),
.B2(n_2),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_9),
.B(n_12),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_3),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_65),
.B1(n_5),
.B2(n_6),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_18),
.B1(n_38),
.B2(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_13),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_4),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_94),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_5),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_90),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_7),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_14),
.C(n_15),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_76),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_94),
.B1(n_93),
.B2(n_87),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_84),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_17),
.B(n_19),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_16),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_107),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_83),
.B(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_110),
.B(n_22),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_20),
.B(n_21),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_95),
.C(n_110),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_112),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_118),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_115),
.C(n_117),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_95),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_97),
.C(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_122),
.B(n_116),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_98),
.B(n_104),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_25),
.C(n_26),
.Y(n_125)
);

OAI211xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_41),
.Y(n_127)
);


endmodule