module fake_netlist_1_12246_n_45 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_45);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_30;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
BUFx10_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_9), .Y(n_18) );
CKINVDCx20_ASAP7_75t_R g19 ( .A(n_6), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_8), .Y(n_20) );
OAI22xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_12), .B(n_11), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_12), .B(n_2), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_13), .Y(n_25) );
BUFx2_ASAP7_75t_L g26 ( .A(n_18), .Y(n_26) );
AND2x4_ASAP7_75t_L g27 ( .A(n_15), .B(n_3), .Y(n_27) );
BUFx3_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_26), .B(n_18), .Y(n_29) );
OAI21xp5_ASAP7_75t_L g30 ( .A1(n_24), .A2(n_17), .B(n_19), .Y(n_30) );
AOI21xp5_ASAP7_75t_L g31 ( .A1(n_24), .A2(n_14), .B(n_16), .Y(n_31) );
AOI22xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_27), .B1(n_23), .B2(n_22), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_28), .B(n_25), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_28), .A2(n_27), .B1(n_25), .B2(n_21), .Y(n_34) );
NAND2xp33_ASAP7_75t_R g35 ( .A(n_33), .B(n_30), .Y(n_35) );
OR2x2_ASAP7_75t_L g36 ( .A(n_34), .B(n_30), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_36), .B(n_32), .Y(n_37) );
AND2x2_ASAP7_75t_L g38 ( .A(n_35), .B(n_27), .Y(n_38) );
AOI22xp5_ASAP7_75t_L g39 ( .A1(n_37), .A2(n_31), .B1(n_27), .B2(n_16), .Y(n_39) );
OAI22xp5_ASAP7_75t_SL g40 ( .A1(n_38), .A2(n_16), .B1(n_5), .B2(n_6), .Y(n_40) );
OAI22xp5_ASAP7_75t_L g41 ( .A1(n_38), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_41) );
OAI22xp5_ASAP7_75t_L g42 ( .A1(n_40), .A2(n_10), .B1(n_4), .B2(n_9), .Y(n_42) );
OR2x2_ASAP7_75t_L g43 ( .A(n_41), .B(n_10), .Y(n_43) );
INVx1_ASAP7_75t_SL g44 ( .A(n_43), .Y(n_44) );
AOI22xp5_ASAP7_75t_L g45 ( .A1(n_44), .A2(n_39), .B1(n_42), .B2(n_40), .Y(n_45) );
endmodule