module real_aes_6752_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_725;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_1), .A2(n_140), .B(n_143), .C(n_223), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_2), .A2(n_169), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g470 ( .A(n_3), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_4), .B(n_199), .Y(n_198) );
AOI21xp33_ASAP7_75t_L g453 ( .A1(n_5), .A2(n_169), .B(n_454), .Y(n_453) );
AND2x6_ASAP7_75t_L g140 ( .A(n_6), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g236 ( .A(n_7), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_8), .B(n_40), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_9), .A2(n_168), .B(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_10), .B(n_152), .Y(n_225) );
INVx1_ASAP7_75t_L g458 ( .A(n_11), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_12), .B(n_193), .Y(n_493) );
INVx1_ASAP7_75t_L g132 ( .A(n_13), .Y(n_132) );
INVx1_ASAP7_75t_L g505 ( .A(n_14), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_15), .A2(n_177), .B(n_258), .C(n_260), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_16), .B(n_199), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_17), .B(n_436), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_18), .B(n_169), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_19), .B(n_183), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_20), .A2(n_193), .B(n_244), .C(n_246), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_21), .B(n_199), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_22), .B(n_152), .Y(n_151) );
AOI22xp33_ASAP7_75t_SL g99 ( .A1(n_23), .A2(n_100), .B1(n_722), .B2(n_727), .Y(n_99) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_24), .A2(n_179), .B(n_260), .C(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_25), .B(n_152), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_26), .Y(n_134) );
INVx1_ASAP7_75t_L g206 ( .A(n_27), .Y(n_206) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_28), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_29), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_30), .B(n_152), .Y(n_471) );
INVx1_ASAP7_75t_L g175 ( .A(n_31), .Y(n_175) );
INVx1_ASAP7_75t_L g448 ( .A(n_32), .Y(n_448) );
INVx2_ASAP7_75t_L g138 ( .A(n_33), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_34), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_35), .A2(n_193), .B(n_194), .C(n_196), .Y(n_192) );
INVxp67_ASAP7_75t_L g178 ( .A(n_36), .Y(n_178) );
CKINVDCx14_ASAP7_75t_R g191 ( .A(n_37), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_38), .A2(n_143), .B(n_205), .C(n_209), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_39), .A2(n_140), .B(n_143), .C(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g447 ( .A(n_41), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_42), .A2(n_154), .B(n_234), .C(n_235), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_43), .B(n_152), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_44), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_45), .Y(n_171) );
INVx1_ASAP7_75t_L g242 ( .A(n_46), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g449 ( .A(n_47), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_48), .B(n_169), .Y(n_495) );
AOI222xp33_ASAP7_75t_L g114 ( .A1(n_49), .A2(n_76), .B1(n_115), .B2(n_709), .C1(n_711), .C2(n_712), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_50), .A2(n_143), .B1(n_246), .B2(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_51), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_52), .Y(n_467) );
CKINVDCx14_ASAP7_75t_R g232 ( .A(n_53), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_54), .A2(n_196), .B(n_234), .C(n_457), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_55), .Y(n_517) );
INVx1_ASAP7_75t_L g455 ( .A(n_56), .Y(n_455) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_57), .A2(n_116), .B1(n_710), .B2(n_719), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_57), .Y(n_719) );
INVx1_ASAP7_75t_L g141 ( .A(n_58), .Y(n_141) );
INVx1_ASAP7_75t_L g131 ( .A(n_59), .Y(n_131) );
INVx1_ASAP7_75t_SL g195 ( .A(n_60), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_61), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_62), .B(n_199), .Y(n_248) );
INVx1_ASAP7_75t_L g147 ( .A(n_63), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_SL g435 ( .A1(n_64), .A2(n_196), .B(n_436), .C(n_437), .Y(n_435) );
INVxp67_ASAP7_75t_L g438 ( .A(n_65), .Y(n_438) );
INVx1_ASAP7_75t_L g725 ( .A(n_66), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_67), .A2(n_169), .B(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_68), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_69), .A2(n_169), .B(n_255), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_70), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_71), .Y(n_107) );
INVx1_ASAP7_75t_L g511 ( .A(n_72), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_73), .A2(n_168), .B(n_170), .Y(n_167) );
CKINVDCx16_ASAP7_75t_R g203 ( .A(n_74), .Y(n_203) );
INVx1_ASAP7_75t_L g256 ( .A(n_75), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_76), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_77), .A2(n_140), .B(n_143), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_78), .A2(n_169), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g259 ( .A(n_79), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_80), .B(n_176), .Y(n_482) );
INVx2_ASAP7_75t_L g129 ( .A(n_81), .Y(n_129) );
INVx1_ASAP7_75t_L g224 ( .A(n_82), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_83), .B(n_436), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_84), .A2(n_140), .B(n_143), .C(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g109 ( .A(n_85), .B(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g422 ( .A(n_85), .B(n_111), .Y(n_422) );
INVx2_ASAP7_75t_L g708 ( .A(n_85), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_86), .A2(n_143), .B(n_146), .C(n_156), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_87), .B(n_161), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_88), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_89), .A2(n_140), .B(n_143), .C(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_90), .Y(n_497) );
INVx1_ASAP7_75t_L g434 ( .A(n_91), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_92), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_93), .B(n_176), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_94), .B(n_127), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_95), .B(n_127), .Y(n_506) );
INVx2_ASAP7_75t_L g245 ( .A(n_96), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_97), .A2(n_169), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_98), .B(n_725), .Y(n_724) );
BUFx3_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_114), .B1(n_715), .B2(n_717), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
BUFx2_ASAP7_75t_L g716 ( .A(n_104), .Y(n_716) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_106), .A2(n_718), .B(n_720), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g721 ( .A(n_108), .Y(n_721) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2x2_ASAP7_75t_L g714 ( .A(n_110), .B(n_708), .Y(n_714) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g707 ( .A(n_111), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
OAI22xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_422), .B1(n_423), .B2(n_705), .Y(n_115) );
INVx2_ASAP7_75t_L g710 ( .A(n_116), .Y(n_710) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_356), .Y(n_116) );
NAND5xp2_ASAP7_75t_L g117 ( .A(n_118), .B(n_285), .C(n_315), .D(n_336), .E(n_342), .Y(n_117) );
AOI221xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_215), .B1(n_249), .B2(n_251), .C(n_262), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_212), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_184), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_SL g336 ( .A1(n_123), .A2(n_200), .B(n_337), .C(n_340), .Y(n_336) );
AND2x2_ASAP7_75t_L g406 ( .A(n_123), .B(n_201), .Y(n_406) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_162), .Y(n_123) );
AND2x2_ASAP7_75t_L g264 ( .A(n_124), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g268 ( .A(n_124), .B(n_265), .Y(n_268) );
OR2x2_ASAP7_75t_L g294 ( .A(n_124), .B(n_201), .Y(n_294) );
AND2x2_ASAP7_75t_L g296 ( .A(n_124), .B(n_187), .Y(n_296) );
AND2x2_ASAP7_75t_L g314 ( .A(n_124), .B(n_186), .Y(n_314) );
INVx1_ASAP7_75t_L g347 ( .A(n_124), .Y(n_347) );
INVx2_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g214 ( .A(n_125), .Y(n_214) );
AND2x2_ASAP7_75t_L g250 ( .A(n_125), .B(n_187), .Y(n_250) );
AND2x2_ASAP7_75t_L g403 ( .A(n_125), .B(n_201), .Y(n_403) );
AO21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_133), .B(n_158), .Y(n_125) );
INVx3_ASAP7_75t_L g199 ( .A(n_126), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_126), .B(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_126), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_SL g484 ( .A(n_126), .B(n_485), .Y(n_484) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_127), .Y(n_188) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_127), .A2(n_432), .B(n_439), .Y(n_431) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g165 ( .A(n_128), .Y(n_165) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_129), .B(n_130), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B(n_142), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_135), .A2(n_161), .B(n_203), .C(n_204), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_135), .A2(n_221), .B(n_222), .Y(n_220) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_135), .A2(n_157), .B1(n_445), .B2(n_449), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_135), .A2(n_467), .B(n_468), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_135), .A2(n_511), .B(n_512), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
AND2x4_ASAP7_75t_L g169 ( .A(n_136), .B(n_140), .Y(n_169) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx1_ASAP7_75t_L g247 ( .A(n_138), .Y(n_247) );
INVx1_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
INVx3_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
INVx1_ASAP7_75t_L g436 ( .A(n_139), .Y(n_436) );
INVx4_ASAP7_75t_SL g157 ( .A(n_140), .Y(n_157) );
BUFx3_ASAP7_75t_L g209 ( .A(n_140), .Y(n_209) );
INVx5_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_144), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .C(n_153), .Y(n_146) );
O2A1O1Ixp5_ASAP7_75t_L g223 ( .A1(n_148), .A2(n_153), .B(n_224), .C(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_149), .A2(n_150), .B1(n_447), .B2(n_448), .Y(n_446) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
INVx4_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
INVx2_ASAP7_75t_L g234 ( .A(n_152), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_153), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_153), .A2(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g260 ( .A(n_155), .Y(n_260) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_SL g170 ( .A1(n_157), .A2(n_171), .B(n_172), .C(n_173), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_157), .A2(n_172), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_SL g231 ( .A1(n_157), .A2(n_172), .B(n_232), .C(n_233), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_157), .A2(n_172), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g255 ( .A1(n_157), .A2(n_172), .B(n_256), .C(n_257), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g433 ( .A1(n_157), .A2(n_172), .B(n_434), .C(n_435), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_157), .A2(n_172), .B(n_455), .C(n_456), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_157), .A2(n_172), .B(n_502), .C(n_503), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx1_ASAP7_75t_L g183 ( .A(n_160), .Y(n_183) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_160), .A2(n_489), .B(n_496), .Y(n_488) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g219 ( .A(n_161), .Y(n_219) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_161), .A2(n_230), .B(n_237), .Y(n_229) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_161), .A2(n_500), .B(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g284 ( .A(n_162), .B(n_185), .Y(n_284) );
OR2x2_ASAP7_75t_L g288 ( .A(n_162), .B(n_201), .Y(n_288) );
AND2x2_ASAP7_75t_L g313 ( .A(n_162), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g360 ( .A(n_162), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_162), .B(n_322), .Y(n_408) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_166), .B(n_181), .Y(n_162) );
INVx1_ASAP7_75t_L g266 ( .A(n_163), .Y(n_266) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_163), .A2(n_510), .B(n_516), .Y(n_509) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_SL g478 ( .A1(n_164), .A2(n_479), .B(n_480), .Y(n_478) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_165), .A2(n_444), .B(n_450), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_165), .B(n_451), .Y(n_450) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_165), .A2(n_466), .B(n_473), .Y(n_465) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_167), .A2(n_182), .B(n_266), .Y(n_265) );
BUFx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_174), .B(n_180), .Y(n_173) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B1(n_178), .B2(n_179), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_176), .A2(n_206), .B(n_207), .C(n_208), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_176), .A2(n_470), .B(n_471), .C(n_472), .Y(n_469) );
INVx5_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_177), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_177), .B(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_177), .B(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_179), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_179), .B(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_179), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g208 ( .A(n_180), .Y(n_208) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OAI322xp33_ASAP7_75t_L g409 ( .A1(n_184), .A2(n_345), .A3(n_368), .B1(n_389), .B2(n_410), .C1(n_412), .C2(n_413), .Y(n_409) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_185), .B(n_265), .Y(n_412) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_200), .Y(n_185) );
AND2x2_ASAP7_75t_L g213 ( .A(n_186), .B(n_214), .Y(n_213) );
AND2x4_ASAP7_75t_L g281 ( .A(n_186), .B(n_201), .Y(n_281) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g322 ( .A(n_187), .B(n_201), .Y(n_322) );
AND2x2_ASAP7_75t_L g366 ( .A(n_187), .B(n_200), .Y(n_366) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_198), .Y(n_187) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_188), .A2(n_240), .B(n_248), .Y(n_239) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_188), .A2(n_254), .B(n_261), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_193), .B(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_197), .Y(n_494) );
OA21x2_ASAP7_75t_L g452 ( .A1(n_199), .A2(n_453), .B(n_459), .Y(n_452) );
AND2x2_ASAP7_75t_L g249 ( .A(n_200), .B(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g267 ( .A(n_200), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_200), .B(n_296), .Y(n_420) );
INVx3_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g212 ( .A(n_201), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_201), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g334 ( .A(n_201), .B(n_265), .Y(n_334) );
AND2x2_ASAP7_75t_L g361 ( .A(n_201), .B(n_296), .Y(n_361) );
OR2x2_ASAP7_75t_L g417 ( .A(n_201), .B(n_268), .Y(n_417) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_210), .Y(n_201) );
INVx1_ASAP7_75t_SL g303 ( .A(n_212), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_213), .B(n_334), .Y(n_335) );
AND2x2_ASAP7_75t_L g369 ( .A(n_213), .B(n_359), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_213), .B(n_292), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_213), .B(n_414), .Y(n_413) );
OAI31xp33_ASAP7_75t_L g387 ( .A1(n_215), .A2(n_249), .A3(n_388), .B(n_390), .Y(n_387) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_228), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_216), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g370 ( .A(n_216), .B(n_305), .Y(n_370) );
OR2x2_ASAP7_75t_L g377 ( .A(n_216), .B(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g389 ( .A(n_216), .B(n_278), .Y(n_389) );
CKINVDCx16_ASAP7_75t_R g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g323 ( .A(n_217), .B(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g251 ( .A(n_218), .B(n_252), .Y(n_251) );
INVx4_ASAP7_75t_L g272 ( .A(n_218), .Y(n_272) );
AND2x2_ASAP7_75t_L g309 ( .A(n_218), .B(n_253), .Y(n_309) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_226), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_219), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_219), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_219), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g308 ( .A(n_228), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g378 ( .A(n_228), .Y(n_378) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_238), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_229), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g278 ( .A(n_229), .B(n_239), .Y(n_278) );
INVx2_ASAP7_75t_L g298 ( .A(n_229), .Y(n_298) );
AND2x2_ASAP7_75t_L g312 ( .A(n_229), .B(n_239), .Y(n_312) );
AND2x2_ASAP7_75t_L g319 ( .A(n_229), .B(n_275), .Y(n_319) );
BUFx3_ASAP7_75t_L g329 ( .A(n_229), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_229), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g274 ( .A(n_238), .Y(n_274) );
AND2x2_ASAP7_75t_L g282 ( .A(n_238), .B(n_272), .Y(n_282) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g252 ( .A(n_239), .B(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_239), .Y(n_306) );
INVx2_ASAP7_75t_L g472 ( .A(n_246), .Y(n_472) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_SL g289 ( .A(n_250), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_250), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_250), .B(n_359), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_251), .B(n_329), .Y(n_382) );
INVx1_ASAP7_75t_SL g416 ( .A(n_251), .Y(n_416) );
INVx1_ASAP7_75t_SL g324 ( .A(n_252), .Y(n_324) );
INVx1_ASAP7_75t_SL g275 ( .A(n_253), .Y(n_275) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_253), .Y(n_286) );
OR2x2_ASAP7_75t_L g297 ( .A(n_253), .B(n_272), .Y(n_297) );
AND2x2_ASAP7_75t_L g311 ( .A(n_253), .B(n_272), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_253), .B(n_301), .Y(n_363) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_267), .B(n_269), .C(n_280), .Y(n_262) );
AOI31xp33_ASAP7_75t_L g379 ( .A1(n_263), .A2(n_380), .A3(n_381), .B(n_382), .Y(n_379) );
AND2x2_ASAP7_75t_L g352 ( .A(n_264), .B(n_281), .Y(n_352) );
BUFx3_ASAP7_75t_L g292 ( .A(n_265), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_265), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g328 ( .A(n_265), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_265), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g283 ( .A(n_268), .Y(n_283) );
OAI222xp33_ASAP7_75t_L g392 ( .A1(n_268), .A2(n_393), .B1(n_396), .B2(n_397), .C1(n_398), .C2(n_399), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_276), .Y(n_269) );
INVx1_ASAP7_75t_L g398 ( .A(n_270), .Y(n_398) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_272), .B(n_275), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_272), .B(n_298), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_272), .B(n_273), .Y(n_368) );
INVx1_ASAP7_75t_L g419 ( .A(n_272), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_273), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g421 ( .A(n_273), .Y(n_421) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g301 ( .A(n_274), .Y(n_301) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_275), .Y(n_344) );
AOI32xp33_ASAP7_75t_L g280 ( .A1(n_276), .A2(n_281), .A3(n_282), .B1(n_283), .B2(n_284), .Y(n_280) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_278), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g355 ( .A(n_278), .Y(n_355) );
OR2x2_ASAP7_75t_L g396 ( .A(n_278), .B(n_297), .Y(n_396) );
INVx1_ASAP7_75t_L g332 ( .A(n_279), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_281), .B(n_292), .Y(n_317) );
INVx3_ASAP7_75t_L g326 ( .A(n_281), .Y(n_326) );
AOI322xp5_ASAP7_75t_L g342 ( .A1(n_281), .A2(n_326), .A3(n_343), .B1(n_345), .B2(n_348), .C1(n_352), .C2(n_353), .Y(n_342) );
AND2x2_ASAP7_75t_L g318 ( .A(n_282), .B(n_319), .Y(n_318) );
INVxp67_ASAP7_75t_L g395 ( .A(n_282), .Y(n_395) );
A2O1A1O1Ixp25_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_290), .C(n_298), .D(n_299), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_286), .B(n_329), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g299 ( .A1(n_288), .A2(n_300), .B1(n_303), .B2(n_304), .C(n_307), .Y(n_299) );
INVx1_ASAP7_75t_SL g414 ( .A(n_288), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_295), .B(n_297), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_292), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OAI221xp5_ASAP7_75t_SL g384 ( .A1(n_294), .A2(n_378), .B1(n_385), .B2(n_386), .C(n_387), .Y(n_384) );
OAI222xp33_ASAP7_75t_L g415 ( .A1(n_295), .A2(n_416), .B1(n_417), .B2(n_418), .C1(n_420), .C2(n_421), .Y(n_415) );
AND2x2_ASAP7_75t_L g373 ( .A(n_296), .B(n_359), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_296), .A2(n_311), .B(n_358), .Y(n_385) );
INVx1_ASAP7_75t_L g399 ( .A(n_296), .Y(n_399) );
INVx2_ASAP7_75t_SL g302 ( .A(n_297), .Y(n_302) );
AND2x2_ASAP7_75t_L g305 ( .A(n_298), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_SL g339 ( .A(n_301), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_301), .B(n_311), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_302), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_302), .B(n_312), .Y(n_341) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI21xp5_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_310), .B(n_313), .Y(n_307) );
INVx1_ASAP7_75t_SL g325 ( .A(n_309), .Y(n_325) );
AND2x2_ASAP7_75t_L g372 ( .A(n_309), .B(n_355), .Y(n_372) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g411 ( .A(n_311), .B(n_329), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_312), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g397 ( .A(n_313), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_318), .B1(n_320), .B2(n_327), .C(n_330), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_323), .B1(n_325), .B2(n_326), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI22xp33_ASAP7_75t_L g330 ( .A1(n_324), .A2(n_331), .B1(n_333), .B2(n_335), .Y(n_330) );
OR2x2_ASAP7_75t_L g401 ( .A(n_325), .B(n_329), .Y(n_401) );
OR2x2_ASAP7_75t_L g404 ( .A(n_325), .B(n_339), .Y(n_404) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_346), .A2(n_401), .B1(n_402), .B2(n_404), .C(n_405), .Y(n_400) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND3xp33_ASAP7_75t_SL g356 ( .A(n_357), .B(n_371), .C(n_383), .Y(n_356) );
AOI222xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_362), .B1(n_364), .B2(n_367), .C1(n_369), .C2(n_370), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_359), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g381 ( .A(n_361), .Y(n_381) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_374), .B2(n_376), .C(n_379), .Y(n_371) );
INVx1_ASAP7_75t_L g386 ( .A(n_372), .Y(n_386) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI21xp33_ASAP7_75t_L g405 ( .A1(n_376), .A2(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
NOR5xp2_ASAP7_75t_L g383 ( .A(n_384), .B(n_392), .C(n_400), .D(n_409), .E(n_415), .Y(n_383) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI22xp5_ASAP7_75t_SL g709 ( .A1(n_422), .A2(n_424), .B1(n_705), .B2(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_SL g424 ( .A(n_425), .B(n_642), .Y(n_424) );
NOR4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_572), .C(n_603), .D(n_622), .Y(n_425) );
NAND4xp25_ASAP7_75t_L g426 ( .A(n_427), .B(n_530), .C(n_545), .D(n_563), .Y(n_426) );
AOI222xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_475), .B1(n_507), .B2(n_518), .C1(n_523), .C2(n_525), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_460), .Y(n_428) );
INVx1_ASAP7_75t_L g586 ( .A(n_429), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_440), .Y(n_429) );
AND2x2_ASAP7_75t_L g461 ( .A(n_430), .B(n_452), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_430), .B(n_464), .Y(n_615) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g522 ( .A(n_431), .B(n_442), .Y(n_522) );
AND2x2_ASAP7_75t_L g531 ( .A(n_431), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g557 ( .A(n_431), .Y(n_557) );
AND2x2_ASAP7_75t_L g578 ( .A(n_431), .B(n_442), .Y(n_578) );
BUFx2_ASAP7_75t_L g601 ( .A(n_431), .Y(n_601) );
AND2x2_ASAP7_75t_L g625 ( .A(n_431), .B(n_443), .Y(n_625) );
AND2x2_ASAP7_75t_L g689 ( .A(n_431), .B(n_452), .Y(n_689) );
AND2x2_ASAP7_75t_L g590 ( .A(n_440), .B(n_521), .Y(n_590) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_441), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_452), .Y(n_441) );
OR2x2_ASAP7_75t_L g550 ( .A(n_442), .B(n_465), .Y(n_550) );
AND2x2_ASAP7_75t_L g562 ( .A(n_442), .B(n_521), .Y(n_562) );
BUFx2_ASAP7_75t_L g694 ( .A(n_442), .Y(n_694) );
INVx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g463 ( .A(n_443), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g544 ( .A(n_443), .B(n_465), .Y(n_544) );
AND2x2_ASAP7_75t_L g597 ( .A(n_443), .B(n_452), .Y(n_597) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_443), .Y(n_633) );
AND2x2_ASAP7_75t_L g520 ( .A(n_452), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_SL g532 ( .A(n_452), .Y(n_532) );
INVx2_ASAP7_75t_L g543 ( .A(n_452), .Y(n_543) );
BUFx2_ASAP7_75t_L g567 ( .A(n_452), .Y(n_567) );
AND2x2_ASAP7_75t_SL g624 ( .A(n_452), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
AOI332xp33_ASAP7_75t_L g545 ( .A1(n_461), .A2(n_546), .A3(n_550), .B1(n_551), .B2(n_555), .B3(n_558), .C1(n_559), .C2(n_561), .Y(n_545) );
NAND2x1_ASAP7_75t_L g630 ( .A(n_461), .B(n_521), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_461), .B(n_535), .Y(n_681) );
A2O1A1Ixp33_ASAP7_75t_SL g563 ( .A1(n_462), .A2(n_564), .B(n_567), .C(n_568), .Y(n_563) );
AND2x2_ASAP7_75t_L g702 ( .A(n_462), .B(n_543), .Y(n_702) );
INVx3_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g599 ( .A(n_463), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g604 ( .A(n_463), .B(n_601), .Y(n_604) );
INVx1_ASAP7_75t_L g535 ( .A(n_464), .Y(n_535) );
AND2x2_ASAP7_75t_L g638 ( .A(n_464), .B(n_597), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_464), .B(n_578), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_464), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_464), .B(n_556), .Y(n_664) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx3_ASAP7_75t_L g521 ( .A(n_465), .Y(n_521) );
OAI31xp33_ASAP7_75t_L g703 ( .A1(n_475), .A2(n_624), .A3(n_631), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
AND2x2_ASAP7_75t_L g507 ( .A(n_476), .B(n_508), .Y(n_507) );
NAND2x1_ASAP7_75t_SL g526 ( .A(n_476), .B(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_476), .Y(n_613) );
AND2x2_ASAP7_75t_L g618 ( .A(n_476), .B(n_529), .Y(n_618) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_477), .A2(n_531), .B(n_533), .C(n_536), .Y(n_530) );
OR2x2_ASAP7_75t_L g547 ( .A(n_477), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g560 ( .A(n_477), .Y(n_560) );
AND2x2_ASAP7_75t_L g566 ( .A(n_477), .B(n_509), .Y(n_566) );
INVx2_ASAP7_75t_L g584 ( .A(n_477), .Y(n_584) );
AND2x2_ASAP7_75t_L g595 ( .A(n_477), .B(n_549), .Y(n_595) );
AND2x2_ASAP7_75t_L g627 ( .A(n_477), .B(n_585), .Y(n_627) );
AND2x2_ASAP7_75t_L g631 ( .A(n_477), .B(n_554), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_477), .B(n_486), .Y(n_636) );
AND2x2_ASAP7_75t_L g670 ( .A(n_477), .B(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_477), .B(n_573), .Y(n_704) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_484), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_486), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g612 ( .A(n_486), .Y(n_612) );
AND2x2_ASAP7_75t_L g674 ( .A(n_486), .B(n_595), .Y(n_674) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
OR2x2_ASAP7_75t_L g528 ( .A(n_487), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g538 ( .A(n_487), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_487), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g646 ( .A(n_487), .Y(n_646) );
AND2x2_ASAP7_75t_L g663 ( .A(n_487), .B(n_509), .Y(n_663) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g554 ( .A(n_488), .B(n_498), .Y(n_554) );
AND2x2_ASAP7_75t_L g583 ( .A(n_488), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g594 ( .A(n_488), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_488), .B(n_549), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_495), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g508 ( .A(n_499), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g529 ( .A(n_499), .Y(n_529) );
AND2x2_ASAP7_75t_L g585 ( .A(n_499), .B(n_549), .Y(n_585) );
INVx1_ASAP7_75t_L g687 ( .A(n_507), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_508), .Y(n_691) );
INVx2_ASAP7_75t_L g549 ( .A(n_509), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_522), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_520), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_520), .B(n_625), .Y(n_683) );
OR2x2_ASAP7_75t_L g524 ( .A(n_521), .B(n_522), .Y(n_524) );
INVx1_ASAP7_75t_SL g576 ( .A(n_521), .Y(n_576) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_527), .A2(n_580), .B1(n_582), .B2(n_586), .C(n_587), .Y(n_579) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g607 ( .A(n_528), .B(n_571), .Y(n_607) );
INVx2_ASAP7_75t_L g539 ( .A(n_529), .Y(n_539) );
INVx1_ASAP7_75t_L g565 ( .A(n_529), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_529), .B(n_549), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_529), .B(n_552), .Y(n_659) );
INVx1_ASAP7_75t_L g667 ( .A(n_529), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_531), .B(n_535), .Y(n_581) );
AND2x4_ASAP7_75t_L g556 ( .A(n_532), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g669 ( .A(n_535), .B(n_625), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_538), .B(n_570), .Y(n_569) );
INVxp67_ASAP7_75t_L g677 ( .A(n_539), .Y(n_677) );
INVxp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g577 ( .A(n_543), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g649 ( .A(n_543), .B(n_625), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_543), .B(n_562), .Y(n_655) );
AOI322xp5_ASAP7_75t_L g609 ( .A1(n_544), .A2(n_578), .A3(n_585), .B1(n_610), .B2(n_613), .C1(n_614), .C2(n_616), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_544), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g675 ( .A(n_547), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g621 ( .A(n_548), .Y(n_621) );
INVx2_ASAP7_75t_L g552 ( .A(n_549), .Y(n_552) );
INVx1_ASAP7_75t_L g611 ( .A(n_549), .Y(n_611) );
CKINVDCx16_ASAP7_75t_R g558 ( .A(n_550), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g647 ( .A(n_552), .B(n_560), .Y(n_647) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g559 ( .A(n_554), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g602 ( .A(n_554), .B(n_595), .Y(n_602) );
AND2x2_ASAP7_75t_L g606 ( .A(n_554), .B(n_566), .Y(n_606) );
OAI21xp33_ASAP7_75t_SL g616 ( .A1(n_555), .A2(n_617), .B(n_619), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g686 ( .A1(n_555), .A2(n_687), .B1(n_688), .B2(n_690), .Y(n_686) );
INVx3_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g561 ( .A(n_556), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_556), .B(n_576), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_558), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g698 ( .A(n_565), .Y(n_698) );
INVx4_ASAP7_75t_L g571 ( .A(n_566), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_566), .B(n_593), .Y(n_641) );
INVx1_ASAP7_75t_SL g653 ( .A(n_567), .Y(n_653) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR2xp67_ASAP7_75t_L g666 ( .A(n_571), .B(n_667), .Y(n_666) );
OAI211xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_574), .B(n_579), .C(n_596), .Y(n_572) );
OAI221xp5_ASAP7_75t_SL g692 ( .A1(n_574), .A2(n_612), .B1(n_691), .B2(n_693), .C(n_695), .Y(n_692) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_576), .B(n_689), .Y(n_688) );
OAI31xp33_ASAP7_75t_L g668 ( .A1(n_577), .A2(n_654), .A3(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g608 ( .A(n_578), .Y(n_608) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g658 ( .A(n_583), .Y(n_658) );
AND2x2_ASAP7_75t_L g671 ( .A(n_585), .B(n_594), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_591), .Y(n_587) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_595), .B(n_698), .Y(n_697) );
OAI21xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_602), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI221xp5_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_605), .B1(n_607), .B2(n_608), .C(n_609), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_604), .A2(n_673), .B(n_675), .C(n_678), .Y(n_672) );
CKINVDCx16_ASAP7_75t_R g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_607), .B(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g634 ( .A(n_615), .Y(n_634) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g620 ( .A(n_618), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g662 ( .A(n_618), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI211xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B(n_628), .C(n_637), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_626), .A2(n_636), .B1(n_700), .B2(n_701), .C(n_703), .Y(n_699) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B1(n_632), .B2(n_635), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_SL g700 ( .A(n_639), .Y(n_700) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NOR4xp25_ASAP7_75t_L g642 ( .A(n_643), .B(n_672), .C(n_692), .D(n_699), .Y(n_642) );
OAI211xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_648), .B(n_650), .C(n_668), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVxp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B(n_656), .C(n_660), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g679 ( .A(n_657), .Y(n_679) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
OR2x2_ASAP7_75t_L g690 ( .A(n_658), .B(n_691), .Y(n_690) );
OAI21xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B(n_665), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_682), .B2(n_684), .C(n_686), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_689), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx3_ASAP7_75t_SL g726 ( .A(n_714), .Y(n_726) );
INVx2_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g728 ( .A(n_723), .Y(n_728) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
endmodule