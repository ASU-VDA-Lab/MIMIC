module fake_netlist_6_2846_n_1982 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1982);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1982;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_41),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_130),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_68),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_97),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_61),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_158),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_101),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_73),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_10),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_52),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_32),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_145),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_92),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_175),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_54),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_108),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_35),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_141),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_28),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_112),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_69),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_77),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_168),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_182),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_140),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_143),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_110),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_134),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_106),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_123),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_65),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_94),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_122),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_124),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_69),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_135),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_60),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_71),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_65),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_116),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_120),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_6),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_99),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_72),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_32),
.Y(n_249)
);

BUFx2_ASAP7_75t_SL g250 ( 
.A(n_142),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_153),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_88),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_128),
.Y(n_254)
);

BUFx8_ASAP7_75t_SL g255 ( 
.A(n_177),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_186),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_104),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_192),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_139),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_16),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_150),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_76),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_100),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_163),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_190),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_87),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_137),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_48),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_6),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_76),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_52),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_165),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_38),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_91),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_63),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_174),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_7),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_2),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_49),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_152),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_151),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_25),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_12),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_162),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_51),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_67),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_185),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_68),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_38),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_29),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_46),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_20),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_114),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_48),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_90),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_67),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_51),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_178),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_180),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_95),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_41),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_144),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_119),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_138),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_0),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_115),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_28),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_9),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_42),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_31),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_154),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_46),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_63),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_66),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_125),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_44),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_79),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_156),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_74),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_4),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_43),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_33),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_131),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_169),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_89),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_1),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_29),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_57),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_18),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_30),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_107),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_34),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_11),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_64),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_136),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_1),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_7),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_33),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_113),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_82),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_183),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_167),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_34),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_66),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_14),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_37),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_194),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_85),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_73),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_105),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_31),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_118),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_56),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_18),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_111),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_55),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_62),
.Y(n_358)
);

BUFx8_ASAP7_75t_SL g359 ( 
.A(n_30),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_155),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_42),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_64),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_27),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_9),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_109),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_62),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_21),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_22),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_117),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_70),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_16),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_84),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_44),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_166),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_189),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_83),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_127),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_70),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_2),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_98),
.Y(n_380)
);

BUFx8_ASAP7_75t_SL g381 ( 
.A(n_129),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_58),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_43),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_102),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_57),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_20),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_226),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_359),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_287),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_270),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_270),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_286),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_286),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_298),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_298),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_384),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_257),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_195),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_195),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_199),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_0),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_208),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_199),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_265),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_R g405 ( 
.A(n_208),
.B(n_3),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_325),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_377),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_200),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_384),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_255),
.Y(n_410)
);

INVxp33_ASAP7_75t_SL g411 ( 
.A(n_382),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_200),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_382),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_381),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_316),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_201),
.B(n_3),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_201),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_308),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_205),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_196),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_308),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_328),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_276),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_205),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_206),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_206),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_328),
.Y(n_427)
);

BUFx6f_ASAP7_75t_SL g428 ( 
.A(n_280),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_334),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_334),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_212),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_219),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_219),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_326),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_350),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_229),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_350),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_212),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_236),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_207),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_229),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_216),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_218),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_230),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_220),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_230),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_231),
.B(n_4),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_302),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_302),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_222),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_R g451 ( 
.A(n_197),
.B(n_5),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_231),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_232),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_233),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_232),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_238),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_242),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_244),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_302),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_244),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_316),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_245),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_245),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_247),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_243),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_374),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_247),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_311),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_249),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_196),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_311),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_311),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_252),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_252),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_267),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_246),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_267),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_198),
.B(n_5),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_262),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_272),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_269),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_272),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_374),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_271),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_198),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_264),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_275),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_203),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_282),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_278),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_279),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_283),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_290),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_448),
.B(n_322),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_415),
.B(n_289),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_431),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_431),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_431),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_411),
.A2(n_315),
.B1(n_335),
.B2(n_295),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_473),
.B(n_223),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_387),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_431),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_396),
.B(n_204),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_438),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_409),
.B(n_213),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_398),
.B(n_223),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_438),
.B(n_215),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_438),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_438),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_468),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_449),
.B(n_210),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_468),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_471),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_399),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_410),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_471),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_414),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_488),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_397),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_389),
.B(n_280),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_459),
.B(n_224),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_472),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_388),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_388),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_400),
.B(n_322),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_403),
.B(n_225),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_472),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_404),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_423),
.B(n_210),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_408),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_412),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_435),
.B(n_321),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_419),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_424),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_406),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_425),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_426),
.B(n_322),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_432),
.B(n_433),
.Y(n_541)
);

OA21x2_ASAP7_75t_L g542 ( 
.A1(n_436),
.A2(n_347),
.B(n_339),
.Y(n_542)
);

OA21x2_ASAP7_75t_L g543 ( 
.A1(n_441),
.A2(n_347),
.B(n_339),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_390),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_390),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_407),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_440),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_391),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_391),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_440),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_444),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_466),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_443),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_452),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_453),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_434),
.B(n_339),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_392),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_455),
.B(n_227),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_458),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_SL g561 ( 
.A(n_405),
.B(n_344),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_460),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_462),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_463),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_443),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_445),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_483),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_442),
.B(n_211),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_464),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_467),
.B(n_228),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_445),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_474),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_450),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_475),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_392),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_477),
.Y(n_576)
);

AND3x1_ASAP7_75t_L g577 ( 
.A(n_416),
.B(n_378),
.C(n_347),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_480),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_482),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_501),
.A2(n_447),
.B1(n_413),
.B2(n_402),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_505),
.B(n_486),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_512),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_533),
.Y(n_583)
);

BUFx8_ASAP7_75t_SL g584 ( 
.A(n_502),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_512),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_506),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_533),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_536),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_513),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_512),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_L g591 ( 
.A(n_505),
.B(n_212),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_506),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_512),
.Y(n_593)
);

AND3x2_ASAP7_75t_L g594 ( 
.A(n_544),
.B(n_376),
.C(n_304),
.Y(n_594)
);

OR2x6_ASAP7_75t_L g595 ( 
.A(n_494),
.B(n_478),
.Y(n_595)
);

AND2x6_ASAP7_75t_L g596 ( 
.A(n_501),
.B(n_304),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_536),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_512),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_507),
.B(n_439),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_506),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_512),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_507),
.B(n_389),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_534),
.B(n_469),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_539),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_539),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_509),
.B(n_489),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_L g607 ( 
.A(n_523),
.B(n_304),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_523),
.B(n_450),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_506),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_520),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_516),
.Y(n_611)
);

INVx4_ASAP7_75t_SL g612 ( 
.A(n_506),
.Y(n_612)
);

INVx5_ASAP7_75t_L g613 ( 
.A(n_506),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_501),
.B(n_454),
.Y(n_614)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_534),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_515),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_515),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_516),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_568),
.B(n_461),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_513),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_515),
.Y(n_621)
);

NOR2x1p5_ASAP7_75t_L g622 ( 
.A(n_525),
.B(n_393),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_501),
.B(n_454),
.Y(n_623)
);

AND2x2_ASAP7_75t_SL g624 ( 
.A(n_577),
.B(n_376),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_511),
.Y(n_625)
);

INVx4_ASAP7_75t_SL g626 ( 
.A(n_510),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_551),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_551),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_531),
.A2(n_401),
.B1(n_378),
.B2(n_478),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_515),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_494),
.B(n_456),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_511),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_521),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_577),
.B(n_234),
.Y(n_634)
);

BUFx4f_ASAP7_75t_L g635 ( 
.A(n_542),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_561),
.A2(n_394),
.B1(n_395),
.B2(n_393),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_494),
.B(n_528),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g638 ( 
.A(n_528),
.B(n_376),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_557),
.B(n_234),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_559),
.B(n_456),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_526),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_531),
.B(n_481),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_557),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_553),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_553),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_516),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_511),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_555),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_570),
.B(n_457),
.Y(n_649)
);

OR2x6_ASAP7_75t_L g650 ( 
.A(n_544),
.B(n_250),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_570),
.B(n_235),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_542),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_510),
.B(n_465),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_511),
.B(n_476),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_496),
.B(n_476),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_SL g656 ( 
.A(n_522),
.B(n_451),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_575),
.B(n_250),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_495),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_555),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_496),
.B(n_497),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_SL g661 ( 
.A(n_500),
.B(n_357),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_556),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_547),
.B(n_479),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_556),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_497),
.B(n_479),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_575),
.B(n_481),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_498),
.B(n_499),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_514),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_508),
.A2(n_378),
.B1(n_368),
.B2(n_354),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_535),
.B(n_235),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_560),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_545),
.B(n_484),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_560),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_542),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_495),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_542),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_542),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_550),
.B(n_484),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_508),
.A2(n_363),
.B1(n_209),
.B2(n_202),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_508),
.A2(n_363),
.B1(n_209),
.B2(n_202),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_562),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_514),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_562),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_554),
.A2(n_422),
.B1(n_418),
.B2(n_421),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_565),
.B(n_487),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_545),
.B(n_487),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_543),
.Y(n_687)
);

INVx5_ASAP7_75t_L g688 ( 
.A(n_537),
.Y(n_688)
);

AND2x2_ASAP7_75t_SL g689 ( 
.A(n_543),
.B(n_380),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_548),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_498),
.B(n_490),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_548),
.B(n_420),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_499),
.B(n_490),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_564),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_530),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_535),
.B(n_380),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_566),
.B(n_491),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_L g698 ( 
.A(n_537),
.B(n_380),
.Y(n_698)
);

OR2x6_ASAP7_75t_L g699 ( 
.A(n_549),
.B(n_558),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_543),
.Y(n_700)
);

AND3x4_ASAP7_75t_L g701 ( 
.A(n_500),
.B(n_395),
.C(n_394),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_564),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_518),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_518),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_503),
.B(n_492),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_574),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_549),
.B(n_418),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_524),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_504),
.B(n_492),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_574),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_576),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_543),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_524),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_504),
.B(n_493),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_529),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_538),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_535),
.B(n_493),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_535),
.B(n_217),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_558),
.B(n_421),
.Y(n_719)
);

AND2x6_ASAP7_75t_L g720 ( 
.A(n_527),
.B(n_282),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_543),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_541),
.B(n_470),
.Y(n_722)
);

AND3x1_ASAP7_75t_L g723 ( 
.A(n_527),
.B(n_248),
.C(n_241),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_571),
.B(n_422),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_527),
.A2(n_352),
.B1(n_241),
.B2(n_248),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_573),
.B(n_427),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_540),
.A2(n_284),
.B1(n_379),
.B2(n_373),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_583),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_587),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_637),
.B(n_537),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_588),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_668),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_643),
.B(n_537),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_635),
.A2(n_676),
.B(n_652),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_584),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_589),
.A2(n_620),
.B1(n_643),
.B2(n_623),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_668),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_589),
.B(n_620),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_631),
.B(n_427),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_606),
.B(n_537),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_603),
.B(n_429),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_625),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_624),
.A2(n_333),
.B1(n_323),
.B2(n_352),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_614),
.A2(n_214),
.B1(n_372),
.B2(n_318),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_642),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_682),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_595),
.A2(n_372),
.B1(n_348),
.B2(n_343),
.Y(n_747)
);

NAND3xp33_ASAP7_75t_L g748 ( 
.A(n_580),
.B(n_430),
.C(n_429),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_625),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_634),
.A2(n_541),
.B(n_578),
.C(n_576),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_724),
.B(n_517),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_608),
.B(n_569),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_635),
.B(n_674),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_640),
.B(n_430),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_635),
.A2(n_676),
.B(n_652),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_584),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_666),
.B(n_437),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_674),
.B(n_687),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_674),
.B(n_569),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_677),
.B(n_569),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_699),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_682),
.Y(n_762)
);

BUFx12f_ASAP7_75t_L g763 ( 
.A(n_641),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_677),
.A2(n_563),
.B(n_532),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_718),
.B(n_569),
.Y(n_765)
);

INVx8_ASAP7_75t_L g766 ( 
.A(n_650),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_649),
.B(n_581),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_597),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_655),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_719),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_674),
.B(n_687),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_SL g772 ( 
.A(n_610),
.B(n_519),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_703),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_687),
.B(n_569),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_687),
.B(n_221),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_634),
.A2(n_303),
.B(n_348),
.C(n_356),
.Y(n_776)
);

NOR2x1p5_ASAP7_75t_L g777 ( 
.A(n_602),
.B(n_437),
.Y(n_777)
);

AOI221xp5_ASAP7_75t_L g778 ( 
.A1(n_661),
.A2(n_485),
.B1(n_366),
.B2(n_277),
.C(n_284),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_625),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_721),
.B(n_532),
.Y(n_780)
);

O2A1O1Ixp5_ASAP7_75t_L g781 ( 
.A1(n_651),
.A2(n_700),
.B(n_639),
.C(n_670),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_703),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_604),
.Y(n_783)
);

INVx8_ASAP7_75t_L g784 ( 
.A(n_650),
.Y(n_784)
);

NOR2x1p5_ASAP7_75t_L g785 ( 
.A(n_707),
.B(n_291),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_605),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_656),
.A2(n_259),
.B1(n_261),
.B2(n_281),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_627),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_624),
.B(n_572),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_704),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_689),
.B(n_572),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_629),
.A2(n_712),
.B(n_656),
.C(n_607),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_615),
.B(n_672),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_704),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_628),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_717),
.B(n_578),
.C(n_297),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_689),
.B(n_365),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_610),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_700),
.B(n_572),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_712),
.B(n_700),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_708),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_599),
.B(n_579),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_717),
.A2(n_351),
.B1(n_312),
.B2(n_239),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_708),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_713),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_644),
.B(n_579),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_645),
.B(n_579),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_648),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_692),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_611),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_713),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_619),
.B(n_428),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_659),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_591),
.B(n_306),
.C(n_292),
.Y(n_814)
);

INVx5_ASAP7_75t_L g815 ( 
.A(n_596),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_722),
.B(n_428),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_722),
.B(n_428),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_611),
.B(n_237),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_722),
.B(n_309),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_618),
.B(n_240),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_662),
.B(n_540),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_664),
.B(n_540),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_671),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_715),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_646),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_673),
.Y(n_826)
);

HB1xp67_ASAP7_75t_SL g827 ( 
.A(n_663),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_681),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_654),
.A2(n_529),
.B(n_305),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_665),
.B(n_251),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_722),
.B(n_310),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_632),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_683),
.B(n_694),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_702),
.B(n_303),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_706),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_710),
.B(n_305),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_711),
.B(n_595),
.Y(n_837)
);

NOR3xp33_ASAP7_75t_L g838 ( 
.A(n_661),
.B(n_320),
.C(n_313),
.Y(n_838)
);

NOR3xp33_ASAP7_75t_L g839 ( 
.A(n_678),
.B(n_329),
.C(n_327),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_715),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_691),
.B(n_253),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_596),
.B(n_318),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_SL g843 ( 
.A1(n_701),
.A2(n_567),
.B1(n_552),
.B2(n_546),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_616),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_591),
.A2(n_260),
.B(n_268),
.C(n_273),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_596),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_596),
.B(n_319),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_596),
.B(n_336),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_633),
.Y(n_849)
);

INVx8_ASAP7_75t_L g850 ( 
.A(n_650),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_660),
.Y(n_851)
);

NOR3xp33_ASAP7_75t_L g852 ( 
.A(n_685),
.B(n_386),
.C(n_385),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_633),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_667),
.Y(n_854)
);

INVxp33_ASAP7_75t_L g855 ( 
.A(n_615),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_616),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_617),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_632),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_617),
.Y(n_859)
);

NAND2xp33_ASAP7_75t_L g860 ( 
.A(n_720),
.B(n_254),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_621),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_621),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_693),
.B(n_256),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_630),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_630),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_647),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_651),
.B(n_349),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_647),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_639),
.B(n_356),
.Y(n_869)
);

NAND2xp33_ASAP7_75t_L g870 ( 
.A(n_653),
.B(n_258),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_699),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_705),
.B(n_360),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_582),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_709),
.B(n_360),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_714),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_696),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_595),
.B(n_636),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_595),
.B(n_330),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_638),
.A2(n_324),
.B1(n_263),
.B2(n_375),
.Y(n_879)
);

INVxp33_ASAP7_75t_L g880 ( 
.A(n_686),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_626),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_696),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_650),
.A2(n_266),
.B1(n_274),
.B2(n_285),
.Y(n_883)
);

NAND2x1_ASAP7_75t_L g884 ( 
.A(n_632),
.B(n_260),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_792),
.A2(n_690),
.B1(n_657),
.B2(n_697),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_767),
.B(n_607),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_781),
.A2(n_638),
.B(n_670),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_846),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_793),
.Y(n_889)
);

AO21x1_ASAP7_75t_L g890 ( 
.A1(n_797),
.A2(n_698),
.B(n_585),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_745),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_743),
.A2(n_727),
.B1(n_725),
.B2(n_669),
.Y(n_892)
);

AOI21x1_ASAP7_75t_L g893 ( 
.A1(n_759),
.A2(n_585),
.B(n_582),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_855),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_742),
.A2(n_592),
.B(n_586),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_881),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_815),
.B(n_726),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_742),
.A2(n_592),
.B(n_586),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_825),
.B(n_723),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_767),
.B(n_641),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_732),
.Y(n_901)
);

NOR2x1_ASAP7_75t_L g902 ( 
.A(n_751),
.B(n_622),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_880),
.B(n_692),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_770),
.B(n_692),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_789),
.A2(n_684),
.B(n_679),
.C(n_680),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_797),
.A2(n_877),
.B1(n_875),
.B2(n_769),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_749),
.A2(n_586),
.B(n_592),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_873),
.Y(n_908)
);

NAND2xp33_ASAP7_75t_L g909 ( 
.A(n_846),
.B(n_586),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_732),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_851),
.B(n_657),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_854),
.B(n_657),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_846),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_749),
.A2(n_592),
.B(n_688),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_739),
.B(n_692),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_779),
.A2(n_688),
.B(n_593),
.Y(n_916)
);

NAND2x1p5_ASAP7_75t_L g917 ( 
.A(n_881),
.B(n_688),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_739),
.B(n_699),
.Y(n_918)
);

AOI21x1_ASAP7_75t_L g919 ( 
.A1(n_759),
.A2(n_590),
.B(n_593),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_791),
.A2(n_699),
.B1(n_701),
.B2(n_590),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_754),
.B(n_641),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_SL g922 ( 
.A(n_778),
.B(n_337),
.C(n_338),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_754),
.B(n_594),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_738),
.B(n_600),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_771),
.B(n_600),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_743),
.A2(n_598),
.B1(n_601),
.B2(n_609),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_849),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_846),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_730),
.B(n_609),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_873),
.Y(n_930)
);

AND2x2_ASAP7_75t_SL g931 ( 
.A(n_877),
.B(n_268),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_757),
.B(n_658),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_744),
.A2(n_273),
.B(n_277),
.C(n_355),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_750),
.A2(n_601),
.B(n_598),
.C(n_609),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_736),
.A2(n_301),
.B1(n_342),
.B2(n_340),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_832),
.A2(n_688),
.B(n_613),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_837),
.A2(n_300),
.B1(n_353),
.B2(n_332),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_737),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_832),
.B(n_858),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_858),
.A2(n_688),
.B(n_613),
.Y(n_940)
);

AOI21x1_ASAP7_75t_L g941 ( 
.A1(n_774),
.A2(n_612),
.B(n_626),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_872),
.B(n_612),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_775),
.A2(n_288),
.B1(n_294),
.B2(n_296),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_798),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_809),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_780),
.A2(n_613),
.B(n_612),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_734),
.A2(n_613),
.B(n_299),
.Y(n_947)
);

OAI21xp33_ASAP7_75t_L g948 ( 
.A1(n_787),
.A2(n_345),
.B(n_346),
.Y(n_948)
);

NAND2x1p5_ASAP7_75t_L g949 ( 
.A(n_815),
.B(n_613),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_837),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_SL g951 ( 
.A1(n_776),
.A2(n_293),
.B(n_379),
.C(n_373),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_819),
.B(n_675),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_837),
.A2(n_802),
.B1(n_796),
.B2(n_753),
.Y(n_953)
);

BUFx4f_ASAP7_75t_L g954 ( 
.A(n_763),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_746),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_748),
.B(n_331),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_845),
.A2(n_323),
.B(n_362),
.C(n_314),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_874),
.B(n_307),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_825),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_762),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_762),
.Y(n_961)
);

O2A1O1Ixp5_ASAP7_75t_L g962 ( 
.A1(n_802),
.A2(n_364),
.B(n_314),
.C(n_317),
.Y(n_962)
);

OR2x6_ASAP7_75t_SL g963 ( 
.A(n_853),
.B(n_358),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_775),
.A2(n_341),
.B1(n_369),
.B2(n_383),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_741),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_758),
.A2(n_364),
.B(n_333),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_845),
.A2(n_362),
.B(n_317),
.C(n_355),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_758),
.A2(n_370),
.B(n_371),
.Y(n_968)
);

AOI21x1_ASAP7_75t_L g969 ( 
.A1(n_774),
.A2(n_370),
.B(n_157),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_773),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_755),
.A2(n_367),
.B(n_361),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_810),
.B(n_716),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_753),
.A2(n_716),
.B1(n_695),
.B2(n_147),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_819),
.B(n_695),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_815),
.A2(n_132),
.B(n_184),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_815),
.B(n_280),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_752),
.A2(n_126),
.B(n_181),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_831),
.B(n_280),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_821),
.B(n_8),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_876),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_773),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_831),
.B(n_12),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_760),
.A2(n_179),
.B(n_176),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_822),
.B(n_13),
.Y(n_984)
);

NAND2xp33_ASAP7_75t_L g985 ( 
.A(n_842),
.B(n_173),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_782),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_800),
.B(n_14),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_765),
.A2(n_171),
.B(n_170),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_799),
.A2(n_161),
.B(n_159),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_740),
.A2(n_133),
.B(n_121),
.Y(n_990)
);

OR2x6_ASAP7_75t_SL g991 ( 
.A(n_735),
.B(n_15),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_747),
.A2(n_15),
.B1(n_17),
.B2(n_19),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_728),
.B(n_17),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_729),
.B(n_19),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_782),
.Y(n_995)
);

NOR2x1p5_ASAP7_75t_L g996 ( 
.A(n_763),
.B(n_21),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_733),
.A2(n_103),
.B(n_96),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_810),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_882),
.A2(n_93),
.B1(n_86),
.B2(n_81),
.Y(n_999)
);

AO22x1_ASAP7_75t_L g1000 ( 
.A1(n_838),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_1000)
);

O2A1O1Ixp5_ASAP7_75t_L g1001 ( 
.A1(n_867),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_878),
.A2(n_80),
.B1(n_27),
.B2(n_35),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_761),
.B(n_26),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_790),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_SL g1005 ( 
.A1(n_847),
.A2(n_26),
.B(n_36),
.C(n_37),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_731),
.B(n_36),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_768),
.B(n_39),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_756),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_790),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_764),
.A2(n_40),
.B(n_45),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_783),
.B(n_45),
.Y(n_1011)
);

CKINVDCx11_ASAP7_75t_R g1012 ( 
.A(n_871),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_786),
.B(n_47),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_788),
.B(n_47),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_827),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_878),
.B(n_75),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_794),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_869),
.A2(n_50),
.B(n_53),
.C(n_54),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_795),
.B(n_50),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_833),
.A2(n_53),
.B(n_55),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_834),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_766),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_808),
.B(n_59),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_836),
.A2(n_60),
.B(n_61),
.C(n_71),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_813),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_785),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_812),
.B(n_777),
.Y(n_1027)
);

OAI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_823),
.A2(n_828),
.B1(n_826),
.B2(n_835),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_860),
.A2(n_848),
.B(n_807),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_818),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_806),
.A2(n_830),
.B(n_863),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_772),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_812),
.B(n_840),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_844),
.A2(n_857),
.B(n_824),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_841),
.A2(n_844),
.B(n_857),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_801),
.Y(n_1036)
);

NOR2xp67_ASAP7_75t_L g1037 ( 
.A(n_814),
.B(n_803),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_801),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_804),
.B(n_824),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_766),
.Y(n_1040)
);

CKINVDCx10_ASAP7_75t_R g1041 ( 
.A(n_843),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_804),
.A2(n_811),
.B(n_805),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_805),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_811),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_818),
.B(n_820),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_866),
.A2(n_868),
.B(n_859),
.Y(n_1046)
);

AND2x6_ASAP7_75t_SL g1047 ( 
.A(n_816),
.B(n_817),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_856),
.A2(n_861),
.B(n_862),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_864),
.Y(n_1049)
);

AOI21x1_ASAP7_75t_L g1050 ( 
.A1(n_884),
.A2(n_865),
.B(n_829),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_816),
.B(n_817),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_870),
.A2(n_879),
.B(n_883),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_766),
.A2(n_784),
.B(n_850),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_839),
.B(n_852),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_784),
.A2(n_767),
.B(n_792),
.C(n_781),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_784),
.B(n_850),
.Y(n_1056)
);

OAI21xp33_ASAP7_75t_L g1057 ( 
.A1(n_850),
.A2(n_568),
.B(n_580),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_767),
.B(n_851),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_L g1059 ( 
.A(n_778),
.B(n_561),
.C(n_748),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_SL g1060 ( 
.A(n_1008),
.B(n_944),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_1058),
.B(n_931),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1055),
.A2(n_886),
.B(n_987),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_906),
.A2(n_953),
.B1(n_892),
.B2(n_921),
.Y(n_1064)
);

AND3x4_ASAP7_75t_L g1065 ( 
.A(n_972),
.B(n_1059),
.C(n_899),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_888),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_901),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_939),
.A2(n_1029),
.B(n_909),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_969),
.A2(n_1035),
.B(n_1050),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_941),
.A2(n_1042),
.B(n_1034),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_921),
.B(n_931),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_892),
.A2(n_915),
.B1(n_911),
.B2(n_912),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_L g1073 ( 
.A(n_1030),
.B(n_965),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_889),
.B(n_932),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_888),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_925),
.A2(n_898),
.B(n_895),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_982),
.A2(n_1045),
.B(n_922),
.C(n_915),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_889),
.B(n_952),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_907),
.A2(n_1048),
.B(n_1046),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1030),
.B(n_1028),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_890),
.A2(n_1031),
.B(n_929),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1028),
.B(n_1045),
.Y(n_1082)
);

AOI221xp5_ASAP7_75t_SL g1083 ( 
.A1(n_982),
.A2(n_933),
.B1(n_885),
.B2(n_968),
.C(n_992),
.Y(n_1083)
);

AOI211x1_ASAP7_75t_L g1084 ( 
.A1(n_922),
.A2(n_1000),
.B(n_920),
.C(n_966),
.Y(n_1084)
);

NOR2x1_ASAP7_75t_L g1085 ( 
.A(n_902),
.B(n_896),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_998),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_905),
.A2(n_926),
.B(n_934),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_918),
.B(n_1033),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_918),
.B(n_959),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_1022),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_959),
.B(n_1059),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1016),
.B(n_979),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_946),
.A2(n_940),
.B(n_936),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_914),
.A2(n_924),
.B(n_949),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_894),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_900),
.B(n_1057),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_916),
.A2(n_1010),
.B(n_1039),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_927),
.B(n_974),
.Y(n_1098)
);

AND2x6_ASAP7_75t_SL g1099 ( 
.A(n_972),
.B(n_956),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_984),
.B(n_978),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1037),
.A2(n_1052),
.B(n_962),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_950),
.A2(n_888),
.B1(n_913),
.B2(n_928),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1019),
.B(n_1023),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_891),
.B(n_904),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1038),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_888),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1019),
.B(n_1023),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_958),
.B(n_993),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_891),
.B(n_903),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_994),
.B(n_1006),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1007),
.B(n_1011),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_899),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_950),
.B(n_1054),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1013),
.B(n_1014),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_903),
.B(n_904),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_910),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_950),
.B(n_1049),
.Y(n_1117)
);

NAND2x1_ASAP7_75t_SL g1118 ( 
.A(n_1027),
.B(n_896),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_980),
.A2(n_1020),
.A3(n_956),
.B(n_961),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_942),
.A2(n_897),
.B(n_947),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_897),
.A2(n_917),
.B(n_913),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_945),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1022),
.Y(n_1123)
);

AOI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_923),
.A2(n_971),
.B(n_964),
.Y(n_1124)
);

O2A1O1Ixp5_ASAP7_75t_L g1125 ( 
.A1(n_962),
.A2(n_923),
.B(n_976),
.C(n_973),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_908),
.A2(n_930),
.B(n_989),
.Y(n_1126)
);

AO21x2_ASAP7_75t_L g1127 ( 
.A1(n_995),
.A2(n_1017),
.B(n_1036),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_913),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1044),
.A2(n_981),
.B(n_1043),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_SL g1130 ( 
.A1(n_957),
.A2(n_967),
.B(n_977),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_917),
.A2(n_913),
.B(n_928),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_928),
.A2(n_985),
.B(n_998),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1032),
.B(n_945),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_928),
.A2(n_998),
.B(n_955),
.Y(n_1134)
);

NAND2x1p5_ASAP7_75t_L g1135 ( 
.A(n_998),
.B(n_1022),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_938),
.B(n_1009),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_960),
.B(n_970),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1022),
.B(n_1056),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_1025),
.A2(n_999),
.A3(n_1004),
.B(n_986),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_990),
.A2(n_988),
.A3(n_983),
.B(n_997),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_908),
.A2(n_930),
.B(n_975),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_992),
.A2(n_1002),
.B(n_1001),
.C(n_1018),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1051),
.A2(n_1001),
.B(n_1024),
.Y(n_1143)
);

NAND3xp33_ASAP7_75t_L g1144 ( 
.A(n_948),
.B(n_937),
.C(n_935),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1021),
.A2(n_943),
.B(n_1003),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1026),
.A2(n_954),
.B(n_1040),
.C(n_1015),
.Y(n_1146)
);

AO31x2_ASAP7_75t_L g1147 ( 
.A1(n_1005),
.A2(n_951),
.A3(n_1047),
.B(n_963),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_996),
.A2(n_1012),
.B(n_954),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1041),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_991),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1058),
.B(n_767),
.Y(n_1153)
);

NAND2x1_ASAP7_75t_L g1154 ( 
.A(n_888),
.B(n_742),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1008),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1038),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_944),
.Y(n_1158)
);

NAND2x1_ASAP7_75t_L g1159 ( 
.A(n_888),
.B(n_742),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_889),
.B(n_793),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_894),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1058),
.A2(n_906),
.B1(n_1055),
.B2(n_886),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_894),
.B(n_603),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_896),
.B(n_998),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1058),
.B(n_767),
.Y(n_1166)
);

NOR2x1_ASAP7_75t_SL g1167 ( 
.A(n_888),
.B(n_913),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_894),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1058),
.B(n_767),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1058),
.A2(n_982),
.B(n_892),
.C(n_767),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1058),
.B(n_767),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_901),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_894),
.Y(n_1173)
);

AOI21xp33_ASAP7_75t_L g1174 ( 
.A1(n_921),
.A2(n_619),
.B(n_880),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1058),
.B(n_906),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_889),
.B(n_793),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1058),
.B(n_767),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_893),
.A2(n_919),
.B(n_1035),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_889),
.B(n_793),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1008),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1058),
.A2(n_982),
.B(n_892),
.C(n_767),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_890),
.A2(n_1055),
.A3(n_792),
.B(n_982),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1058),
.B(n_906),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1058),
.A2(n_906),
.B1(n_1055),
.B2(n_886),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_1012),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1058),
.B(n_767),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_894),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_SL g1189 ( 
.A1(n_982),
.A2(n_743),
.B1(n_778),
.B2(n_744),
.C(n_933),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_888),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_889),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_894),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1058),
.B(n_767),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1197)
);

OAI22x1_ASAP7_75t_L g1198 ( 
.A1(n_921),
.A2(n_701),
.B1(n_982),
.B2(n_915),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_893),
.A2(n_919),
.B(n_887),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_894),
.B(n_603),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1164),
.B(n_1200),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1166),
.B(n_1153),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_1158),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1158),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1169),
.B(n_1171),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_1186),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1178),
.B(n_1187),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1173),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1095),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1090),
.Y(n_1210)
);

BUFx10_ASAP7_75t_L g1211 ( 
.A(n_1156),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1090),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1123),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1095),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1196),
.A2(n_1182),
.B1(n_1170),
.B2(n_1107),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1061),
.B(n_1088),
.Y(n_1216)
);

CKINVDCx16_ASAP7_75t_R g1217 ( 
.A(n_1060),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1156),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1078),
.B(n_1074),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1067),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1116),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1086),
.Y(n_1222)
);

INVxp67_ASAP7_75t_SL g1223 ( 
.A(n_1193),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1068),
.A2(n_1063),
.B(n_1163),
.Y(n_1224)
);

NAND3xp33_ASAP7_75t_L g1225 ( 
.A(n_1103),
.B(n_1077),
.C(n_1174),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1061),
.A2(n_1124),
.B1(n_1071),
.B2(n_1144),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1161),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1185),
.A2(n_1120),
.B(n_1101),
.Y(n_1228)
);

NOR2xp67_ASAP7_75t_L g1229 ( 
.A(n_1181),
.B(n_1168),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1160),
.B(n_1176),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1064),
.A2(n_1100),
.B(n_1082),
.C(n_1142),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1195),
.B(n_1115),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_L g1233 ( 
.A(n_1181),
.B(n_1188),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1175),
.B(n_1184),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1096),
.B(n_1189),
.C(n_1083),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1133),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1138),
.B(n_1180),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1123),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1109),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1065),
.A2(n_1198),
.B1(n_1096),
.B2(n_1098),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1112),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1175),
.B(n_1184),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1142),
.A2(n_1080),
.B1(n_1065),
.B2(n_1092),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1066),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1186),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1193),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1138),
.B(n_1085),
.Y(n_1247)
);

INVx3_ASAP7_75t_SL g1248 ( 
.A(n_1149),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1091),
.A2(n_1111),
.B1(n_1114),
.B2(n_1110),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1172),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1108),
.A2(n_1072),
.B(n_1125),
.C(n_1104),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1138),
.B(n_1073),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1084),
.A2(n_1087),
.B1(n_1089),
.B2(n_1104),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1086),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_SL g1255 ( 
.A1(n_1113),
.A2(n_1159),
.B(n_1154),
.C(n_1146),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1066),
.Y(n_1256)
);

INVx3_ASAP7_75t_SL g1257 ( 
.A(n_1150),
.Y(n_1257)
);

OR2x4_ASAP7_75t_L g1258 ( 
.A(n_1066),
.B(n_1075),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1148),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1118),
.Y(n_1260)
);

OR2x2_ASAP7_75t_SL g1261 ( 
.A(n_1150),
.B(n_1099),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1113),
.B(n_1105),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1136),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1122),
.B(n_1117),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1146),
.A2(n_1145),
.B1(n_1148),
.B2(n_1102),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1135),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1157),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1157),
.B(n_1137),
.Y(n_1268)
);

CKINVDCx11_ASAP7_75t_R g1269 ( 
.A(n_1066),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1075),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1106),
.B(n_1191),
.Y(n_1271)
);

BUFx12f_ASAP7_75t_L g1272 ( 
.A(n_1135),
.Y(n_1272)
);

INVx3_ASAP7_75t_SL g1273 ( 
.A(n_1075),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1147),
.B(n_1119),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1165),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1147),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1075),
.A2(n_1165),
.B1(n_1129),
.B2(n_1131),
.Y(n_1277)
);

OAI21xp33_ASAP7_75t_L g1278 ( 
.A1(n_1145),
.A2(n_1143),
.B(n_1121),
.Y(n_1278)
);

OR2x6_ASAP7_75t_L g1279 ( 
.A(n_1134),
.B(n_1132),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1130),
.A2(n_1127),
.B1(n_1143),
.B2(n_1106),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1128),
.B(n_1191),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1128),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1147),
.B(n_1119),
.Y(n_1283)
);

INVx8_ASAP7_75t_L g1284 ( 
.A(n_1167),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_L g1285 ( 
.A(n_1147),
.Y(n_1285)
);

NAND3xp33_ASAP7_75t_L g1286 ( 
.A(n_1094),
.B(n_1119),
.C(n_1183),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1081),
.A2(n_1062),
.B(n_1199),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1183),
.B(n_1139),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1139),
.B(n_1141),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1183),
.B(n_1139),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1141),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1079),
.A2(n_1081),
.B(n_1076),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1183),
.B(n_1070),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1126),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1062),
.B(n_1162),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1140),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1140),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1070),
.B(n_1177),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1140),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1151),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1069),
.A2(n_1199),
.B(n_1194),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1093),
.B(n_1177),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1097),
.A2(n_1197),
.B1(n_1194),
.B2(n_1151),
.Y(n_1303)
);

OAI21xp33_ASAP7_75t_L g1304 ( 
.A1(n_1152),
.A2(n_1155),
.B(n_1190),
.Y(n_1304)
);

OR2x6_ASAP7_75t_L g1305 ( 
.A(n_1152),
.B(n_1155),
.Y(n_1305)
);

NAND2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1192),
.B(n_1197),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1179),
.B(n_1093),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1166),
.B(n_1153),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1095),
.Y(n_1309)
);

BUFx10_ASAP7_75t_L g1310 ( 
.A(n_1156),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1090),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1078),
.B(n_1074),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1061),
.B(n_1174),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1166),
.A2(n_1153),
.B1(n_1171),
.B2(n_1169),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1186),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1158),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1067),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1086),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1158),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1158),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1090),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1086),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1067),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1166),
.B(n_1153),
.Y(n_1324)
);

CKINVDCx8_ASAP7_75t_R g1325 ( 
.A(n_1156),
.Y(n_1325)
);

OR2x6_ASAP7_75t_L g1326 ( 
.A(n_1158),
.B(n_1053),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1086),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1064),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1166),
.B(n_1153),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1078),
.B(n_1074),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_1195),
.Y(n_1331)
);

NAND2x1p5_ASAP7_75t_L g1332 ( 
.A(n_1086),
.B(n_1090),
.Y(n_1332)
);

INVxp67_ASAP7_75t_SL g1333 ( 
.A(n_1095),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1164),
.B(n_1200),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1067),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1158),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1078),
.B(n_1074),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1166),
.B(n_1153),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1158),
.Y(n_1339)
);

AND2x4_ASAP7_75t_SL g1340 ( 
.A(n_1095),
.B(n_1022),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1166),
.B(n_1153),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1067),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1195),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1195),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1138),
.B(n_1022),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1061),
.A2(n_397),
.B1(n_404),
.B2(n_387),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1166),
.A2(n_1153),
.B1(n_1171),
.B2(n_1169),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1309),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1225),
.A2(n_1328),
.B(n_1231),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1284),
.Y(n_1350)
);

INVx6_ASAP7_75t_L g1351 ( 
.A(n_1272),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1315),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1202),
.A2(n_1324),
.B1(n_1329),
.B2(n_1341),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1202),
.A2(n_1324),
.B1(n_1329),
.B2(n_1341),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1328),
.A2(n_1251),
.B(n_1226),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1249),
.A2(n_1313),
.B(n_1228),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1216),
.B(n_1243),
.Y(n_1357)
);

CKINVDCx6p67_ASAP7_75t_R g1358 ( 
.A(n_1248),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1220),
.Y(n_1359)
);

INVx6_ASAP7_75t_L g1360 ( 
.A(n_1203),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1243),
.A2(n_1235),
.B1(n_1249),
.B2(n_1240),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1218),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1250),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1319),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1308),
.A2(n_1338),
.B1(n_1346),
.B2(n_1205),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1258),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1228),
.A2(n_1242),
.B(n_1234),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1215),
.A2(n_1232),
.B1(n_1216),
.B2(n_1237),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1325),
.Y(n_1369)
);

AO21x1_ASAP7_75t_L g1370 ( 
.A1(n_1215),
.A2(n_1253),
.B(n_1224),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1317),
.Y(n_1371)
);

BUFx12f_ASAP7_75t_L g1372 ( 
.A(n_1206),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1308),
.A2(n_1338),
.B1(n_1205),
.B2(n_1207),
.Y(n_1373)
);

AO21x1_ASAP7_75t_L g1374 ( 
.A1(n_1253),
.A2(n_1224),
.B(n_1234),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1284),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1230),
.B(n_1314),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1237),
.A2(n_1285),
.B1(n_1347),
.B2(n_1314),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1201),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1269),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1323),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1335),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1285),
.A2(n_1347),
.B1(n_1334),
.B2(n_1259),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_1333),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1331),
.B(n_1343),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1207),
.B(n_1219),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1342),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1217),
.A2(n_1242),
.B1(n_1239),
.B2(n_1236),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1267),
.Y(n_1388)
);

INVx4_ASAP7_75t_L g1389 ( 
.A(n_1284),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1279),
.Y(n_1390)
);

AO21x1_ASAP7_75t_SL g1391 ( 
.A1(n_1274),
.A2(n_1290),
.B(n_1265),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1331),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1279),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1239),
.B(n_1283),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1262),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1312),
.B(n_1330),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1343),
.B(n_1344),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1337),
.B(n_1236),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1262),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1263),
.Y(n_1400)
);

NOR2x1_ASAP7_75t_R g1401 ( 
.A(n_1245),
.B(n_1203),
.Y(n_1401)
);

INVx6_ASAP7_75t_L g1402 ( 
.A(n_1210),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1344),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1208),
.A2(n_1241),
.B1(n_1276),
.B2(n_1209),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1289),
.Y(n_1405)
);

AO21x1_ASAP7_75t_SL g1406 ( 
.A1(n_1290),
.A2(n_1280),
.B(n_1293),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_1244),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1289),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1282),
.Y(n_1409)
);

BUFx4f_ASAP7_75t_L g1410 ( 
.A(n_1210),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1296),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1268),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1320),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1246),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1256),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1256),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1204),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1261),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1303),
.A2(n_1307),
.B(n_1287),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1270),
.Y(n_1420)
);

INVxp67_ASAP7_75t_SL g1421 ( 
.A(n_1214),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1264),
.B(n_1252),
.Y(n_1422)
);

BUFx2_ASAP7_75t_R g1423 ( 
.A(n_1257),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1270),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1271),
.Y(n_1425)
);

BUFx2_ASAP7_75t_R g1426 ( 
.A(n_1273),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1210),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1211),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1300),
.B(n_1299),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1279),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1307),
.A2(n_1287),
.B(n_1306),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1297),
.A2(n_1252),
.B1(n_1326),
.B2(n_1247),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1326),
.A2(n_1260),
.B1(n_1229),
.B2(n_1233),
.Y(n_1433)
);

AND2x4_ASAP7_75t_SL g1434 ( 
.A(n_1211),
.B(n_1310),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1286),
.A2(n_1277),
.B(n_1278),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1326),
.A2(n_1247),
.B1(n_1345),
.B2(n_1227),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_SL g1437 ( 
.A(n_1310),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1316),
.B(n_1339),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1271),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1336),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1345),
.B(n_1281),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1340),
.A2(n_1275),
.B1(n_1266),
.B2(n_1288),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1212),
.Y(n_1443)
);

INVxp33_ASAP7_75t_L g1444 ( 
.A(n_1212),
.Y(n_1444)
);

BUFx12f_ASAP7_75t_L g1445 ( 
.A(n_1212),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1332),
.A2(n_1327),
.B1(n_1222),
.B2(n_1322),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1213),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1295),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1332),
.A2(n_1327),
.B1(n_1222),
.B2(n_1322),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1293),
.B(n_1281),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1244),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1213),
.A2(n_1238),
.B1(n_1311),
.B2(n_1321),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1305),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1298),
.A2(n_1294),
.B(n_1304),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1213),
.Y(n_1455)
);

NAND2x1p5_ASAP7_75t_L g1456 ( 
.A(n_1291),
.B(n_1302),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1305),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1305),
.Y(n_1458)
);

BUFx2_ASAP7_75t_R g1459 ( 
.A(n_1254),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1318),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1311),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1311),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1321),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1302),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1291),
.A2(n_1069),
.B(n_1292),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1255),
.B(n_1291),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1220),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1328),
.A2(n_931),
.B1(n_982),
.B2(n_922),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1220),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1292),
.A2(n_1069),
.B(n_1301),
.Y(n_1470)
);

AO21x1_ASAP7_75t_SL g1471 ( 
.A1(n_1274),
.A2(n_1242),
.B(n_1234),
.Y(n_1471)
);

OR2x6_ASAP7_75t_L g1472 ( 
.A(n_1231),
.B(n_1251),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1223),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1220),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1284),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1221),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1346),
.A2(n_567),
.B1(n_552),
.B2(n_397),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1220),
.Y(n_1478)
);

INVx5_ASAP7_75t_L g1479 ( 
.A(n_1284),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1220),
.Y(n_1480)
);

CKINVDCx14_ASAP7_75t_R g1481 ( 
.A(n_1315),
.Y(n_1481)
);

AOI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1228),
.A2(n_1292),
.B(n_1224),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1220),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1220),
.Y(n_1484)
);

AO21x1_ASAP7_75t_L g1485 ( 
.A1(n_1328),
.A2(n_1064),
.B(n_1243),
.Y(n_1485)
);

INVxp67_ASAP7_75t_SL g1486 ( 
.A(n_1383),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1468),
.A2(n_1485),
.B1(n_1361),
.B2(n_1355),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1395),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1485),
.A2(n_1472),
.B1(n_1357),
.B2(n_1349),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1464),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1448),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1448),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1395),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1473),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1390),
.B(n_1393),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1399),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1422),
.B(n_1477),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1365),
.B(n_1387),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1473),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1348),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1450),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1360),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1403),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1450),
.Y(n_1504)
);

BUFx8_ASAP7_75t_L g1505 ( 
.A(n_1437),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1360),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1392),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1453),
.Y(n_1508)
);

AO21x1_ASAP7_75t_SL g1509 ( 
.A1(n_1356),
.A2(n_1435),
.B(n_1466),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1453),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1394),
.B(n_1357),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1457),
.Y(n_1512)
);

AOI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1482),
.A2(n_1472),
.B(n_1470),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1457),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1423),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1373),
.B(n_1353),
.Y(n_1516)
);

OR2x6_ASAP7_75t_L g1517 ( 
.A(n_1390),
.B(n_1393),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1368),
.A2(n_1354),
.B1(n_1472),
.B2(n_1376),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1458),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1458),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1411),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1394),
.B(n_1376),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1411),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1367),
.B(n_1472),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1414),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1429),
.Y(n_1526)
);

INVxp67_ASAP7_75t_SL g1527 ( 
.A(n_1388),
.Y(n_1527)
);

INVx4_ASAP7_75t_SL g1528 ( 
.A(n_1437),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1471),
.B(n_1405),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1378),
.B(n_1385),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1454),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1412),
.B(n_1398),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1454),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1400),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1471),
.B(n_1405),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1479),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1408),
.B(n_1391),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1421),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1391),
.B(n_1406),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1374),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1374),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1430),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1384),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1430),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1370),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1434),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1370),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1431),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1382),
.A2(n_1377),
.B1(n_1418),
.B2(n_1432),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1465),
.A2(n_1431),
.B(n_1419),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1359),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1397),
.Y(n_1552)
);

AO21x2_ASAP7_75t_L g1553 ( 
.A1(n_1363),
.A2(n_1484),
.B(n_1483),
.Y(n_1553)
);

AOI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1433),
.A2(n_1446),
.B(n_1449),
.Y(n_1554)
);

BUFx4f_ASAP7_75t_SL g1555 ( 
.A(n_1369),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1406),
.B(n_1396),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1371),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1456),
.A2(n_1476),
.B(n_1375),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1380),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1381),
.Y(n_1560)
);

AOI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1386),
.A2(n_1467),
.B(n_1469),
.Y(n_1561)
);

INVx5_ASAP7_75t_L g1562 ( 
.A(n_1479),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1474),
.B(n_1478),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1480),
.B(n_1409),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1415),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1440),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1441),
.B(n_1362),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1416),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1441),
.B(n_1439),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1350),
.A2(n_1375),
.B(n_1475),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1420),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1462),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1424),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1460),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1350),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1404),
.B(n_1436),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1441),
.B(n_1425),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1418),
.A2(n_1437),
.B1(n_1369),
.B2(n_1358),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1366),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1434),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1366),
.A2(n_1463),
.B(n_1452),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1501),
.B(n_1504),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1559),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1552),
.B(n_1442),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1499),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1501),
.B(n_1451),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1504),
.B(n_1451),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1561),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1511),
.B(n_1379),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1559),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1517),
.B(n_1350),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1522),
.B(n_1379),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1538),
.Y(n_1593)
);

INVx4_ASAP7_75t_L g1594 ( 
.A(n_1562),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1561),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_SL g1596 ( 
.A(n_1487),
.B(n_1455),
.C(n_1362),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1553),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1553),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1524),
.B(n_1438),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1494),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1553),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1494),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_1486),
.Y(n_1603)
);

AND2x4_ASAP7_75t_SL g1604 ( 
.A(n_1536),
.B(n_1379),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1517),
.B(n_1375),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1551),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1524),
.B(n_1379),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1503),
.B(n_1461),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1522),
.B(n_1379),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1556),
.B(n_1444),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1517),
.Y(n_1611)
);

OR2x6_ASAP7_75t_L g1612 ( 
.A(n_1517),
.B(n_1389),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1498),
.A2(n_1428),
.B1(n_1481),
.B2(n_1372),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1556),
.B(n_1444),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1491),
.B(n_1461),
.Y(n_1615)
);

NOR2xp67_ASAP7_75t_L g1616 ( 
.A(n_1562),
.B(n_1475),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1491),
.B(n_1417),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1492),
.B(n_1417),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1517),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1540),
.B(n_1413),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1540),
.B(n_1413),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1495),
.Y(n_1622)
);

NAND2x1p5_ASAP7_75t_SL g1623 ( 
.A(n_1539),
.B(n_1459),
.Y(n_1623)
);

NAND4xp25_ASAP7_75t_L g1624 ( 
.A(n_1530),
.B(n_1364),
.C(n_1427),
.D(n_1389),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1500),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1550),
.A2(n_1455),
.B(n_1407),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1525),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1543),
.B(n_1447),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1546),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1516),
.B(n_1364),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1527),
.B(n_1443),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1546),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1489),
.A2(n_1428),
.B1(n_1481),
.B2(n_1372),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1541),
.B(n_1358),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1534),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1532),
.B(n_1443),
.Y(n_1636)
);

NAND4xp25_ASAP7_75t_L g1637 ( 
.A(n_1497),
.B(n_1401),
.C(n_1352),
.D(n_1447),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1580),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1549),
.A2(n_1426),
.B1(n_1351),
.B2(n_1360),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_SL g1640 ( 
.A1(n_1554),
.A2(n_1518),
.B(n_1579),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1633),
.B(n_1518),
.C(n_1566),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1599),
.B(n_1557),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1599),
.B(n_1560),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1582),
.B(n_1537),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1613),
.B(n_1528),
.Y(n_1645)
);

OAI21xp33_ASAP7_75t_L g1646 ( 
.A1(n_1596),
.A2(n_1576),
.B(n_1545),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1593),
.B(n_1496),
.Y(n_1647)
);

OAI21xp33_ASAP7_75t_L g1648 ( 
.A1(n_1639),
.A2(n_1576),
.B(n_1545),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1625),
.B(n_1496),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1589),
.B(n_1537),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1584),
.A2(n_1578),
.B1(n_1351),
.B2(n_1515),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1603),
.B(n_1508),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1630),
.B(n_1528),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1635),
.B(n_1510),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1627),
.B(n_1510),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1611),
.B(n_1529),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1619),
.B(n_1529),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1585),
.B(n_1512),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1607),
.B(n_1512),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1640),
.A2(n_1507),
.B1(n_1547),
.B2(n_1572),
.C(n_1519),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1607),
.A2(n_1509),
.B1(n_1555),
.B2(n_1569),
.Y(n_1661)
);

NOR3xp33_ASAP7_75t_L g1662 ( 
.A(n_1624),
.B(n_1554),
.C(n_1575),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1583),
.B(n_1535),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1583),
.B(n_1542),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1637),
.A2(n_1578),
.B(n_1567),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1634),
.B(n_1528),
.Y(n_1666)
);

OAI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1634),
.A2(n_1562),
.B1(n_1495),
.B2(n_1536),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1636),
.B(n_1514),
.Y(n_1668)
);

NAND3xp33_ASAP7_75t_L g1669 ( 
.A(n_1620),
.B(n_1547),
.C(n_1505),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1617),
.B(n_1514),
.Y(n_1670)
);

NAND4xp25_ASAP7_75t_SL g1671 ( 
.A(n_1592),
.B(n_1609),
.C(n_1610),
.D(n_1614),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1617),
.B(n_1519),
.Y(n_1672)
);

NAND3xp33_ASAP7_75t_L g1673 ( 
.A(n_1620),
.B(n_1544),
.C(n_1520),
.Y(n_1673)
);

NAND3xp33_ASAP7_75t_L g1674 ( 
.A(n_1621),
.B(n_1505),
.C(n_1579),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1590),
.B(n_1520),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1618),
.B(n_1631),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1590),
.B(n_1509),
.Y(n_1677)
);

OAI21xp33_ASAP7_75t_L g1678 ( 
.A1(n_1628),
.A2(n_1563),
.B(n_1564),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1618),
.B(n_1563),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1640),
.A2(n_1577),
.B1(n_1569),
.B2(n_1505),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1586),
.B(n_1564),
.Y(n_1681)
);

AOI221x1_ASAP7_75t_SL g1682 ( 
.A1(n_1608),
.A2(n_1574),
.B1(n_1571),
.B2(n_1521),
.C(n_1523),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_SL g1683 ( 
.A1(n_1604),
.A2(n_1609),
.B(n_1592),
.Y(n_1683)
);

AOI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1588),
.A2(n_1574),
.B1(n_1571),
.B2(n_1577),
.C(n_1533),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1622),
.B(n_1548),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1621),
.B(n_1581),
.C(n_1505),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1604),
.A2(n_1351),
.B1(n_1580),
.B2(n_1490),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1610),
.B(n_1580),
.Y(n_1688)
);

NAND4xp25_ASAP7_75t_L g1689 ( 
.A(n_1588),
.B(n_1573),
.C(n_1565),
.D(n_1568),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1586),
.B(n_1488),
.Y(n_1690)
);

NAND3xp33_ASAP7_75t_L g1691 ( 
.A(n_1595),
.B(n_1581),
.C(n_1526),
.Y(n_1691)
);

NOR3xp33_ASAP7_75t_L g1692 ( 
.A(n_1594),
.B(n_1575),
.C(n_1506),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1614),
.A2(n_1351),
.B1(n_1528),
.B2(n_1581),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1595),
.B(n_1581),
.C(n_1526),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1587),
.B(n_1493),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1600),
.B(n_1493),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1629),
.A2(n_1490),
.B1(n_1632),
.B2(n_1638),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1629),
.B(n_1402),
.Y(n_1698)
);

AOI221x1_ASAP7_75t_SL g1699 ( 
.A1(n_1606),
.A2(n_1523),
.B1(n_1521),
.B2(n_1531),
.C(n_1533),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1616),
.A2(n_1570),
.B(n_1558),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1644),
.B(n_1626),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1644),
.B(n_1626),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1648),
.A2(n_1646),
.B1(n_1641),
.B2(n_1645),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1664),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1663),
.B(n_1626),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1685),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1675),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1675),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1642),
.B(n_1597),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1677),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1682),
.B(n_1597),
.Y(n_1711)
);

INVxp67_ASAP7_75t_SL g1712 ( 
.A(n_1691),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1647),
.Y(n_1713)
);

NOR2x1p5_ASAP7_75t_L g1714 ( 
.A(n_1641),
.B(n_1632),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1690),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1659),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1643),
.B(n_1598),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1699),
.B(n_1598),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1700),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1692),
.B(n_1612),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1654),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1656),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1657),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1676),
.B(n_1601),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1649),
.B(n_1601),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1655),
.B(n_1658),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1650),
.B(n_1602),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1695),
.B(n_1606),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1696),
.Y(n_1729)
);

AO22x1_ASAP7_75t_L g1730 ( 
.A1(n_1662),
.A2(n_1638),
.B1(n_1562),
.B2(n_1594),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1650),
.B(n_1591),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1693),
.B(n_1591),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1693),
.B(n_1591),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1652),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1670),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1672),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1686),
.B(n_1594),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1724),
.B(n_1681),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1704),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1721),
.Y(n_1740)
);

INVxp67_ASAP7_75t_SL g1741 ( 
.A(n_1714),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1724),
.B(n_1679),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1722),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1734),
.B(n_1678),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1721),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1728),
.Y(n_1746)
);

NAND3xp33_ASAP7_75t_L g1747 ( 
.A(n_1703),
.B(n_1660),
.C(n_1648),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1726),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1704),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1728),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1726),
.B(n_1665),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1729),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1709),
.B(n_1694),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1734),
.B(n_1352),
.Y(n_1754)
);

INVxp67_ASAP7_75t_SL g1755 ( 
.A(n_1714),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1709),
.B(n_1712),
.Y(n_1756)
);

NOR2x1p5_ASAP7_75t_SL g1757 ( 
.A(n_1725),
.B(n_1513),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1722),
.B(n_1688),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1706),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1713),
.B(n_1651),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1729),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1727),
.Y(n_1762)
);

OAI33xp33_ASAP7_75t_L g1763 ( 
.A1(n_1711),
.A2(n_1678),
.A3(n_1668),
.B1(n_1689),
.B2(n_1646),
.B3(n_1673),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1713),
.B(n_1684),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1703),
.B(n_1671),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1722),
.B(n_1683),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1722),
.B(n_1591),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1707),
.Y(n_1768)
);

OAI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1719),
.A2(n_1669),
.B1(n_1674),
.B2(n_1653),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1716),
.B(n_1666),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1723),
.B(n_1605),
.Y(n_1771)
);

OR2x6_ASAP7_75t_L g1772 ( 
.A(n_1730),
.B(n_1669),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1723),
.B(n_1605),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1723),
.B(n_1605),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1707),
.Y(n_1775)
);

NAND3xp33_ASAP7_75t_L g1776 ( 
.A(n_1712),
.B(n_1661),
.C(n_1674),
.Y(n_1776)
);

AND2x4_ASAP7_75t_SL g1777 ( 
.A(n_1737),
.B(n_1605),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1706),
.Y(n_1778)
);

INVx2_ASAP7_75t_SL g1779 ( 
.A(n_1723),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1716),
.B(n_1615),
.Y(n_1780)
);

A2O1A1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1719),
.A2(n_1680),
.B(n_1623),
.C(n_1698),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1708),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1760),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1768),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1751),
.B(n_1735),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1777),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1777),
.B(n_1701),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1744),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1754),
.B(n_1763),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1756),
.B(n_1711),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1741),
.B(n_1701),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1748),
.B(n_1736),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1747),
.B(n_1736),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1755),
.B(n_1701),
.Y(n_1794)
);

NAND2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1766),
.B(n_1737),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1775),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1756),
.B(n_1718),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1739),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1782),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1752),
.Y(n_1800)
);

AND2x4_ASAP7_75t_SL g1801 ( 
.A(n_1772),
.B(n_1737),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1739),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1759),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1765),
.A2(n_1737),
.B1(n_1720),
.B2(n_1732),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1749),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1766),
.B(n_1720),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1778),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1764),
.B(n_1710),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1770),
.B(n_1710),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1746),
.B(n_1715),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1761),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1767),
.B(n_1702),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1767),
.B(n_1702),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1750),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1740),
.B(n_1715),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1771),
.B(n_1702),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1753),
.B(n_1718),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1771),
.B(n_1705),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1772),
.Y(n_1819)
);

AOI21xp33_ASAP7_75t_L g1820 ( 
.A1(n_1776),
.A2(n_1667),
.B(n_1720),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1753),
.B(n_1717),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1745),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1742),
.B(n_1717),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1769),
.B(n_1731),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1781),
.A2(n_1730),
.B(n_1720),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1772),
.Y(n_1826)
);

INVxp67_ASAP7_75t_L g1827 ( 
.A(n_1780),
.Y(n_1827)
);

NAND2x2_ASAP7_75t_L g1828 ( 
.A(n_1781),
.B(n_1743),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1784),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1812),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1784),
.Y(n_1831)
);

INVx5_ASAP7_75t_L g1832 ( 
.A(n_1819),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1789),
.B(n_1762),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1812),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1796),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1819),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1793),
.A2(n_1826),
.B1(n_1783),
.B2(n_1788),
.C(n_1820),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1796),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1785),
.B(n_1758),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1826),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1813),
.Y(n_1841)
);

INVxp67_ASAP7_75t_SL g1842 ( 
.A(n_1803),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1801),
.B(n_1772),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1797),
.B(n_1749),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1799),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1800),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1800),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1807),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1801),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1799),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1808),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1811),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1811),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1791),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1813),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1822),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1817),
.B(n_1758),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1791),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1797),
.B(n_1742),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1790),
.B(n_1738),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1816),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1822),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1790),
.B(n_1738),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1814),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1795),
.B(n_1773),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1814),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1816),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1829),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1829),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1842),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1854),
.B(n_1817),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1831),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1831),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1836),
.B(n_1824),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1837),
.A2(n_1828),
.B1(n_1825),
.B2(n_1806),
.Y(n_1875)
);

NAND2x1_ASAP7_75t_L g1876 ( 
.A(n_1843),
.B(n_1786),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1833),
.A2(n_1804),
.B1(n_1827),
.B2(n_1821),
.C(n_1794),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1849),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1832),
.B(n_1828),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1840),
.B(n_1809),
.Y(n_1880)
);

BUFx2_ASAP7_75t_SL g1881 ( 
.A(n_1832),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1848),
.B(n_1851),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1843),
.B(n_1786),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1832),
.A2(n_1806),
.B1(n_1821),
.B2(n_1795),
.Y(n_1884)
);

INVx2_ASAP7_75t_SL g1885 ( 
.A(n_1832),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1835),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1858),
.B(n_1795),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1835),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1832),
.Y(n_1889)
);

O2A1O1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1856),
.A2(n_1792),
.B(n_1794),
.C(n_1806),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1839),
.B(n_1823),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1857),
.B(n_1823),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1865),
.B(n_1787),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1838),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1866),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1838),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1885),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1883),
.B(n_1865),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1889),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1878),
.B(n_1867),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1870),
.B(n_1867),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1874),
.B(n_1830),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1883),
.B(n_1830),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1877),
.B(n_1846),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1893),
.B(n_1834),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1895),
.B(n_1847),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1880),
.B(n_1834),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1871),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1882),
.B(n_1856),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1893),
.B(n_1841),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1887),
.B(n_1841),
.Y(n_1911)
);

INVx1_ASAP7_75t_SL g1912 ( 
.A(n_1881),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1885),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1887),
.B(n_1864),
.Y(n_1914)
);

NAND2xp33_ASAP7_75t_L g1915 ( 
.A(n_1884),
.B(n_1859),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1876),
.B(n_1855),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1876),
.B(n_1855),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1871),
.Y(n_1918)
);

BUFx2_ASAP7_75t_L g1919 ( 
.A(n_1875),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1879),
.A2(n_1861),
.B1(n_1863),
.B2(n_1860),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1919),
.A2(n_1879),
.B1(n_1884),
.B2(n_1892),
.Y(n_1921)
);

BUFx2_ASAP7_75t_L g1922 ( 
.A(n_1918),
.Y(n_1922)
);

AOI222xp33_ASAP7_75t_L g1923 ( 
.A1(n_1919),
.A2(n_1891),
.B1(n_1894),
.B2(n_1896),
.C1(n_1868),
.C2(n_1888),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_SL g1924 ( 
.A(n_1912),
.B(n_1898),
.Y(n_1924)
);

AOI211xp5_ASAP7_75t_L g1925 ( 
.A1(n_1904),
.A2(n_1890),
.B(n_1886),
.C(n_1873),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1915),
.A2(n_1862),
.B(n_1864),
.Y(n_1926)
);

NAND2x1p5_ASAP7_75t_L g1927 ( 
.A(n_1912),
.B(n_1410),
.Y(n_1927)
);

AOI221xp5_ASAP7_75t_L g1928 ( 
.A1(n_1904),
.A2(n_1920),
.B1(n_1909),
.B2(n_1908),
.C(n_1900),
.Y(n_1928)
);

NOR4xp25_ASAP7_75t_SL g1929 ( 
.A(n_1908),
.B(n_1872),
.C(n_1869),
.D(n_1862),
.Y(n_1929)
);

NAND4xp75_ASAP7_75t_L g1930 ( 
.A(n_1916),
.B(n_1917),
.C(n_1899),
.D(n_1918),
.Y(n_1930)
);

AOI21xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1918),
.A2(n_1902),
.B(n_1901),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1909),
.A2(n_1906),
.B1(n_1899),
.B2(n_1907),
.C(n_1913),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1897),
.Y(n_1933)
);

NOR2x1_ASAP7_75t_L g1934 ( 
.A(n_1897),
.B(n_1845),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1924),
.B(n_1906),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1928),
.B(n_1903),
.Y(n_1936)
);

NOR4xp75_ASAP7_75t_L g1937 ( 
.A(n_1930),
.B(n_1911),
.C(n_1903),
.D(n_1898),
.Y(n_1937)
);

OA22x2_ASAP7_75t_L g1938 ( 
.A1(n_1921),
.A2(n_1917),
.B1(n_1916),
.B2(n_1914),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1922),
.B(n_1905),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1923),
.B(n_1897),
.Y(n_1940)
);

NAND3xp33_ASAP7_75t_SL g1941 ( 
.A(n_1929),
.B(n_1910),
.C(n_1905),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1933),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1934),
.Y(n_1943)
);

AND5x1_ASAP7_75t_L g1944 ( 
.A(n_1932),
.B(n_1910),
.C(n_1914),
.D(n_1861),
.E(n_1863),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1931),
.B(n_1914),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1925),
.B(n_1914),
.Y(n_1946)
);

NAND3xp33_ASAP7_75t_L g1947 ( 
.A(n_1940),
.B(n_1926),
.C(n_1850),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1939),
.Y(n_1948)
);

OAI311xp33_ASAP7_75t_L g1949 ( 
.A1(n_1936),
.A2(n_1860),
.A3(n_1859),
.B1(n_1927),
.C1(n_1844),
.Y(n_1949)
);

INVxp33_ASAP7_75t_SL g1950 ( 
.A(n_1935),
.Y(n_1950)
);

NOR3xp33_ASAP7_75t_L g1951 ( 
.A(n_1946),
.B(n_1850),
.C(n_1845),
.Y(n_1951)
);

NOR3xp33_ASAP7_75t_SL g1952 ( 
.A(n_1941),
.B(n_1853),
.C(n_1852),
.Y(n_1952)
);

NOR2x1_ASAP7_75t_L g1953 ( 
.A(n_1943),
.B(n_1852),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1948),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1947),
.B(n_1942),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1953),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1952),
.B(n_1945),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1951),
.Y(n_1958)
);

INVx2_ASAP7_75t_SL g1959 ( 
.A(n_1950),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1949),
.Y(n_1960)
);

AOI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1960),
.A2(n_1942),
.B1(n_1944),
.B2(n_1937),
.C(n_1938),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1955),
.Y(n_1962)
);

OAI21xp33_ASAP7_75t_L g1963 ( 
.A1(n_1959),
.A2(n_1853),
.B(n_1844),
.Y(n_1963)
);

NOR3x2_ASAP7_75t_L g1964 ( 
.A(n_1957),
.B(n_1528),
.C(n_1445),
.Y(n_1964)
);

NAND5xp2_ASAP7_75t_L g1965 ( 
.A(n_1954),
.B(n_1787),
.C(n_1733),
.D(n_1732),
.E(n_1818),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_1956),
.Y(n_1966)
);

NAND2x1p5_ASAP7_75t_L g1967 ( 
.A(n_1966),
.B(n_1958),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1963),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_SL g1969 ( 
.A1(n_1962),
.A2(n_1957),
.B1(n_1445),
.B2(n_1779),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1964),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1967),
.A2(n_1961),
.B1(n_1798),
.B2(n_1805),
.Y(n_1971)
);

XNOR2x1_ASAP7_75t_L g1972 ( 
.A(n_1971),
.B(n_1968),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1972),
.A2(n_1969),
.B(n_1970),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1972),
.Y(n_1974)
);

NAND3xp33_ASAP7_75t_L g1975 ( 
.A(n_1973),
.B(n_1965),
.C(n_1802),
.Y(n_1975)
);

OAI21x1_ASAP7_75t_SL g1976 ( 
.A1(n_1974),
.A2(n_1802),
.B(n_1798),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1975),
.B(n_1805),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1976),
.B(n_1815),
.Y(n_1978)
);

AOI222xp33_ASAP7_75t_L g1979 ( 
.A1(n_1977),
.A2(n_1810),
.B1(n_1757),
.B2(n_1818),
.C1(n_1743),
.C2(n_1779),
.Y(n_1979)
);

AOI222xp33_ASAP7_75t_L g1980 ( 
.A1(n_1979),
.A2(n_1978),
.B1(n_1757),
.B2(n_1410),
.C1(n_1774),
.C2(n_1773),
.Y(n_1980)
);

OAI221xp5_ASAP7_75t_L g1981 ( 
.A1(n_1980),
.A2(n_1410),
.B1(n_1402),
.B2(n_1443),
.C(n_1502),
.Y(n_1981)
);

AOI211xp5_ASAP7_75t_L g1982 ( 
.A1(n_1981),
.A2(n_1687),
.B(n_1536),
.C(n_1697),
.Y(n_1982)
);


endmodule