module real_aes_8441_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_0), .B(n_111), .C(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g122 ( .A(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g535 ( .A(n_1), .Y(n_535) );
INVx1_ASAP7_75t_L g156 ( .A(n_2), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_3), .A2(n_38), .B1(n_181), .B2(n_481), .Y(n_504) );
AOI21xp33_ASAP7_75t_L g188 ( .A1(n_4), .A2(n_172), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_5), .B(n_170), .Y(n_547) );
AND2x6_ASAP7_75t_L g149 ( .A(n_6), .B(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_7), .A2(n_259), .B(n_260), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_8), .B(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_8), .B(n_39), .Y(n_123) );
INVx1_ASAP7_75t_L g194 ( .A(n_9), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_10), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g141 ( .A(n_11), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_12), .B(n_162), .Y(n_490) );
INVx1_ASAP7_75t_L g265 ( .A(n_13), .Y(n_265) );
INVx1_ASAP7_75t_L g529 ( .A(n_14), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_15), .B(n_137), .Y(n_518) );
AO32x2_ASAP7_75t_L g502 ( .A1(n_16), .A2(n_136), .A3(n_170), .B1(n_483), .B2(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_17), .B(n_181), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_18), .B(n_177), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_19), .B(n_137), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_20), .A2(n_49), .B1(n_181), .B2(n_481), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_21), .B(n_172), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_22), .A2(n_98), .B1(n_737), .B2(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_22), .Y(n_738) );
AOI22xp33_ASAP7_75t_SL g482 ( .A1(n_23), .A2(n_75), .B1(n_162), .B2(n_181), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_24), .B(n_181), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_25), .B(n_184), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_26), .A2(n_263), .B(n_264), .C(n_266), .Y(n_262) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_27), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_28), .B(n_167), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_29), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_30), .B(n_117), .Y(n_443) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_31), .A2(n_87), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_31), .Y(n_127) );
INVx1_ASAP7_75t_L g209 ( .A(n_32), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_33), .B(n_167), .Y(n_474) );
INVx2_ASAP7_75t_L g147 ( .A(n_34), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_35), .B(n_181), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_36), .B(n_167), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_37), .A2(n_149), .B(n_152), .C(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g109 ( .A(n_39), .Y(n_109) );
INVx1_ASAP7_75t_L g207 ( .A(n_40), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_41), .B(n_160), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_42), .B(n_181), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_43), .A2(n_85), .B1(n_229), .B2(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_44), .B(n_181), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_45), .B(n_181), .Y(n_530) );
CKINVDCx16_ASAP7_75t_R g210 ( .A(n_46), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_47), .B(n_534), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_48), .B(n_172), .Y(n_253) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_50), .A2(n_60), .B1(n_162), .B2(n_181), .Y(n_522) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_51), .A2(n_735), .B1(n_736), .B2(n_739), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_51), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_52), .A2(n_152), .B1(n_162), .B2(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_53), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_54), .B(n_181), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g143 ( .A(n_55), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_56), .B(n_181), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_57), .A2(n_180), .B(n_192), .C(n_193), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_58), .Y(n_242) );
INVx1_ASAP7_75t_L g190 ( .A(n_59), .Y(n_190) );
INVx1_ASAP7_75t_L g150 ( .A(n_61), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_62), .B(n_181), .Y(n_536) );
INVx1_ASAP7_75t_L g140 ( .A(n_63), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_64), .Y(n_446) );
AO32x2_ASAP7_75t_L g478 ( .A1(n_65), .A2(n_170), .A3(n_245), .B1(n_479), .B2(n_483), .Y(n_478) );
INVx1_ASAP7_75t_L g554 ( .A(n_66), .Y(n_554) );
INVx1_ASAP7_75t_L g469 ( .A(n_67), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_68), .A2(n_125), .B1(n_441), .B2(n_442), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_68), .Y(n_441) );
A2O1A1Ixp33_ASAP7_75t_SL g176 ( .A1(n_69), .A2(n_177), .B(n_178), .C(n_180), .Y(n_176) );
INVxp67_ASAP7_75t_L g179 ( .A(n_70), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_71), .B(n_162), .Y(n_470) );
INVx1_ASAP7_75t_L g114 ( .A(n_72), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_73), .Y(n_212) );
INVx1_ASAP7_75t_L g235 ( .A(n_74), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_76), .A2(n_149), .B(n_152), .C(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_77), .B(n_481), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_78), .B(n_162), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_79), .B(n_157), .Y(n_225) );
INVx2_ASAP7_75t_L g138 ( .A(n_80), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_81), .B(n_177), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_82), .B(n_162), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_83), .A2(n_149), .B(n_152), .C(n_155), .Y(n_151) );
INVx2_ASAP7_75t_L g111 ( .A(n_84), .Y(n_111) );
OR2x2_ASAP7_75t_L g119 ( .A(n_84), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g452 ( .A(n_84), .B(n_121), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_86), .A2(n_102), .B1(n_162), .B2(n_163), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_87), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_88), .B(n_167), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_89), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_90), .A2(n_149), .B(n_152), .C(n_248), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_91), .Y(n_255) );
INVx1_ASAP7_75t_L g175 ( .A(n_92), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_93), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_94), .B(n_157), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_95), .A2(n_104), .B1(n_115), .B2(n_745), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_96), .B(n_162), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_97), .B(n_170), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_98), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_100), .A2(n_172), .B(n_173), .Y(n_171) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_101), .A2(n_449), .B1(n_733), .B2(n_734), .C1(n_740), .C2(n_743), .Y(n_448) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g746 ( .A(n_107), .Y(n_746) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
OR2x2_ASAP7_75t_L g456 ( .A(n_111), .B(n_121), .Y(n_456) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_111), .B(n_120), .Y(n_742) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AO21x1_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_444), .B(n_447), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_124), .B(n_443), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g442 ( .A(n_125), .Y(n_442) );
XNOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
INVx1_ASAP7_75t_L g453 ( .A(n_129), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_129), .A2(n_454), .B1(n_458), .B2(n_744), .Y(n_743) );
NAND2x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_357), .Y(n_129) );
NOR5xp2_ASAP7_75t_L g130 ( .A(n_131), .B(n_280), .C(n_312), .D(n_327), .E(n_344), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_196), .B(n_217), .C(n_268), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_168), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_133), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_133), .B(n_332), .Y(n_395) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_134), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_134), .B(n_214), .Y(n_281) );
AND2x2_ASAP7_75t_L g322 ( .A(n_134), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_134), .B(n_291), .Y(n_326) );
OR2x2_ASAP7_75t_L g363 ( .A(n_134), .B(n_202), .Y(n_363) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g201 ( .A(n_135), .B(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g271 ( .A(n_135), .Y(n_271) );
OR2x2_ASAP7_75t_L g434 ( .A(n_135), .B(n_274), .Y(n_434) );
AO21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_142), .B(n_164), .Y(n_135) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_136), .A2(n_203), .B(n_211), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_136), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g230 ( .A(n_136), .Y(n_230) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_137), .Y(n_170) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_138), .B(n_139), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_151), .Y(n_142) );
OAI22xp33_ASAP7_75t_L g203 ( .A1(n_144), .A2(n_182), .B1(n_204), .B2(n_210), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_144), .A2(n_235), .B(n_236), .Y(n_234) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
AND2x4_ASAP7_75t_L g172 ( .A(n_145), .B(n_149), .Y(n_172) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g534 ( .A(n_146), .Y(n_534) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
INVx1_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx3_ASAP7_75t_L g158 ( .A(n_148), .Y(n_158) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_148), .Y(n_160) );
INVx1_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_148), .Y(n_206) );
INVx4_ASAP7_75t_SL g182 ( .A(n_149), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_149), .A2(n_468), .B(n_471), .Y(n_467) );
BUFx3_ASAP7_75t_L g483 ( .A(n_149), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_149), .A2(n_488), .B(n_492), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_149), .A2(n_528), .B(n_532), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_149), .A2(n_541), .B(n_544), .Y(n_540) );
INVx5_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
BUFx3_ASAP7_75t_L g229 ( .A(n_153), .Y(n_229) );
INVx1_ASAP7_75t_L g481 ( .A(n_153), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_159), .C(n_161), .Y(n_155) );
O2A1O1Ixp5_ASAP7_75t_SL g468 ( .A1(n_157), .A2(n_180), .B(n_469), .C(n_470), .Y(n_468) );
INVx2_ASAP7_75t_L g505 ( .A(n_157), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_157), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_157), .A2(n_551), .B(n_552), .Y(n_550) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_158), .B(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_158), .B(n_194), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g479 ( .A1(n_158), .A2(n_160), .B1(n_480), .B2(n_482), .Y(n_479) );
INVx2_ASAP7_75t_L g192 ( .A(n_160), .Y(n_192) );
INVx4_ASAP7_75t_L g251 ( .A(n_160), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_160), .A2(n_504), .B1(n_505), .B2(n_506), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_160), .A2(n_505), .B1(n_521), .B2(n_522), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_161), .A2(n_529), .B(n_530), .C(n_531), .Y(n_528) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_166), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_166), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g245 ( .A(n_167), .Y(n_245) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_167), .A2(n_258), .B(n_267), .Y(n_257) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_167), .A2(n_467), .B(n_474), .Y(n_466) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_167), .A2(n_487), .B(n_495), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_168), .A2(n_337), .B1(n_338), .B2(n_341), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_168), .B(n_271), .Y(n_420) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_186), .Y(n_168) );
AND2x2_ASAP7_75t_L g216 ( .A(n_169), .B(n_202), .Y(n_216) );
AND2x2_ASAP7_75t_L g273 ( .A(n_169), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g278 ( .A(n_169), .Y(n_278) );
INVx3_ASAP7_75t_L g291 ( .A(n_169), .Y(n_291) );
OR2x2_ASAP7_75t_L g311 ( .A(n_169), .B(n_274), .Y(n_311) );
AND2x2_ASAP7_75t_L g330 ( .A(n_169), .B(n_187), .Y(n_330) );
BUFx2_ASAP7_75t_L g362 ( .A(n_169), .Y(n_362) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_183), .Y(n_169) );
INVx4_ASAP7_75t_L g185 ( .A(n_170), .Y(n_185) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_170), .A2(n_540), .B(n_547), .Y(n_539) );
BUFx2_ASAP7_75t_L g259 ( .A(n_172), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_182), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_174), .A2(n_182), .B(n_190), .C(n_191), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_174), .A2(n_182), .B(n_261), .C(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g491 ( .A(n_177), .Y(n_491) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_181), .Y(n_252) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_184), .A2(n_188), .B(n_195), .Y(n_187) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_SL g231 ( .A(n_185), .B(n_232), .Y(n_231) );
NAND3xp33_ASAP7_75t_L g519 ( .A(n_185), .B(n_483), .C(n_520), .Y(n_519) );
AO21x1_ASAP7_75t_L g609 ( .A1(n_185), .A2(n_520), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g277 ( .A(n_186), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
BUFx2_ASAP7_75t_L g200 ( .A(n_187), .Y(n_200) );
INVx2_ASAP7_75t_L g215 ( .A(n_187), .Y(n_215) );
OR2x2_ASAP7_75t_L g293 ( .A(n_187), .B(n_274), .Y(n_293) );
AND2x2_ASAP7_75t_L g323 ( .A(n_187), .B(n_202), .Y(n_323) );
AND2x2_ASAP7_75t_L g340 ( .A(n_187), .B(n_271), .Y(n_340) );
AND2x2_ASAP7_75t_L g380 ( .A(n_187), .B(n_291), .Y(n_380) );
AND2x2_ASAP7_75t_SL g416 ( .A(n_187), .B(n_216), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_192), .A2(n_493), .B(n_494), .Y(n_492) );
O2A1O1Ixp5_ASAP7_75t_L g553 ( .A1(n_192), .A2(n_533), .B(n_554), .C(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp33_ASAP7_75t_SL g197 ( .A(n_198), .B(n_213), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_201), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_199), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
OAI21xp33_ASAP7_75t_L g354 ( .A1(n_200), .A2(n_216), .B(n_355), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_200), .B(n_202), .Y(n_410) );
AND2x2_ASAP7_75t_L g346 ( .A(n_201), .B(n_347), .Y(n_346) );
INVx3_ASAP7_75t_L g274 ( .A(n_202), .Y(n_274) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_202), .Y(n_372) );
OAI22xp5_ASAP7_75t_SL g205 ( .A1(n_206), .A2(n_207), .B1(n_208), .B2(n_209), .Y(n_205) );
INVx2_ASAP7_75t_L g208 ( .A(n_206), .Y(n_208) );
INVx4_ASAP7_75t_L g263 ( .A(n_206), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_213), .B(n_271), .Y(n_439) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_214), .A2(n_382), .B1(n_383), .B2(n_388), .Y(n_381) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
AND2x2_ASAP7_75t_L g272 ( .A(n_215), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g310 ( .A(n_215), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_SL g347 ( .A(n_215), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_216), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g401 ( .A(n_216), .Y(n_401) );
CKINVDCx16_ASAP7_75t_R g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_243), .Y(n_218) );
INVx4_ASAP7_75t_L g287 ( .A(n_219), .Y(n_287) );
AND2x2_ASAP7_75t_L g365 ( .A(n_219), .B(n_332), .Y(n_365) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_233), .Y(n_219) );
INVx3_ASAP7_75t_L g284 ( .A(n_220), .Y(n_284) );
AND2x2_ASAP7_75t_L g298 ( .A(n_220), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g302 ( .A(n_220), .Y(n_302) );
INVx2_ASAP7_75t_L g316 ( .A(n_220), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_220), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g373 ( .A(n_220), .B(n_368), .Y(n_373) );
AND2x2_ASAP7_75t_L g438 ( .A(n_220), .B(n_408), .Y(n_438) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_231), .Y(n_220) );
AOI21xp5_ASAP7_75t_SL g221 ( .A1(n_222), .A2(n_223), .B(n_230), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_227), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_227), .A2(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g266 ( .A(n_229), .Y(n_266) );
INVx1_ASAP7_75t_L g240 ( .A(n_230), .Y(n_240) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_230), .A2(n_527), .B(n_537), .Y(n_526) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_230), .A2(n_549), .B(n_556), .Y(n_548) );
AND2x2_ASAP7_75t_L g279 ( .A(n_233), .B(n_257), .Y(n_279) );
INVx2_ASAP7_75t_L g299 ( .A(n_233), .Y(n_299) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_240), .B(n_241), .Y(n_233) );
INVx1_ASAP7_75t_L g304 ( .A(n_243), .Y(n_304) );
AND2x2_ASAP7_75t_L g350 ( .A(n_243), .B(n_298), .Y(n_350) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_256), .Y(n_243) );
INVx2_ASAP7_75t_L g289 ( .A(n_244), .Y(n_289) );
INVx1_ASAP7_75t_L g297 ( .A(n_244), .Y(n_297) );
AND2x2_ASAP7_75t_L g315 ( .A(n_244), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_244), .B(n_299), .Y(n_353) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_254), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_253), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B(n_252), .Y(n_248) );
AND2x2_ASAP7_75t_L g332 ( .A(n_256), .B(n_289), .Y(n_332) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g285 ( .A(n_257), .Y(n_285) );
AND2x2_ASAP7_75t_L g368 ( .A(n_257), .B(n_299), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_263), .B(n_265), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_263), .A2(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g531 ( .A(n_263), .Y(n_531) );
OAI21xp5_ASAP7_75t_SL g268 ( .A1(n_269), .A2(n_275), .B(n_279), .Y(n_268) );
INVx1_ASAP7_75t_SL g313 ( .A(n_269), .Y(n_313) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_270), .B(n_277), .Y(n_370) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g319 ( .A(n_271), .B(n_274), .Y(n_319) );
AND2x2_ASAP7_75t_L g348 ( .A(n_271), .B(n_292), .Y(n_348) );
OR2x2_ASAP7_75t_L g351 ( .A(n_271), .B(n_311), .Y(n_351) );
AOI222xp33_ASAP7_75t_L g415 ( .A1(n_272), .A2(n_364), .B1(n_416), .B2(n_417), .C1(n_419), .C2(n_421), .Y(n_415) );
BUFx2_ASAP7_75t_L g329 ( .A(n_274), .Y(n_329) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g318 ( .A(n_277), .B(n_319), .Y(n_318) );
INVx3_ASAP7_75t_SL g335 ( .A(n_277), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_277), .B(n_329), .Y(n_389) );
AND2x2_ASAP7_75t_L g324 ( .A(n_279), .B(n_284), .Y(n_324) );
INVx1_ASAP7_75t_L g343 ( .A(n_279), .Y(n_343) );
OAI221xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_282), .B1(n_286), .B2(n_290), .C(n_294), .Y(n_280) );
OR2x2_ASAP7_75t_L g352 ( .A(n_282), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g337 ( .A(n_284), .B(n_307), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_284), .B(n_297), .Y(n_377) );
AND2x2_ASAP7_75t_L g382 ( .A(n_284), .B(n_332), .Y(n_382) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_284), .Y(n_392) );
NAND2x1_ASAP7_75t_SL g403 ( .A(n_284), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g288 ( .A(n_285), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g308 ( .A(n_285), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_285), .B(n_303), .Y(n_334) );
INVx1_ASAP7_75t_L g400 ( .A(n_285), .Y(n_400) );
INVx1_ASAP7_75t_L g375 ( .A(n_286), .Y(n_375) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g387 ( .A(n_287), .Y(n_387) );
NOR2xp67_ASAP7_75t_L g399 ( .A(n_287), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g404 ( .A(n_288), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_288), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g307 ( .A(n_289), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_289), .B(n_299), .Y(n_320) );
INVx1_ASAP7_75t_L g386 ( .A(n_289), .Y(n_386) );
INVx1_ASAP7_75t_L g407 ( .A(n_290), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI21xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_300), .B(n_309), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
AND2x2_ASAP7_75t_L g440 ( .A(n_296), .B(n_373), .Y(n_440) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g408 ( .A(n_297), .B(n_368), .Y(n_408) );
AOI32xp33_ASAP7_75t_L g321 ( .A1(n_298), .A2(n_304), .A3(n_322), .B1(n_324), .B2(n_325), .Y(n_321) );
AOI322xp5_ASAP7_75t_L g423 ( .A1(n_298), .A2(n_330), .A3(n_413), .B1(n_424), .B2(n_425), .C1(n_426), .C2(n_428), .Y(n_423) );
INVx2_ASAP7_75t_L g303 ( .A(n_299), .Y(n_303) );
INVx1_ASAP7_75t_L g413 ( .A(n_299), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .B1(n_305), .B2(n_306), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_301), .B(n_307), .Y(n_356) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_302), .B(n_368), .Y(n_418) );
INVx1_ASAP7_75t_L g305 ( .A(n_303), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_303), .B(n_332), .Y(n_422) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_311), .B(n_406), .Y(n_405) );
OAI221xp5_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_314), .B1(n_317), .B2(n_320), .C(n_321), .Y(n_312) );
OR2x2_ASAP7_75t_L g333 ( .A(n_314), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g342 ( .A(n_314), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g367 ( .A(n_315), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g371 ( .A(n_325), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI221xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_331), .B1(n_333), .B2(n_335), .C(n_336), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_329), .A2(n_360), .B1(n_364), .B2(n_365), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_330), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g435 ( .A(n_330), .Y(n_435) );
INVx1_ASAP7_75t_L g429 ( .A(n_332), .Y(n_429) );
INVx1_ASAP7_75t_SL g364 ( .A(n_333), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_335), .B(n_363), .Y(n_425) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_340), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g406 ( .A(n_340), .Y(n_406) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
OAI221xp5_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_349), .B1(n_351), .B2(n_352), .C(n_354), .Y(n_344) );
NOR2xp33_ASAP7_75t_SL g345 ( .A(n_346), .B(n_348), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_346), .A2(n_364), .B1(n_410), .B2(n_411), .Y(n_409) );
CKINVDCx14_ASAP7_75t_R g349 ( .A(n_350), .Y(n_349) );
OAI21xp33_ASAP7_75t_L g428 ( .A1(n_351), .A2(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR3xp33_ASAP7_75t_SL g357 ( .A(n_358), .B(n_390), .C(n_414), .Y(n_357) );
NAND4xp25_ASAP7_75t_L g358 ( .A(n_359), .B(n_366), .C(n_374), .D(n_381), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g437 ( .A(n_362), .Y(n_437) );
INVx3_ASAP7_75t_SL g431 ( .A(n_363), .Y(n_431) );
OR2x2_ASAP7_75t_L g436 ( .A(n_363), .B(n_437), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B1(n_371), .B2(n_373), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_368), .B(n_386), .Y(n_427) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI21xp5_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_376), .B(n_378), .Y(n_374) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI211xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_393), .B(n_396), .C(n_409), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g424 ( .A(n_395), .Y(n_424) );
AOI222xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_401), .B1(n_402), .B2(n_405), .C1(n_407), .C2(n_408), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND4xp25_ASAP7_75t_SL g433 ( .A(n_406), .B(n_434), .C(n_435), .D(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND3xp33_ASAP7_75t_SL g414 ( .A(n_415), .B(n_423), .C(n_432), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_438), .B1(n_439), .B2(n_440), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g447 ( .A1(n_443), .A2(n_444), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_453), .B1(n_454), .B2(n_457), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g744 ( .A(n_451), .Y(n_744) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_654), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_603), .C(n_645), .Y(n_459) );
AOI211xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_512), .B(n_557), .C(n_579), .Y(n_460) );
OAI211xp5_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_475), .B(n_496), .C(n_507), .Y(n_461) );
INVxp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_463), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g666 ( .A(n_463), .B(n_583), .Y(n_666) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g568 ( .A(n_464), .B(n_499), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_464), .B(n_486), .Y(n_685) );
INVx1_ASAP7_75t_L g703 ( .A(n_464), .Y(n_703) );
AND2x2_ASAP7_75t_L g712 ( .A(n_464), .B(n_600), .Y(n_712) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g595 ( .A(n_465), .B(n_486), .Y(n_595) );
AND2x2_ASAP7_75t_L g653 ( .A(n_465), .B(n_600), .Y(n_653) );
INVx1_ASAP7_75t_L g697 ( .A(n_465), .Y(n_697) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g574 ( .A(n_466), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g582 ( .A(n_466), .Y(n_582) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_466), .Y(n_622) );
INVxp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_484), .Y(n_476) );
AND2x2_ASAP7_75t_L g561 ( .A(n_477), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g594 ( .A(n_477), .Y(n_594) );
OR2x2_ASAP7_75t_L g720 ( .A(n_477), .B(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_477), .B(n_486), .Y(n_724) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g499 ( .A(n_478), .Y(n_499) );
INVx1_ASAP7_75t_L g510 ( .A(n_478), .Y(n_510) );
AND2x2_ASAP7_75t_L g583 ( .A(n_478), .B(n_501), .Y(n_583) );
AND2x2_ASAP7_75t_L g623 ( .A(n_478), .B(n_502), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_483), .A2(n_550), .B(n_553), .Y(n_549) );
INVxp67_ASAP7_75t_L g665 ( .A(n_484), .Y(n_665) );
AND2x4_ASAP7_75t_L g690 ( .A(n_484), .B(n_583), .Y(n_690) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_SL g581 ( .A(n_485), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g500 ( .A(n_486), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g569 ( .A(n_486), .B(n_502), .Y(n_569) );
INVx1_ASAP7_75t_L g575 ( .A(n_486), .Y(n_575) );
INVx2_ASAP7_75t_L g601 ( .A(n_486), .Y(n_601) );
AND2x2_ASAP7_75t_L g617 ( .A(n_486), .B(n_618), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_491), .Y(n_488) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_497), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g572 ( .A(n_499), .Y(n_572) );
AND2x2_ASAP7_75t_L g680 ( .A(n_499), .B(n_501), .Y(n_680) );
AND2x2_ASAP7_75t_L g597 ( .A(n_500), .B(n_582), .Y(n_597) );
AND2x2_ASAP7_75t_L g696 ( .A(n_500), .B(n_697), .Y(n_696) );
NOR2xp67_ASAP7_75t_L g618 ( .A(n_501), .B(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g721 ( .A(n_501), .B(n_582), .Y(n_721) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g511 ( .A(n_502), .Y(n_511) );
AND2x2_ASAP7_75t_L g600 ( .A(n_502), .B(n_601), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_505), .A2(n_533), .B(n_535), .C(n_536), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_505), .A2(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
AND2x2_ASAP7_75t_L g646 ( .A(n_509), .B(n_581), .Y(n_646) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_510), .B(n_582), .Y(n_631) );
INVx2_ASAP7_75t_L g630 ( .A(n_511), .Y(n_630) );
OAI222xp33_ASAP7_75t_L g634 ( .A1(n_511), .A2(n_574), .B1(n_635), .B2(n_637), .C1(n_638), .C2(n_641), .Y(n_634) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_523), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g559 ( .A(n_516), .Y(n_559) );
OR2x2_ASAP7_75t_L g670 ( .A(n_516), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g592 ( .A(n_517), .Y(n_592) );
NOR2x1_ASAP7_75t_L g643 ( .A(n_517), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g649 ( .A(n_517), .B(n_563), .Y(n_649) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g610 ( .A(n_518), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_523), .A2(n_613), .B1(n_652), .B2(n_653), .Y(n_651) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_538), .Y(n_523) );
INVx3_ASAP7_75t_L g585 ( .A(n_524), .Y(n_585) );
OR2x2_ASAP7_75t_L g718 ( .A(n_524), .B(n_594), .Y(n_718) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g591 ( .A(n_525), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g607 ( .A(n_525), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g615 ( .A(n_525), .B(n_563), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_525), .B(n_539), .Y(n_671) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g562 ( .A(n_526), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g566 ( .A(n_526), .B(n_539), .Y(n_566) );
AND2x2_ASAP7_75t_L g642 ( .A(n_526), .B(n_589), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_526), .B(n_548), .Y(n_682) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_538), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g598 ( .A(n_538), .B(n_559), .Y(n_598) );
AND2x2_ASAP7_75t_L g602 ( .A(n_538), .B(n_592), .Y(n_602) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_548), .Y(n_538) );
INVx3_ASAP7_75t_L g563 ( .A(n_539), .Y(n_563) );
AND2x2_ASAP7_75t_L g588 ( .A(n_539), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g723 ( .A(n_539), .B(n_706), .Y(n_723) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_548), .Y(n_577) );
INVx2_ASAP7_75t_L g589 ( .A(n_548), .Y(n_589) );
AND2x2_ASAP7_75t_L g633 ( .A(n_548), .B(n_609), .Y(n_633) );
INVx1_ASAP7_75t_L g676 ( .A(n_548), .Y(n_676) );
OR2x2_ASAP7_75t_L g707 ( .A(n_548), .B(n_609), .Y(n_707) );
AND2x2_ASAP7_75t_L g727 ( .A(n_548), .B(n_563), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_560), .B(n_564), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g565 ( .A(n_559), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_559), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g684 ( .A(n_561), .Y(n_684) );
INVx2_ASAP7_75t_SL g578 ( .A(n_562), .Y(n_578) );
AND2x2_ASAP7_75t_L g698 ( .A(n_562), .B(n_592), .Y(n_698) );
INVx2_ASAP7_75t_L g644 ( .A(n_563), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_563), .B(n_676), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_567), .B1(n_570), .B2(n_576), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_566), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g732 ( .A(n_566), .Y(n_732) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g657 ( .A(n_568), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_568), .B(n_600), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_569), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g673 ( .A(n_569), .B(n_622), .Y(n_673) );
INVx2_ASAP7_75t_L g729 ( .A(n_569), .Y(n_729) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AND2x2_ASAP7_75t_L g599 ( .A(n_572), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_572), .B(n_617), .Y(n_650) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_574), .B(n_594), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g711 ( .A(n_577), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_SL g661 ( .A1(n_578), .A2(n_662), .B(n_664), .C(n_667), .Y(n_661) );
OR2x2_ASAP7_75t_L g688 ( .A(n_578), .B(n_592), .Y(n_688) );
OAI221xp5_ASAP7_75t_SL g579 ( .A1(n_580), .A2(n_584), .B1(n_586), .B2(n_593), .C(n_596), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_581), .B(n_583), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_581), .B(n_630), .Y(n_637) );
AND2x2_ASAP7_75t_L g679 ( .A(n_581), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g715 ( .A(n_581), .Y(n_715) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_582), .Y(n_606) );
INVx1_ASAP7_75t_L g619 ( .A(n_582), .Y(n_619) );
NOR2xp67_ASAP7_75t_L g639 ( .A(n_585), .B(n_640), .Y(n_639) );
INVxp67_ASAP7_75t_L g693 ( .A(n_585), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_585), .B(n_633), .Y(n_709) );
INVx2_ASAP7_75t_L g695 ( .A(n_586), .Y(n_695) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g636 ( .A(n_588), .B(n_607), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_588), .A2(n_604), .B(n_646), .C(n_647), .Y(n_645) );
AND2x2_ASAP7_75t_L g614 ( .A(n_589), .B(n_609), .Y(n_614) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_593), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
OR2x2_ASAP7_75t_L g662 ( .A(n_594), .B(n_663), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_599), .B2(n_602), .Y(n_596) );
INVx1_ASAP7_75t_L g716 ( .A(n_598), .Y(n_716) );
INVx1_ASAP7_75t_L g663 ( .A(n_600), .Y(n_663) );
INVx1_ASAP7_75t_L g714 ( .A(n_602), .Y(n_714) );
AOI211xp5_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_607), .B(n_611), .C(n_634), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g626 ( .A(n_606), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g677 ( .A(n_607), .Y(n_677) );
AND2x2_ASAP7_75t_L g726 ( .A(n_607), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_616), .B(n_624), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx2_ASAP7_75t_L g640 ( .A(n_614), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_614), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g632 ( .A(n_615), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g708 ( .A(n_615), .Y(n_708) );
OAI32xp33_ASAP7_75t_L g719 ( .A1(n_615), .A2(n_667), .A3(n_674), .B1(n_715), .B2(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_SL g616 ( .A(n_617), .B(n_620), .Y(n_616) );
INVx1_ASAP7_75t_SL g687 ( .A(n_617), .Y(n_687) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g627 ( .A(n_623), .Y(n_627) );
OAI21xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_628), .B(n_632), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g699 ( .A1(n_626), .A2(n_674), .B1(n_700), .B2(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_630), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g667 ( .A(n_633), .Y(n_667) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g660 ( .A(n_644), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_650), .B(n_651), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_653), .A2(n_695), .B1(n_696), .B2(n_698), .C(n_699), .Y(n_694) );
NAND5xp2_ASAP7_75t_L g654 ( .A(n_655), .B(n_678), .C(n_694), .D(n_704), .E(n_722), .Y(n_654) );
AOI211xp5_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_658), .B(n_661), .C(n_668), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g725 ( .A(n_662), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_672), .B2(n_674), .Y(n_668) );
INVx1_ASAP7_75t_SL g701 ( .A(n_671), .Y(n_701) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI322xp33_ASAP7_75t_L g683 ( .A1(n_674), .A2(n_684), .A3(n_685), .B1(n_686), .B2(n_687), .C1(n_688), .C2(n_689), .Y(n_683) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g686 ( .A(n_676), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_676), .B(n_701), .Y(n_700) );
AOI211xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_681), .B(n_683), .C(n_691), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_687), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_713) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g730 ( .A(n_697), .Y(n_730) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_712), .B1(n_713), .B2(n_717), .C(n_719), .Y(n_704) );
OAI211xp5_ASAP7_75t_SL g705 ( .A1(n_706), .A2(n_708), .B(n_709), .C(n_710), .Y(n_705) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g731 ( .A(n_707), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_725), .B2(n_726), .C(n_728), .Y(n_722) );
AOI21xp33_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_730), .B(n_731), .Y(n_728) );
CKINVDCx16_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
endmodule