module fake_jpeg_26249_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_22),
.B(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_68),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_71),
.B(n_57),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_63),
.B1(n_60),
.B2(n_46),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_79),
.B1(n_1),
.B2(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_60),
.B1(n_63),
.B2(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_55),
.B1(n_61),
.B2(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_80),
.A2(n_82),
.B1(n_86),
.B2(n_49),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_54),
.B1(n_58),
.B2(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_53),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_50),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_93),
.B1(n_98),
.B2(n_102),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_91),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_49),
.B(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_94),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_50),
.B1(n_64),
.B2(n_3),
.Y(n_93)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_83),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_97),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_73),
.B1(n_79),
.B2(n_3),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_103),
.B1(n_2),
.B2(n_4),
.Y(n_112)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_38),
.B1(n_35),
.B2(n_33),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_112),
.B1(n_100),
.B2(n_89),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_113),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_96),
.B(n_90),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_117),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_118),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_102),
.B1(n_95),
.B2(n_87),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_120),
.B1(n_107),
.B2(n_110),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_104),
.A2(n_97),
.B(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_107),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_124),
.B(n_128),
.C(n_5),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_112),
.B1(n_111),
.B2(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_100),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_130),
.C(n_27),
.Y(n_132)
);

AOI221xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_131),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_108),
.B1(n_32),
.B2(n_28),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_26),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_132),
.A2(n_133),
.B1(n_128),
.B2(n_7),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_25),
.C(n_24),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);

OAI322xp33_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_127),
.A3(n_129),
.B1(n_128),
.B2(n_20),
.C1(n_18),
.C2(n_16),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_133),
.C(n_134),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_138),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_138),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_137),
.B1(n_8),
.B2(n_9),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_6),
.C(n_8),
.Y(n_144)
);

OAI321xp33_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_10),
.B(n_11),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_12),
.Y(n_148)
);


endmodule