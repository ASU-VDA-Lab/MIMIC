module fake_jpeg_19242_n_166 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_29),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_25),
.B1(n_28),
.B2(n_20),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_19),
.B1(n_16),
.B2(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_38),
.B1(n_25),
.B2(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_24),
.A2(n_16),
.B1(n_19),
.B2(n_18),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_19),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_29),
.C(n_30),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_44),
.B1(n_39),
.B2(n_33),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_11),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_11),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_54),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_26),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

AOI32xp33_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_41),
.A3(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_59),
.Y(n_78)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_62),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_20),
.C(n_41),
.Y(n_62)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_72),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_39),
.B1(n_46),
.B2(n_56),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_23),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_27),
.C(n_30),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_69),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_26),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_86),
.B1(n_37),
.B2(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_26),
.B(n_23),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_26),
.B(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_67),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_67),
.B1(n_72),
.B2(n_59),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_100),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_95),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_62),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_101),
.B1(n_80),
.B2(n_77),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_78),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_37),
.B1(n_33),
.B2(n_51),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_76),
.B(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_17),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_103),
.B(n_105),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_85),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_115),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_88),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_81),
.B1(n_79),
.B2(n_33),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_100),
.B(n_102),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_118),
.B1(n_87),
.B2(n_18),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_95),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_130),
.C(n_131),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_98),
.B1(n_94),
.B2(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_129),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_101),
.B1(n_106),
.B2(n_97),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_118),
.B1(n_42),
.B2(n_27),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_110),
.B1(n_111),
.B2(n_120),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_114),
.C(n_108),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_30),
.C(n_27),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_139),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_137),
.B1(n_15),
.B2(n_14),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_17),
.B(n_1),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_131),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_141),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_130),
.C(n_124),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_122),
.C(n_126),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_143),
.C(n_138),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_15),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_151),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_144),
.A2(n_135),
.B(n_10),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_148),
.B(n_149),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_15),
.C(n_14),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_140),
.B(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_152),
.B(n_14),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_9),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_157),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_0),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_155),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_159),
.A2(n_160),
.B(n_153),
.C(n_158),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.C(n_4),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_4),
.B(n_5),
.Y(n_164)
);

OAI221xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_6),
.Y(n_166)
);


endmodule