module fake_jpeg_14584_n_162 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_162);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_5),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_SL g62 ( 
.A(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_3),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_3),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_15),
.Y(n_58)
);

CKINVDCx9p33_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_17),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_49),
.B1(n_30),
.B2(n_13),
.Y(n_57)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_24),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_6),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_7),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_31),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_17),
.A2(n_8),
.B1(n_11),
.B2(n_29),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_50),
.A2(n_17),
.B1(n_29),
.B2(n_16),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_61),
.B1(n_65),
.B2(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_22),
.B1(n_26),
.B2(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_58),
.B(n_74),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_29),
.B1(n_21),
.B2(n_31),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_21),
.B1(n_13),
.B2(n_18),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_14),
.Y(n_67)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_19),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_33),
.A2(n_19),
.B1(n_22),
.B2(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_93),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_49),
.B(n_46),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_72),
.B(n_63),
.Y(n_102)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_71),
.B1(n_62),
.B2(n_69),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_87),
.B(n_95),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_91),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_20),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_11),
.B1(n_52),
.B2(n_60),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_68),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_62),
.A2(n_60),
.B1(n_54),
.B2(n_77),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_64),
.B1(n_91),
.B2(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_79),
.B(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_59),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_114),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_64),
.B1(n_70),
.B2(n_69),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_87),
.B1(n_94),
.B2(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_89),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_105),
.C(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_117),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_85),
.B1(n_95),
.B2(n_86),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_130),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_101),
.B1(n_127),
.B2(n_129),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_124),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_115),
.B(n_113),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_108),
.B(n_111),
.C(n_116),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_110),
.C(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_126),
.B(n_129),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_103),
.C(n_109),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_121),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_117),
.C(n_108),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_124),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_137),
.Y(n_145)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_123),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_140),
.A2(n_142),
.B1(n_128),
.B2(n_137),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_134),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_125),
.C(n_126),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_146),
.C(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_148),
.A2(n_142),
.B1(n_140),
.B2(n_144),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_152),
.Y(n_157)
);

AND2x4_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_140),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_154),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_143),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.C(n_156),
.Y(n_161)
);

OAI211xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_153),
.B(n_156),
.C(n_140),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);


endmodule