module fake_jpeg_15931_n_275 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_275);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_31),
.Y(n_60)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_17),
.B1(n_25),
.B2(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_59),
.B1(n_26),
.B2(n_25),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_54),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx2_ASAP7_75t_SL g75 ( 
.A(n_55),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_25),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_24),
.B1(n_15),
.B2(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_27),
.C(n_29),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_46),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_73),
.B1(n_19),
.B2(n_16),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_46),
.B1(n_42),
.B2(n_39),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_74),
.B1(n_65),
.B2(n_55),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_17),
.B1(n_19),
.B2(n_16),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_42),
.B1(n_34),
.B2(n_33),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_55),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_80),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_42),
.B1(n_34),
.B2(n_35),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_84),
.B1(n_66),
.B2(n_45),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_52),
.B1(n_55),
.B2(n_66),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_34),
.C(n_13),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_95),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_56),
.B1(n_54),
.B2(n_52),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_107),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_61),
.B1(n_57),
.B2(n_69),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_99),
.B1(n_105),
.B2(n_91),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_57),
.B1(n_69),
.B2(n_67),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_97),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_61),
.B1(n_67),
.B2(n_60),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_103),
.B(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_106),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_68),
.B(n_23),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_13),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_82),
.B(n_81),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_112),
.B(n_98),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_81),
.B(n_80),
.Y(n_112)
);

AO21x2_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_84),
.B(n_74),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_64),
.B(n_50),
.C(n_40),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_119),
.B1(n_95),
.B2(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_15),
.A3(n_24),
.B1(n_19),
.B2(n_16),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_22),
.B(n_14),
.C(n_20),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_35),
.B1(n_30),
.B2(n_88),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_85),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_29),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_27),
.C(n_29),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_128),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_27),
.C(n_29),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_23),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_132),
.A2(n_138),
.B(n_147),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_148),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_140),
.B1(n_152),
.B2(n_131),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_106),
.B1(n_49),
.B2(n_45),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_139),
.B1(n_143),
.B2(n_145),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_108),
.C(n_13),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_138),
.C(n_129),
.Y(n_159)
);

OAI22x1_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_108),
.B1(n_14),
.B2(n_48),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_35),
.B1(n_30),
.B2(n_64),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_15),
.B1(n_24),
.B2(n_49),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_30),
.B1(n_35),
.B2(n_22),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_22),
.Y(n_146)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_45),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_22),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_123),
.B1(n_112),
.B2(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_14),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_121),
.C(n_116),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_162),
.C(n_164),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_171),
.B1(n_177),
.B2(n_20),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_124),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_160),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_122),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_111),
.C(n_125),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_126),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_145),
.B1(n_139),
.B2(n_143),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_132),
.B(n_125),
.CI(n_118),
.CON(n_166),
.SN(n_166)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_11),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_12),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_124),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_176),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_120),
.B(n_48),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NOR4xp25_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_120),
.C(n_48),
.D(n_28),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_120),
.B(n_1),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_162),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_180),
.C(n_181),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_153),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_136),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_156),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_183),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_171),
.B1(n_169),
.B2(n_161),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_163),
.A2(n_145),
.B1(n_30),
.B2(n_64),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_186),
.B1(n_198),
.B2(n_177),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_50),
.C(n_28),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_197),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_173),
.B(n_12),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_50),
.C(n_28),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_155),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_203),
.C(n_209),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_155),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_204),
.B(n_205),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_165),
.B1(n_161),
.B2(n_170),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_180),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_178),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_10),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_210),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_184),
.B(n_194),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_195),
.B(n_1),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_213),
.C(n_201),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_218),
.C(n_219),
.Y(n_234)
);

HAxp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_181),
.CON(n_222),
.SN(n_222)
);

OAI21x1_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_204),
.B(n_202),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_2),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_190),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_229),
.B(n_230),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_197),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_213),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_234),
.C(n_240),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_222),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_241),
.B(n_226),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_0),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_20),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_238),
.B(n_224),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_225),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_3),
.B(n_4),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_20),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_21),
.C(n_20),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_248),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_244),
.A2(n_245),
.B1(n_242),
.B2(n_236),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_223),
.B(n_228),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_217),
.C(n_223),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_249),
.B(n_251),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_20),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_256),
.Y(n_261)
);

AO21x1_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_260),
.B(n_21),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_250),
.B(n_231),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_3),
.B(n_4),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_5),
.B(n_6),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_21),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_248),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_21),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_265),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_6),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_253),
.B(n_260),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_7),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_7),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_268),
.B1(n_7),
.B2(n_8),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_7),
.C(n_8),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_274),
.B(n_8),
.Y(n_275)
);


endmodule