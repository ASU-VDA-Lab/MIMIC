module fake_jpeg_30277_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx8_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_0),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_64),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_2),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_20),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_42),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_55),
.B1(n_46),
.B2(n_52),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_69),
.B1(n_78),
.B2(n_64),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_72),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_52),
.B1(n_49),
.B2(n_48),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_54),
.C(n_53),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_75),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NOR4xp25_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_26),
.C(n_41),
.D(n_40),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_44),
.B(n_4),
.C(n_5),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_56),
.B1(n_51),
.B2(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_43),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_89),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_93),
.B1(n_8),
.B2(n_9),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_6),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_19),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_57),
.B(n_5),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_6),
.B(n_7),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_3),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_21),
.B1(n_37),
.B2(n_35),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_11),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_68),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_102),
.C(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_105),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_10),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_70),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_80),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_90),
.B1(n_89),
.B2(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_112),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_96),
.C(n_98),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_8),
.B(n_9),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_SL g120 ( 
.A(n_115),
.B(n_116),
.C(n_117),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_39),
.B(n_25),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_119),
.A3(n_99),
.B1(n_27),
.B2(n_29),
.C1(n_31),
.C2(n_32),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_121),
.A2(n_116),
.B(n_33),
.C(n_34),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_110),
.C(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_126),
.C(n_127),
.Y(n_128)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_112),
.C(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_116),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_123),
.A3(n_120),
.B1(n_114),
.B2(n_113),
.C1(n_108),
.C2(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_23),
.B(n_120),
.Y(n_133)
);


endmodule