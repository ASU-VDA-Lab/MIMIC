module real_jpeg_24876_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_18),
.B1(n_19),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_1),
.A2(n_22),
.B1(n_27),
.B2(n_32),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_32),
.B1(n_55),
.B2(n_56),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_35),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_4),
.A2(n_37),
.B(n_53),
.C(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_4),
.B(n_22),
.C(n_25),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_18),
.B1(n_19),
.B2(n_54),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_4),
.A2(n_40),
.B(n_46),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_5),
.A2(n_22),
.B1(n_27),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_6),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_20),
.B1(n_22),
.B2(n_27),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_22),
.B1(n_27),
.B2(n_45),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_8),
.A2(n_18),
.B1(n_19),
.B2(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_10),
.A2(n_41),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_77),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_76),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_50),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_15),
.B(n_50),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_33),
.C(n_39),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_16),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_21),
.B(n_28),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_18),
.A2(n_19),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g53 ( 
.A1(n_18),
.A2(n_38),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_54),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_29),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_29),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_31),
.B(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_35),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_38),
.B1(n_55),
.B2(n_56),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_39),
.B(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B(n_46),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_49),
.Y(n_62)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_48),
.B(n_54),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_62),
.B(n_91),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_63),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B(n_62),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_103),
.B(n_108),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_93),
.B(n_102),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_89),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_89),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_98),
.B(n_101),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_107),
.Y(n_108)
);


endmodule