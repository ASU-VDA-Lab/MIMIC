module fake_jpeg_12886_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_7),
.B(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_4),
.B(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_44),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_6),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_45),
.B(n_50),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_49),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_29),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_51),
.B(n_54),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_52),
.B(n_55),
.Y(n_127)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_60),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_5),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_58),
.Y(n_102)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_27),
.B(n_5),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_66),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_27),
.A2(n_8),
.B(n_12),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_69),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_14),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_38),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_14),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_83),
.B(n_11),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_37),
.B1(n_32),
.B2(n_22),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_87),
.A2(n_95),
.B1(n_114),
.B2(n_118),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_49),
.A2(n_24),
.B1(n_42),
.B2(n_37),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_97),
.B(n_101),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_28),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_26),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_103),
.B(n_113),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_48),
.A2(n_16),
.B1(n_24),
.B2(n_36),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_116),
.B1(n_128),
.B2(n_110),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_62),
.A2(n_32),
.B1(n_22),
.B2(n_36),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_125),
.B1(n_134),
.B2(n_121),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_44),
.B(n_37),
.C(n_42),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_121),
.C(n_66),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_46),
.B(n_43),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_65),
.A2(n_42),
.B1(n_37),
.B2(n_40),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_61),
.A2(n_16),
.B1(n_36),
.B2(n_32),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_75),
.A2(n_22),
.B1(n_16),
.B2(n_41),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_46),
.B(n_41),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_119),
.B(n_129),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_40),
.B1(n_34),
.B2(n_35),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_72),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_76),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_4),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_77),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_54),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_135)
);

FAx1_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_98),
.CI(n_126),
.CON(n_154),
.SN(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_11),
.Y(n_138)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_138),
.B(n_143),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_140),
.B(n_157),
.Y(n_198)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_175),
.B1(n_137),
.B2(n_141),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_80),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_82),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_144),
.B(n_162),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_161),
.Y(n_185)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_87),
.B1(n_112),
.B2(n_117),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_159),
.B1(n_146),
.B2(n_172),
.Y(n_183)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_SL g149 ( 
.A(n_102),
.B(n_66),
.C(n_1),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_154),
.C(n_156),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_1),
.B1(n_3),
.B2(n_100),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_167),
.Y(n_188)
);

OA22x2_ASAP7_75t_SL g151 ( 
.A1(n_135),
.A2(n_124),
.B1(n_109),
.B2(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_153),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_SL g200 ( 
.A(n_154),
.B(n_166),
.C(n_173),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_117),
.C(n_123),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_166),
.C(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_112),
.A2(n_106),
.B1(n_123),
.B2(n_85),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_124),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_171),
.Y(n_187)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_86),
.B(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_102),
.B(n_122),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_164),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_94),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_165),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_122),
.C(n_131),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_100),
.A2(n_131),
.B1(n_107),
.B2(n_92),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_169),
.Y(n_211)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_88),
.B(n_120),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_88),
.B(n_85),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_90),
.B(n_104),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_104),
.A2(n_106),
.B1(n_132),
.B2(n_99),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_90),
.B(n_115),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_107),
.B(n_89),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_168),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_209),
.B1(n_213),
.B2(n_211),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_183),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_154),
.B1(n_151),
.B2(n_145),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_182),
.B1(n_201),
.B2(n_185),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_155),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_201),
.C(n_204),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_176),
.B(n_178),
.C(n_171),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_182),
.B(n_212),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_197),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_212),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_170),
.C(n_165),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_148),
.A2(n_153),
.B1(n_152),
.B2(n_161),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_154),
.A2(n_144),
.B(n_151),
.C(n_145),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

AOI221xp5_ASAP7_75t_L g248 ( 
.A1(n_218),
.A2(n_189),
.B1(n_225),
.B2(n_219),
.C(n_220),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_181),
.B1(n_187),
.B2(n_195),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_214),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_200),
.A2(n_202),
.B1(n_206),
.B2(n_199),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_226),
.B1(n_233),
.B2(n_234),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_185),
.A2(n_202),
.B1(n_199),
.B2(n_204),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_206),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_230),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_191),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_188),
.A2(n_190),
.B1(n_198),
.B2(n_208),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_188),
.A2(n_190),
.B1(n_198),
.B2(n_208),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_211),
.B1(n_213),
.B2(n_189),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_238),
.B1(n_236),
.B2(n_226),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_237),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_207),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_184),
.B(n_203),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_239),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_189),
.C(n_203),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g273 ( 
.A1(n_247),
.A2(n_248),
.B(n_252),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_218),
.C(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_251),
.C(n_257),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_231),
.CI(n_216),
.CON(n_250),
.SN(n_250)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_250),
.B(n_227),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_218),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_260),
.B1(n_244),
.B2(n_257),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_234),
.C(n_233),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_228),
.A2(n_215),
.B1(n_223),
.B2(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_266),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_268),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_243),
.A2(n_221),
.B1(n_217),
.B2(n_215),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_224),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_232),
.C(n_237),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_246),
.C(n_255),
.Y(n_289)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_274),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_277),
.B(n_247),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_256),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_260),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_276),
.Y(n_285)
);

OA22x2_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_241),
.B1(n_245),
.B2(n_250),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_277),
.B(n_265),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_249),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_286),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_244),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_276),
.C(n_246),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_293),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_275),
.B1(n_278),
.B2(n_285),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_296),
.B1(n_287),
.B2(n_269),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_270),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_255),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_297),
.Y(n_304)
);

AOI31xp67_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_276),
.A3(n_250),
.B(n_272),
.Y(n_295)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_268),
.B1(n_262),
.B2(n_276),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_299),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_276),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_289),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_305),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_296),
.Y(n_302)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_280),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_302),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_292),
.C(n_294),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_309),
.C(n_305),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_297),
.C(n_291),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_281),
.B(n_274),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_300),
.B(n_303),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_287),
.B1(n_281),
.B2(n_279),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_315),
.A2(n_316),
.B1(n_266),
.B2(n_271),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_295),
.C(n_261),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_320),
.B(n_318),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_267),
.B1(n_245),
.B2(n_263),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_317),
.C(n_312),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_307),
.Y(n_323)
);


endmodule