module fake_ariane_1134_n_2188 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2188);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2188;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_204),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_63),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_85),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_87),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_134),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_63),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_111),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_10),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_1),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_56),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_56),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_88),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_139),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_40),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_138),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_12),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_77),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_195),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_27),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_5),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_98),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_6),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_85),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_93),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_17),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_172),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_106),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_144),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_99),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_142),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_215),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_105),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_118),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_168),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_68),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_129),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_149),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_57),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_153),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_184),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_69),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_179),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_132),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_120),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_114),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_86),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_15),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_191),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_54),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_58),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_81),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_102),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_218),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_42),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_113),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_94),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_147),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_35),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_131),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_154),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_17),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_90),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_32),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_100),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_217),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_7),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_70),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_21),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_45),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_77),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_35),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_31),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_206),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_171),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_159),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_74),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_62),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_44),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_76),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_32),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_156),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_127),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_194),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_20),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_182),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_23),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_41),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_203),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_181),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_167),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_158),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_42),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_33),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_123),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_8),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_9),
.Y(n_320)
);

BUFx8_ASAP7_75t_SL g321 ( 
.A(n_69),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_163),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_200),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_59),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_47),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_13),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_13),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_8),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_96),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_116),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_50),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_178),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_122),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_82),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_173),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_101),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_5),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_188),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_82),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_207),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_70),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_36),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_78),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_19),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_46),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_219),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_146),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_196),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_216),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_212),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_125),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_38),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_110),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_79),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_183),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_137),
.Y(n_356)
);

BUFx10_ASAP7_75t_L g357 ( 
.A(n_34),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_27),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_43),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_119),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_193),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_40),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_73),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_136),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_202),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_3),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_65),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_164),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_91),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_75),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_31),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_26),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_41),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_155),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_198),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_79),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_9),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_185),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_76),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_145),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_24),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_21),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_10),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_117),
.Y(n_384)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_52),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_135),
.Y(n_386)
);

BUFx10_ASAP7_75t_L g387 ( 
.A(n_89),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_133),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_33),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_126),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_4),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_150),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_161),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_44),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_115),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_62),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_18),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_143),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_84),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_50),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_52),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_86),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_103),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_60),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_175),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_75),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_109),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_151),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_199),
.Y(n_409)
);

BUFx10_ASAP7_75t_L g410 ( 
.A(n_104),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_112),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_64),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_130),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_83),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_18),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_148),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_81),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_162),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_46),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_7),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_160),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_30),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_38),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_28),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_30),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_0),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_210),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_97),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_1),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_80),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_141),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_95),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_6),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_366),
.B(n_0),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_264),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_366),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_321),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_275),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_367),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_323),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_385),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_261),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_385),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_385),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_385),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_287),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_261),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_252),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_385),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_407),
.B(n_2),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_335),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_385),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_366),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_353),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_364),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_403),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_366),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_223),
.B(n_2),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_311),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_223),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_325),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_396),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_427),
.B(n_3),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_325),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_337),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_331),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_396),
.Y(n_471)
);

INVxp33_ASAP7_75t_SL g472 ( 
.A(n_316),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_224),
.B(n_11),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_236),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_224),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_399),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_225),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_225),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_337),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_221),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_230),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_229),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_230),
.B(n_11),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_238),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_231),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_228),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_238),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_233),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_237),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_239),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_334),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_252),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_249),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_240),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_242),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_228),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_249),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_251),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_251),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_243),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_259),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_352),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_415),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g504 ( 
.A(n_342),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_259),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_354),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_263),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_245),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g509 ( 
.A(n_246),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_263),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_267),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_342),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_267),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_248),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_271),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_272),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_271),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_359),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_279),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_273),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_383),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_288),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_288),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_274),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_279),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_286),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_288),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_286),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_282),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_305),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_344),
.B(n_12),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_291),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_305),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_288),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_313),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_336),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_292),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_336),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_313),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_293),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_294),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_336),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_376),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_329),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_296),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_300),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_301),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_461),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_461),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_464),
.B(n_475),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_435),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_435),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_442),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_503),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_467),
.B(n_415),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_503),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_442),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_464),
.B(n_475),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_477),
.B(n_329),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_443),
.Y(n_560)
);

BUFx8_ASAP7_75t_L g561 ( 
.A(n_479),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_457),
.B(n_244),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_477),
.B(n_330),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_463),
.B(n_304),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_452),
.B(n_415),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_466),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_443),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_470),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_445),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_457),
.B(n_244),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_445),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_446),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_478),
.B(n_376),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_446),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_447),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_447),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_451),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_451),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_454),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_454),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_456),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_471),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_478),
.B(n_412),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_456),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_449),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_457),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_481),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_481),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_484),
.B(n_412),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_480),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_531),
.B(n_344),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_484),
.Y(n_592)
);

CKINVDCx6p67_ASAP7_75t_R g593 ( 
.A(n_450),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_487),
.B(n_415),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_487),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_493),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_493),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_497),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_497),
.B(n_330),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_498),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_498),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_499),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_474),
.B(n_303),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g604 ( 
.A1(n_491),
.A2(n_414),
.B1(n_226),
.B2(n_258),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_499),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_501),
.B(n_303),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_501),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_505),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_505),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_474),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_507),
.Y(n_611)
);

NOR2x1_ASAP7_75t_L g612 ( 
.A(n_474),
.B(n_236),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_507),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_510),
.B(n_373),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_510),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_511),
.B(n_333),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_511),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_513),
.B(n_373),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_513),
.B(n_336),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_515),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_515),
.B(n_333),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_517),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_517),
.Y(n_623)
);

NOR2x1_ASAP7_75t_L g624 ( 
.A(n_519),
.B(n_347),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_519),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_525),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_525),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_453),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_526),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_526),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_528),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_528),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_530),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_530),
.B(n_356),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_533),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_533),
.B(n_415),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_476),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_SL g638 ( 
.A(n_590),
.B(n_482),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_550),
.B(n_465),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_586),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_590),
.B(n_450),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_586),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_586),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_L g644 ( 
.A(n_551),
.B(n_485),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_587),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_587),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_610),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_619),
.B(n_610),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_585),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_586),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_566),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_587),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_619),
.B(n_468),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_587),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_586),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_586),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_587),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_619),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_590),
.B(n_492),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_587),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_634),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_586),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_610),
.B(n_509),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_587),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_596),
.Y(n_665)
);

AND2x6_ASAP7_75t_L g666 ( 
.A(n_550),
.B(n_340),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_550),
.B(n_437),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_576),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g669 ( 
.A(n_568),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_591),
.A2(n_492),
.B1(n_472),
.B2(n_489),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_L g671 ( 
.A(n_551),
.B(n_488),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_596),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_582),
.B(n_490),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_596),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_576),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_582),
.B(n_494),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_576),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_591),
.A2(n_500),
.B1(n_508),
.B2(n_495),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_596),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_566),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_565),
.B(n_516),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_591),
.A2(n_524),
.B1(n_529),
.B2(n_520),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_565),
.B(n_532),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_L g684 ( 
.A1(n_591),
.A2(n_593),
.B1(n_444),
.B2(n_531),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_578),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_588),
.B(n_537),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_597),
.B(n_588),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_596),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_591),
.A2(n_462),
.B1(n_483),
.B2(n_473),
.Y(n_689)
);

NOR2x1p5_ASAP7_75t_L g690 ( 
.A(n_593),
.B(n_438),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_596),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_591),
.A2(n_539),
.B1(n_544),
.B2(n_535),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_592),
.B(n_540),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_592),
.B(n_541),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_573),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_578),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_552),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_595),
.B(n_545),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_596),
.Y(n_699)
);

AND2x2_ASAP7_75t_SL g700 ( 
.A(n_636),
.B(n_340),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_573),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_568),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_606),
.B(n_469),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_603),
.B(n_504),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_578),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_585),
.B(n_448),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_579),
.Y(n_707)
);

AND2x2_ASAP7_75t_SL g708 ( 
.A(n_594),
.B(n_350),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_558),
.B(n_547),
.C(n_546),
.Y(n_709)
);

BUFx4f_ASAP7_75t_L g710 ( 
.A(n_617),
.Y(n_710)
);

OR2x6_ASAP7_75t_L g711 ( 
.A(n_603),
.B(n_479),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_552),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_579),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_553),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_606),
.B(n_512),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_617),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_579),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_597),
.B(n_535),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_L g719 ( 
.A(n_551),
.B(n_350),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_597),
.B(n_539),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_595),
.B(n_436),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_573),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_617),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_617),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_597),
.B(n_544),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_583),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_553),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_597),
.B(n_439),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_558),
.B(n_441),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_551),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_617),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_603),
.B(n_543),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_593),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_580),
.Y(n_734)
);

CKINVDCx6p67_ASAP7_75t_R g735 ( 
.A(n_628),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_617),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_580),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_580),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_598),
.B(n_455),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_SL g740 ( 
.A(n_598),
.B(n_522),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_601),
.B(n_458),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_601),
.B(n_440),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_617),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_603),
.A2(n_523),
.B1(n_534),
.B2(n_527),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_584),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_548),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_605),
.B(n_459),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_584),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_548),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_628),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_605),
.B(n_536),
.Y(n_751)
);

BUFx6f_ASAP7_75t_SL g752 ( 
.A(n_603),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_606),
.B(n_486),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_584),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_614),
.A2(n_624),
.B1(n_555),
.B2(n_612),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_549),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_549),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_604),
.B(n_496),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_551),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_561),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_551),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_607),
.B(n_434),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_551),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_636),
.B(n_365),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_600),
.Y(n_765)
);

INVx5_ASAP7_75t_L g766 ( 
.A(n_634),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_560),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_600),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_604),
.B(n_514),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_560),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_600),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_602),
.Y(n_772)
);

AND3x2_ASAP7_75t_L g773 ( 
.A(n_637),
.B(n_258),
.C(n_248),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_560),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_607),
.B(n_434),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_602),
.Y(n_776)
);

AND2x6_ASAP7_75t_L g777 ( 
.A(n_636),
.B(n_365),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_560),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_560),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_618),
.B(n_222),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_602),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_611),
.Y(n_782)
);

OR2x6_ASAP7_75t_L g783 ( 
.A(n_618),
.B(n_614),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_560),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_608),
.B(n_538),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_560),
.Y(n_786)
);

AOI21x1_ASAP7_75t_L g787 ( 
.A1(n_557),
.A2(n_390),
.B(n_380),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_618),
.B(n_583),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_614),
.A2(n_542),
.B1(n_270),
.B2(n_276),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_571),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_571),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_571),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_658),
.B(n_608),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_780),
.B(n_583),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_700),
.B(n_557),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_658),
.B(n_609),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_668),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_686),
.B(n_693),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_668),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_694),
.B(n_609),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_706),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_698),
.B(n_653),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_700),
.B(n_567),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_675),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_746),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_785),
.B(n_518),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_675),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_706),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_746),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_700),
.A2(n_561),
.B1(n_624),
.B2(n_555),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_653),
.B(n_615),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_786),
.B(n_567),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_677),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_677),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_685),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_685),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_696),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_696),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_680),
.B(n_460),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_750),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_786),
.B(n_569),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_729),
.B(n_561),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_666),
.A2(n_561),
.B1(n_637),
.B2(n_614),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_721),
.B(n_561),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_786),
.B(n_569),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_742),
.B(n_502),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_653),
.B(n_615),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_765),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_705),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_765),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_681),
.B(n_506),
.Y(n_831)
);

OR2x6_ASAP7_75t_L g832 ( 
.A(n_783),
.B(n_614),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_705),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_689),
.A2(n_623),
.B1(n_626),
.B2(n_622),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_780),
.B(n_622),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_711),
.Y(n_836)
);

INVxp33_ASAP7_75t_L g837 ( 
.A(n_750),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_647),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_L g839 ( 
.A(n_666),
.B(n_571),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_697),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_667),
.A2(n_577),
.B(n_581),
.C(n_572),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_695),
.B(n_623),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_666),
.A2(n_612),
.B1(n_636),
.B2(n_627),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_695),
.B(n_701),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_749),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_663),
.B(n_627),
.C(n_626),
.Y(n_846)
);

BUFx4_ASAP7_75t_L g847 ( 
.A(n_735),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_783),
.B(n_589),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_683),
.B(n_521),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_786),
.B(n_572),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_701),
.B(n_630),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_722),
.B(n_630),
.Y(n_852)
);

INVxp67_ASAP7_75t_SL g853 ( 
.A(n_647),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_728),
.B(n_631),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_756),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_756),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_739),
.B(n_631),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_722),
.B(n_633),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_726),
.B(n_633),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_726),
.B(n_635),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_757),
.Y(n_861)
);

BUFx8_ASAP7_75t_L g862 ( 
.A(n_752),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_666),
.A2(n_636),
.B1(n_635),
.B2(n_589),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_757),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_786),
.B(n_577),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_697),
.A2(n_563),
.B1(n_599),
.B2(n_559),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_666),
.A2(n_589),
.B1(n_613),
.B2(n_611),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_692),
.B(n_611),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_648),
.B(n_613),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_712),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_711),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_741),
.B(n_564),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_666),
.A2(n_620),
.B1(n_625),
.B2(n_613),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_707),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_704),
.B(n_620),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_704),
.B(n_620),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_712),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_704),
.B(n_625),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_790),
.B(n_581),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_714),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_714),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_727),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_711),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_727),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_707),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_747),
.B(n_564),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_751),
.B(n_641),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_669),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_768),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_730),
.A2(n_574),
.B(n_571),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_790),
.B(n_678),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_732),
.B(n_625),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_642),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_788),
.B(n_629),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_702),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_732),
.B(n_629),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_642),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_732),
.B(n_629),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_639),
.B(n_632),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_768),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_713),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_790),
.B(n_571),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_639),
.B(n_632),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_771),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_788),
.B(n_632),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_703),
.B(n_559),
.Y(n_906)
);

AOI221xp5_ASAP7_75t_L g907 ( 
.A1(n_789),
.A2(n_302),
.B1(n_345),
.B2(n_328),
.C(n_324),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_649),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_703),
.B(n_563),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_715),
.B(n_666),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_771),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_772),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_713),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_790),
.B(n_571),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_790),
.B(n_682),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_715),
.B(n_599),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_753),
.B(n_616),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_772),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_783),
.A2(n_621),
.B1(n_616),
.B2(n_319),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_776),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_753),
.B(n_621),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_762),
.B(n_574),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_776),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_781),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_717),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_710),
.B(n_574),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_710),
.B(n_574),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_781),
.Y(n_928)
);

NOR3xp33_ASAP7_75t_L g929 ( 
.A(n_638),
.B(n_270),
.C(n_269),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_783),
.A2(n_320),
.B1(n_326),
.B2(n_317),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_775),
.B(n_574),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_758),
.A2(n_570),
.B1(n_562),
.B2(n_387),
.Y(n_932)
);

O2A1O1Ixp5_ASAP7_75t_L g933 ( 
.A1(n_710),
.A2(n_398),
.B(n_390),
.C(n_380),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_782),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_755),
.B(n_574),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_718),
.B(n_574),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_651),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_720),
.B(n_575),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_717),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_711),
.B(n_269),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_725),
.B(n_687),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_645),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_764),
.A2(n_234),
.B1(n_421),
.B2(n_418),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_659),
.B(n_327),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_651),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_782),
.B(n_575),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_764),
.A2(n_777),
.B1(n_684),
.B2(n_671),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_764),
.B(n_575),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_764),
.B(n_575),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_764),
.B(n_575),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_L g951 ( 
.A(n_642),
.B(n_575),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_764),
.B(n_575),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_764),
.B(n_235),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_709),
.B(n_339),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_651),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_735),
.B(n_276),
.Y(n_956)
);

OAI22xp33_ASAP7_75t_L g957 ( 
.A1(n_670),
.A2(n_324),
.B1(n_310),
.B2(n_308),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_734),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_734),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_737),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_777),
.B(n_250),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_737),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_642),
.B(n_418),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_758),
.B(n_290),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_798),
.B(n_760),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_797),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_941),
.A2(n_671),
.B(n_644),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_836),
.B(n_733),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_936),
.A2(n_644),
.B(n_761),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_802),
.B(n_760),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_906),
.B(n_777),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_955),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_910),
.B(n_642),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_947),
.B(n_763),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_854),
.A2(n_738),
.B(n_748),
.C(n_745),
.Y(n_975)
);

NAND2xp33_ASAP7_75t_L g976 ( 
.A(n_800),
.B(n_759),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_857),
.A2(n_738),
.B(n_748),
.C(n_745),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_938),
.A2(n_767),
.B(n_761),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_909),
.B(n_777),
.Y(n_979)
);

NAND3xp33_ASAP7_75t_L g980 ( 
.A(n_806),
.B(n_819),
.C(n_826),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_926),
.A2(n_774),
.B(n_767),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_824),
.B(n_673),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_917),
.A2(n_921),
.B(n_835),
.C(n_844),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_926),
.A2(n_778),
.B(n_774),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_836),
.B(n_690),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_805),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_890),
.A2(n_754),
.B(n_652),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_838),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_799),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_841),
.A2(n_754),
.B(n_652),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_801),
.B(n_758),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_916),
.A2(n_665),
.B(n_654),
.C(n_657),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_809),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_871),
.B(n_883),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_927),
.A2(n_779),
.B(n_778),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_887),
.A2(n_940),
.B1(n_822),
.B2(n_849),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_794),
.B(n_777),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_794),
.B(n_777),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_927),
.A2(n_784),
.B(n_779),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_811),
.B(n_777),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_831),
.B(n_676),
.Y(n_1001)
);

AOI21x1_ASAP7_75t_L g1002 ( 
.A1(n_902),
.A2(n_914),
.B(n_821),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_827),
.B(n_708),
.Y(n_1003)
);

OAI21xp33_ASAP7_75t_L g1004 ( 
.A1(n_837),
.A2(n_343),
.B(n_341),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_869),
.A2(n_784),
.B(n_759),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_946),
.A2(n_654),
.B(n_646),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_922),
.A2(n_759),
.B(n_763),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_940),
.A2(n_740),
.B1(n_752),
.B2(n_758),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_837),
.B(n_752),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_940),
.A2(n_769),
.B1(n_708),
.B2(n_690),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_808),
.B(n_769),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_894),
.B(n_769),
.Y(n_1012)
);

NAND2x1p5_ASAP7_75t_L g1013 ( 
.A(n_871),
.B(n_645),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_840),
.B(n_763),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_893),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_931),
.A2(n_791),
.B(n_770),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_SL g1017 ( 
.A1(n_812),
.A2(n_657),
.B(n_660),
.C(n_646),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_820),
.B(n_769),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_940),
.B(n_744),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_883),
.B(n_770),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_955),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_804),
.Y(n_1022)
);

NOR2x1p5_ASAP7_75t_SL g1023 ( 
.A(n_828),
.B(n_787),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_832),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_908),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_905),
.A2(n_873),
.B(n_830),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_945),
.B(n_770),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_893),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_840),
.B(n_791),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_828),
.A2(n_664),
.B(n_660),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_964),
.B(n_773),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_845),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_848),
.A2(n_688),
.B1(n_645),
.B2(n_791),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_866),
.A2(n_719),
.B(n_295),
.C(n_302),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_870),
.B(n_792),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_832),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_964),
.B(n_222),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_902),
.A2(n_792),
.B(n_672),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_894),
.B(n_792),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_899),
.B(n_665),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_956),
.B(n_222),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_SL g1042 ( 
.A(n_840),
.B(n_661),
.Y(n_1042)
);

NOR2xp67_ASAP7_75t_L g1043 ( 
.A(n_937),
.B(n_665),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_903),
.B(n_875),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_914),
.A2(n_672),
.B(n_664),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_848),
.A2(n_688),
.B1(n_719),
.B2(n_679),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_876),
.B(n_688),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_878),
.B(n_674),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_830),
.A2(n_679),
.B(n_674),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_892),
.B(n_896),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_855),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_898),
.B(n_691),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_847),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_793),
.B(n_691),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_856),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_919),
.A2(n_295),
.B(n_308),
.C(n_290),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_804),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_832),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_861),
.A2(n_864),
.B(n_954),
.C(n_803),
.Y(n_1059)
);

BUFx4f_ASAP7_75t_L g1060 ( 
.A(n_945),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_862),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_812),
.A2(n_716),
.B(n_699),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_796),
.B(n_699),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_821),
.A2(n_723),
.B(n_716),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_956),
.B(n_222),
.Y(n_1065)
);

AOI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_944),
.A2(n_724),
.B(n_723),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_807),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_842),
.B(n_724),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_851),
.B(n_731),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_795),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_929),
.B(n_328),
.C(n_310),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_SL g1072 ( 
.A1(n_825),
.A2(n_865),
.B(n_879),
.C(n_850),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_825),
.A2(n_736),
.B(n_731),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_877),
.B(n_736),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_850),
.A2(n_743),
.B(n_643),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_848),
.B(n_640),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_807),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_832),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_865),
.A2(n_879),
.B(n_803),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_852),
.B(n_743),
.Y(n_1080)
);

NAND2x1p5_ASAP7_75t_L g1081 ( 
.A(n_838),
.B(n_795),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_880),
.B(n_640),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_839),
.A2(n_650),
.B(n_643),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_858),
.B(n_650),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_881),
.B(n_655),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_859),
.B(n_655),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_839),
.A2(n_662),
.B(n_656),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_882),
.B(n_656),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_848),
.A2(n_662),
.B1(n_421),
.B2(n_431),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_863),
.A2(n_402),
.B1(n_433),
.B2(n_370),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_884),
.B(n_358),
.Y(n_1091)
);

BUFx5_ASAP7_75t_L g1092 ( 
.A(n_900),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_957),
.A2(n_431),
.B1(n_406),
.B2(n_371),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_813),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_893),
.B(n_787),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_860),
.B(n_345),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_907),
.A2(n_868),
.B1(n_823),
.B2(n_810),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_893),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_867),
.B(n_362),
.Y(n_1099)
);

AOI21xp33_ASAP7_75t_L g1100 ( 
.A1(n_953),
.A2(n_381),
.B(n_377),
.Y(n_1100)
);

OAI321xp33_ASAP7_75t_L g1101 ( 
.A1(n_943),
.A2(n_372),
.A3(n_419),
.B1(n_422),
.B2(n_379),
.C(n_362),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_834),
.B(n_363),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_951),
.A2(n_594),
.B(n_227),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_893),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_813),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_900),
.A2(n_918),
.B(n_904),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_951),
.A2(n_241),
.B(n_220),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_888),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_814),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_862),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_935),
.A2(n_556),
.B(n_554),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_846),
.B(n_363),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_897),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_904),
.B(n_372),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_918),
.A2(n_417),
.B1(n_400),
.B2(n_430),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_930),
.A2(n_389),
.B(n_382),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_853),
.B(n_379),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_942),
.A2(n_253),
.B(n_247),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_895),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_942),
.A2(n_255),
.B(n_254),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_942),
.A2(n_260),
.B(n_256),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_889),
.A2(n_920),
.B1(n_911),
.B2(n_923),
.Y(n_1122)
);

AOI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_961),
.A2(n_394),
.B(n_391),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_897),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_912),
.A2(n_928),
.B(n_924),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_933),
.A2(n_570),
.B(n_562),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_934),
.A2(n_404),
.B1(n_401),
.B2(n_429),
.Y(n_1127)
);

BUFx4f_ASAP7_75t_L g1128 ( 
.A(n_847),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_897),
.A2(n_265),
.B(n_262),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_897),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_843),
.B(n_397),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_814),
.B(n_397),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_815),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_891),
.A2(n_419),
.B(n_422),
.C(n_420),
.Y(n_1134)
);

O2A1O1Ixp5_ASAP7_75t_L g1135 ( 
.A1(n_891),
.A2(n_556),
.B(n_554),
.C(n_562),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_815),
.B(n_423),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_816),
.B(n_424),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_915),
.B(n_425),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_948),
.A2(n_570),
.B(n_562),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_862),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_915),
.B(n_661),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_949),
.A2(n_570),
.B(n_562),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_959),
.A2(n_426),
.B(n_368),
.C(n_347),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_872),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_960),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_897),
.A2(n_952),
.B(n_950),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_932),
.B(n_232),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_886),
.B(n_232),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_963),
.A2(n_562),
.B1(n_570),
.B2(n_266),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_816),
.B(n_257),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_817),
.B(n_766),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_817),
.B(n_562),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_818),
.B(n_232),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_818),
.A2(n_277),
.B(n_268),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_829),
.B(n_562),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_967),
.A2(n_833),
.B(n_829),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1044),
.B(n_833),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1037),
.B(n_232),
.Y(n_1158)
);

CKINVDCx12_ASAP7_75t_R g1159 ( 
.A(n_1128),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_980),
.B(n_962),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_1078),
.Y(n_1161)
);

BUFx2_ASAP7_75t_R g1162 ( 
.A(n_1061),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1019),
.A2(n_901),
.B1(n_958),
.B2(n_939),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_976),
.A2(n_885),
.B(n_874),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1026),
.A2(n_885),
.B(n_874),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_966),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1015),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1095),
.A2(n_913),
.B(n_901),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1041),
.B(n_278),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1001),
.A2(n_963),
.B1(n_958),
.B2(n_939),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1078),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_996),
.A2(n_925),
.B1(n_913),
.B2(n_368),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_1119),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1001),
.A2(n_925),
.B1(n_278),
.B2(n_285),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_965),
.B(n_278),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_982),
.A2(n_416),
.B(n_554),
.C(n_556),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1095),
.A2(n_280),
.B(n_281),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_982),
.A2(n_278),
.B1(n_285),
.B2(n_357),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1148),
.B(n_285),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1148),
.B(n_285),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1016),
.A2(n_360),
.B(n_284),
.Y(n_1181)
);

BUFx12f_ASAP7_75t_L g1182 ( 
.A(n_1053),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1059),
.A2(n_361),
.B(n_289),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_SL g1184 ( 
.A1(n_992),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_970),
.B(n_357),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1106),
.A2(n_283),
.B(n_297),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_983),
.B(n_357),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_986),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_993),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1032),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1011),
.A2(n_357),
.B1(n_562),
.B2(n_570),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1015),
.Y(n_1192)
);

AOI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1111),
.A2(n_570),
.B(n_634),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1070),
.B(n_570),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1060),
.B(n_386),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1138),
.A2(n_416),
.B(n_298),
.C(n_374),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1012),
.B(n_570),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_1119),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1015),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1005),
.A2(n_299),
.B(n_306),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1138),
.A2(n_378),
.B(n_309),
.C(n_312),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_971),
.A2(n_634),
.B(n_766),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1021),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1060),
.B(n_386),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1025),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1065),
.B(n_386),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1102),
.A2(n_14),
.B(n_16),
.C(n_19),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1007),
.A2(n_1040),
.B(n_978),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1051),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1153),
.B(n_20),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1056),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1034),
.A2(n_307),
.B(n_314),
.C(n_315),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1011),
.B(n_22),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1144),
.B(n_25),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1019),
.B(n_25),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_989),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1025),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_979),
.A2(n_634),
.B(n_766),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1116),
.A2(n_29),
.B(n_34),
.C(n_36),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1015),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1024),
.B(n_766),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_SL g1222 ( 
.A(n_1128),
.B(n_1108),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1070),
.A2(n_318),
.B(n_322),
.C(n_332),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_972),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1055),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1010),
.B(n_386),
.Y(n_1226)
);

O2A1O1Ixp5_ASAP7_75t_SL g1227 ( 
.A1(n_1066),
.A2(n_410),
.B(n_387),
.C(n_634),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1008),
.B(n_387),
.Y(n_1228)
);

NAND3xp33_ASAP7_75t_SL g1229 ( 
.A(n_1071),
.B(n_1093),
.C(n_1004),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1003),
.B(n_37),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1097),
.A2(n_338),
.B1(n_346),
.B2(n_348),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1110),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1050),
.B(n_37),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_969),
.A2(n_393),
.B(n_351),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1097),
.A2(n_349),
.B1(n_355),
.B2(n_432),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_991),
.B(n_39),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1125),
.A2(n_405),
.B(n_375),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1071),
.A2(n_39),
.B(n_43),
.C(n_45),
.Y(n_1238)
);

INVxp67_ASAP7_75t_SL g1239 ( 
.A(n_1028),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1079),
.A2(n_408),
.B(n_384),
.C(n_388),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1018),
.B(n_392),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1076),
.B(n_766),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1031),
.A2(n_410),
.B1(n_387),
.B2(n_634),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1145),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1092),
.B(n_634),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1096),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1132),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1114),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_968),
.B(n_410),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_968),
.B(n_48),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1022),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1036),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1009),
.A2(n_428),
.B1(n_413),
.B2(n_411),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_SL g1254 ( 
.A1(n_974),
.A2(n_356),
.B(n_369),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_1140),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1076),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1092),
.B(n_634),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1134),
.A2(n_409),
.B(n_395),
.C(n_369),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1028),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1084),
.A2(n_661),
.B(n_369),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1036),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1000),
.A2(n_369),
.B(n_356),
.C(n_661),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_1009),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1135),
.A2(n_661),
.B(n_369),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1092),
.B(n_997),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1100),
.A2(n_1123),
.B(n_1020),
.C(n_998),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1020),
.A2(n_356),
.B(n_410),
.C(n_53),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1057),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1086),
.A2(n_356),
.B(n_121),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1074),
.A2(n_49),
.B(n_51),
.C(n_53),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1067),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1092),
.B(n_1039),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_988),
.B(n_124),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1054),
.A2(n_108),
.B(n_211),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1063),
.A2(n_107),
.B(n_208),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1047),
.A2(n_51),
.B(n_55),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1077),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1094),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1092),
.B(n_988),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1105),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1068),
.A2(n_128),
.B(n_205),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1092),
.B(n_1122),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_985),
.B(n_55),
.Y(n_1283)
);

O2A1O1Ixp5_ASAP7_75t_L g1284 ( 
.A1(n_974),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1058),
.B(n_60),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1109),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1048),
.B(n_61),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1058),
.B(n_61),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_985),
.Y(n_1289)
);

NOR3xp33_ASAP7_75t_SL g1290 ( 
.A(n_1115),
.B(n_64),
.C(n_65),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1052),
.B(n_66),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1074),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1091),
.B(n_67),
.Y(n_1293)
);

NAND2x1_ASAP7_75t_L g1294 ( 
.A(n_1124),
.B(n_166),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1133),
.B(n_71),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1117),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1069),
.B(n_71),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1112),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1136),
.Y(n_1299)
);

INVx5_ASAP7_75t_L g1300 ( 
.A(n_1028),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1081),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1080),
.B(n_72),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1099),
.B(n_72),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1090),
.A2(n_73),
.B1(n_74),
.B2(n_78),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_981),
.A2(n_174),
.B(n_201),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1028),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1081),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1089),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1091),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1098),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1131),
.A2(n_92),
.B1(n_140),
.B2(n_152),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1043),
.A2(n_157),
.B1(n_165),
.B2(n_169),
.Y(n_1312)
);

NOR3xp33_ASAP7_75t_L g1313 ( 
.A(n_1127),
.B(n_170),
.C(n_176),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_994),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1137),
.B(n_177),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_984),
.A2(n_186),
.B(n_187),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1072),
.A2(n_189),
.B(n_190),
.C(n_192),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1147),
.A2(n_197),
.B1(n_214),
.B2(n_1046),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1188),
.Y(n_1319)
);

AOI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1208),
.A2(n_973),
.B(n_1002),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1156),
.A2(n_973),
.B(n_999),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1282),
.A2(n_1030),
.B(n_1049),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1282),
.A2(n_1006),
.B(n_1087),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1272),
.A2(n_1083),
.B(n_1098),
.Y(n_1324)
);

AO32x2_ASAP7_75t_L g1325 ( 
.A1(n_1172),
.A2(n_1124),
.A3(n_1130),
.B1(n_1023),
.B2(n_1101),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1189),
.Y(n_1326)
);

INVx5_ASAP7_75t_L g1327 ( 
.A(n_1300),
.Y(n_1327)
);

NAND2xp33_ASAP7_75t_L g1328 ( 
.A(n_1203),
.B(n_1098),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1179),
.B(n_1150),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1293),
.A2(n_1035),
.B(n_1082),
.C(n_1088),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1190),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1266),
.A2(n_1135),
.B(n_990),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1180),
.B(n_1082),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1248),
.B(n_1113),
.Y(n_1334)
);

NOR2x1_ASAP7_75t_R g1335 ( 
.A(n_1232),
.B(n_1130),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1166),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1272),
.A2(n_1098),
.B(n_1104),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1264),
.A2(n_987),
.B(n_995),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1309),
.A2(n_1035),
.B(n_1088),
.C(n_1085),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1215),
.A2(n_1085),
.B(n_1143),
.C(n_1033),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1224),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1315),
.A2(n_1146),
.B(n_977),
.C(n_975),
.Y(n_1342)
);

AOI221x1_ASAP7_75t_L g1343 ( 
.A1(n_1308),
.A2(n_1045),
.B1(n_1075),
.B2(n_1073),
.C(n_1062),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_1255),
.Y(n_1344)
);

OAI21xp33_ASAP7_75t_L g1345 ( 
.A1(n_1276),
.A2(n_1118),
.B(n_1121),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1168),
.A2(n_1064),
.B(n_1038),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1300),
.B(n_1104),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1296),
.B(n_1113),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1298),
.B(n_1013),
.Y(n_1349)
);

BUFx2_ASAP7_75t_SL g1350 ( 
.A(n_1300),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1162),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1256),
.B(n_1104),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1165),
.A2(n_1155),
.B(n_1152),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1193),
.A2(n_1029),
.B(n_1014),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1263),
.B(n_1027),
.Y(n_1355)
);

OAI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1178),
.A2(n_1013),
.B1(n_1149),
.B2(n_1126),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1205),
.B(n_1173),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1157),
.A2(n_1164),
.B(n_1279),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1157),
.B(n_1104),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1198),
.B(n_1129),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1172),
.A2(n_1154),
.A3(n_1103),
.B(n_1120),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1216),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1260),
.A2(n_1014),
.B(n_1029),
.Y(n_1363)
);

AND3x4_ASAP7_75t_L g1364 ( 
.A(n_1290),
.B(n_1141),
.C(n_1017),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1229),
.A2(n_1139),
.B(n_1142),
.C(n_1107),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1247),
.A2(n_1141),
.B(n_1151),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1305),
.A2(n_1316),
.B(n_1269),
.Y(n_1367)
);

AO31x2_ASAP7_75t_L g1368 ( 
.A1(n_1262),
.A2(n_1042),
.A3(n_1151),
.B(n_1267),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1187),
.A2(n_1302),
.B(n_1297),
.Y(n_1369)
);

AND3x2_ASAP7_75t_L g1370 ( 
.A(n_1222),
.B(n_1158),
.C(n_1169),
.Y(n_1370)
);

BUFx12f_ASAP7_75t_L g1371 ( 
.A(n_1182),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1206),
.B(n_1299),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1289),
.Y(n_1373)
);

AO21x1_ASAP7_75t_L g1374 ( 
.A1(n_1219),
.A2(n_1213),
.B(n_1303),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1265),
.A2(n_1227),
.B(n_1317),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1297),
.A2(n_1302),
.B(n_1233),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1174),
.A2(n_1308),
.B1(n_1236),
.B2(n_1214),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1231),
.A2(n_1235),
.B1(n_1304),
.B2(n_1288),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1287),
.A2(n_1291),
.B(n_1245),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1209),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1285),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1287),
.A2(n_1291),
.B(n_1245),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1301),
.A2(n_1307),
.A3(n_1258),
.B(n_1240),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1230),
.A2(n_1303),
.B(n_1197),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1241),
.B(n_1225),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1196),
.A2(n_1210),
.B(n_1211),
.C(n_1318),
.Y(n_1386)
);

O2A1O1Ixp5_ASAP7_75t_SL g1387 ( 
.A1(n_1160),
.A2(n_1228),
.B(n_1185),
.C(n_1226),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1159),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1311),
.A2(n_1295),
.A3(n_1268),
.B(n_1278),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1244),
.Y(n_1390)
);

INVx5_ASAP7_75t_L g1391 ( 
.A(n_1300),
.Y(n_1391)
);

NAND3x1_ASAP7_75t_L g1392 ( 
.A(n_1249),
.B(n_1175),
.C(n_1313),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1194),
.A2(n_1295),
.B(n_1176),
.Y(n_1393)
);

AOI222xp33_ASAP7_75t_L g1394 ( 
.A1(n_1285),
.A2(n_1283),
.B1(n_1231),
.B2(n_1235),
.C1(n_1292),
.C2(n_1270),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1238),
.A2(n_1217),
.B(n_1207),
.C(n_1201),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1212),
.A2(n_1170),
.B1(n_1246),
.B2(n_1250),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1274),
.A2(n_1281),
.B(n_1275),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1257),
.A2(n_1273),
.B(n_1294),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1194),
.A2(n_1284),
.B(n_1183),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1195),
.B(n_1204),
.Y(n_1400)
);

NOR4xp25_ASAP7_75t_L g1401 ( 
.A(n_1184),
.B(n_1311),
.C(n_1223),
.D(n_1163),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1257),
.A2(n_1218),
.B(n_1202),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_SL g1403 ( 
.A1(n_1177),
.A2(n_1186),
.B(n_1181),
.C(n_1239),
.Y(n_1403)
);

CKINVDCx11_ASAP7_75t_R g1404 ( 
.A(n_1167),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1254),
.A2(n_1234),
.B(n_1200),
.Y(n_1405)
);

BUFx10_ASAP7_75t_L g1406 ( 
.A(n_1167),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1252),
.A2(n_1261),
.B(n_1237),
.C(n_1314),
.Y(n_1407)
);

BUFx8_ASAP7_75t_L g1408 ( 
.A(n_1167),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1192),
.A2(n_1220),
.B(n_1306),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1256),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1171),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1161),
.B(n_1171),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1192),
.A2(n_1259),
.B(n_1310),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1271),
.A2(n_1277),
.B1(n_1251),
.B2(n_1286),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1161),
.B(n_1280),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1253),
.A2(n_1191),
.B1(n_1312),
.B2(n_1273),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1192),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1199),
.A2(n_1220),
.B(n_1259),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1199),
.A2(n_1220),
.B(n_1259),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1199),
.B(n_1306),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1306),
.Y(n_1421)
);

AOI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1221),
.A2(n_1310),
.B(n_1242),
.Y(n_1422)
);

AO31x2_ASAP7_75t_L g1423 ( 
.A1(n_1243),
.A2(n_1310),
.A3(n_1242),
.B(n_1221),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1203),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_SL g1425 ( 
.A1(n_1293),
.A2(n_1211),
.B1(n_1276),
.B2(n_1238),
.C(n_689),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1208),
.A2(n_1111),
.B(n_1156),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1293),
.A2(n_798),
.B(n_980),
.C(n_982),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1208),
.A2(n_1282),
.B(n_1165),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1282),
.A2(n_798),
.B(n_967),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1188),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1166),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1208),
.A2(n_1111),
.B(n_1156),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1179),
.B(n_798),
.Y(n_1433)
);

INVx5_ASAP7_75t_L g1434 ( 
.A(n_1300),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1166),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1208),
.A2(n_1111),
.B(n_1156),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1282),
.A2(n_798),
.B(n_967),
.Y(n_1437)
);

AO31x2_ASAP7_75t_L g1438 ( 
.A1(n_1208),
.A2(n_1165),
.A3(n_1282),
.B(n_1059),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1166),
.Y(n_1439)
);

INVxp67_ASAP7_75t_SL g1440 ( 
.A(n_1173),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1282),
.A2(n_1059),
.B(n_798),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1188),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1161),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1203),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1282),
.A2(n_798),
.B(n_967),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1293),
.A2(n_798),
.B(n_980),
.C(n_1001),
.Y(n_1446)
);

BUFx12f_ASAP7_75t_L g1447 ( 
.A(n_1203),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1309),
.B(n_996),
.Y(n_1448)
);

AND2x6_ASAP7_75t_L g1449 ( 
.A(n_1285),
.B(n_1256),
.Y(n_1449)
);

NOR2xp67_ASAP7_75t_SL g1450 ( 
.A(n_1203),
.B(n_955),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1208),
.A2(n_1111),
.B(n_1156),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1208),
.A2(n_1111),
.B(n_1156),
.Y(n_1452)
);

AO32x2_ASAP7_75t_L g1453 ( 
.A1(n_1172),
.A2(n_1308),
.A3(n_689),
.B1(n_1235),
.B2(n_1231),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1179),
.B(n_798),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1282),
.A2(n_798),
.B(n_967),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1203),
.Y(n_1456)
);

BUFx10_ASAP7_75t_L g1457 ( 
.A(n_1203),
.Y(n_1457)
);

AO31x2_ASAP7_75t_L g1458 ( 
.A1(n_1208),
.A2(n_1165),
.A3(n_1282),
.B(n_1059),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1179),
.B(n_798),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1282),
.A2(n_798),
.B(n_967),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1179),
.B(n_798),
.Y(n_1461)
);

BUFx12f_ASAP7_75t_L g1462 ( 
.A(n_1203),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1188),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1309),
.B(n_996),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1179),
.B(n_798),
.Y(n_1465)
);

AO31x2_ASAP7_75t_L g1466 ( 
.A1(n_1208),
.A2(n_1165),
.A3(n_1282),
.B(n_1059),
.Y(n_1466)
);

A2O1A1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1293),
.A2(n_798),
.B(n_980),
.C(n_982),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1248),
.B(n_1157),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1248),
.B(n_1157),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1248),
.B(n_1157),
.Y(n_1470)
);

AOI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1293),
.A2(n_980),
.B1(n_1001),
.B2(n_826),
.C(n_806),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1282),
.A2(n_1059),
.B(n_798),
.Y(n_1472)
);

BUFx8_ASAP7_75t_SL g1473 ( 
.A(n_1255),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1179),
.B(n_798),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1208),
.A2(n_1165),
.A3(n_1282),
.B(n_1059),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1300),
.Y(n_1476)
);

AO22x2_ASAP7_75t_L g1477 ( 
.A1(n_1229),
.A2(n_980),
.B1(n_1215),
.B2(n_1226),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1188),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1224),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1203),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1179),
.B(n_798),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1282),
.A2(n_798),
.B(n_967),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1179),
.B(n_798),
.Y(n_1483)
);

O2A1O1Ixp33_ASAP7_75t_SL g1484 ( 
.A1(n_1282),
.A2(n_798),
.B(n_1293),
.C(n_1279),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1293),
.A2(n_798),
.B1(n_996),
.B2(n_1309),
.Y(n_1485)
);

AO32x2_ASAP7_75t_L g1486 ( 
.A1(n_1172),
.A2(n_1308),
.A3(n_689),
.B1(n_1235),
.B2(n_1231),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_SL g1487 ( 
.A1(n_1282),
.A2(n_798),
.B(n_1293),
.C(n_1279),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1208),
.A2(n_1111),
.B(n_1156),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1282),
.A2(n_798),
.B(n_967),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1166),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1158),
.B(n_801),
.Y(n_1491)
);

O2A1O1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1293),
.A2(n_798),
.B(n_980),
.C(n_1001),
.Y(n_1492)
);

O2A1O1Ixp5_ASAP7_75t_L g1493 ( 
.A1(n_1179),
.A2(n_1180),
.B(n_798),
.C(n_1293),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1471),
.A2(n_1378),
.B1(n_1485),
.B2(n_1454),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1378),
.A2(n_1485),
.B1(n_1433),
.B2(n_1459),
.Y(n_1495)
);

BUFx10_ASAP7_75t_L g1496 ( 
.A(n_1351),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1477),
.A2(n_1461),
.B1(n_1465),
.B2(n_1483),
.Y(n_1497)
);

INVx6_ASAP7_75t_L g1498 ( 
.A(n_1408),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1394),
.A2(n_1377),
.B1(n_1474),
.B2(n_1481),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1473),
.Y(n_1500)
);

CKINVDCx11_ASAP7_75t_R g1501 ( 
.A(n_1344),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1319),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1388),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1394),
.A2(n_1477),
.B1(n_1464),
.B2(n_1448),
.Y(n_1504)
);

CKINVDCx11_ASAP7_75t_R g1505 ( 
.A(n_1371),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1326),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1333),
.A2(n_1329),
.B1(n_1374),
.B2(n_1370),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1426),
.A2(n_1436),
.B(n_1432),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1327),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1385),
.A2(n_1372),
.B1(n_1396),
.B2(n_1376),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1362),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1331),
.Y(n_1512)
);

CKINVDCx11_ASAP7_75t_R g1513 ( 
.A(n_1457),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1380),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_SL g1515 ( 
.A(n_1457),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1408),
.Y(n_1516)
);

BUFx2_ASAP7_75t_SL g1517 ( 
.A(n_1456),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1327),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1427),
.A2(n_1467),
.B1(n_1492),
.B2(n_1446),
.Y(n_1519)
);

OAI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1381),
.A2(n_1441),
.B1(n_1472),
.B2(n_1416),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1390),
.Y(n_1521)
);

INVx5_ASAP7_75t_L g1522 ( 
.A(n_1449),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1396),
.A2(n_1449),
.B1(n_1472),
.B2(n_1441),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1449),
.A2(n_1469),
.B1(n_1468),
.B2(n_1470),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1430),
.Y(n_1525)
);

INVx6_ASAP7_75t_L g1526 ( 
.A(n_1391),
.Y(n_1526)
);

INVx6_ASAP7_75t_L g1527 ( 
.A(n_1391),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1424),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1447),
.Y(n_1529)
);

INVx8_ASAP7_75t_L g1530 ( 
.A(n_1449),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1386),
.A2(n_1330),
.B1(n_1364),
.B2(n_1392),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1391),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1442),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1341),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1438),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1416),
.A2(n_1453),
.B1(n_1486),
.B2(n_1325),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1440),
.B(n_1357),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1463),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1355),
.A2(n_1339),
.B1(n_1395),
.B2(n_1493),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1479),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1468),
.B(n_1469),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1425),
.A2(n_1400),
.B1(n_1479),
.B2(n_1356),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1360),
.A2(n_1340),
.B1(n_1322),
.B2(n_1470),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1453),
.A2(n_1486),
.B1(n_1325),
.B2(n_1369),
.Y(n_1544)
);

BUFx12f_ASAP7_75t_L g1545 ( 
.A(n_1404),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1462),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1478),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1453),
.A2(n_1486),
.B1(n_1325),
.B2(n_1369),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1384),
.A2(n_1490),
.B1(n_1439),
.B2(n_1431),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1384),
.A2(n_1435),
.B1(n_1345),
.B2(n_1334),
.Y(n_1550)
);

BUFx10_ASAP7_75t_L g1551 ( 
.A(n_1480),
.Y(n_1551)
);

OAI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1334),
.A2(n_1348),
.B1(n_1359),
.B2(n_1349),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_SL g1553 ( 
.A1(n_1332),
.A2(n_1425),
.B1(n_1393),
.B2(n_1401),
.Y(n_1553)
);

BUFx12f_ASAP7_75t_L g1554 ( 
.A(n_1444),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1345),
.A2(n_1414),
.B1(n_1332),
.B2(n_1373),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1415),
.B(n_1412),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1421),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1365),
.A2(n_1443),
.B1(n_1407),
.B2(n_1382),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1443),
.A2(n_1379),
.B1(n_1482),
.B2(n_1437),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1489),
.A2(n_1455),
.B1(n_1429),
.B2(n_1460),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1393),
.A2(n_1399),
.B1(n_1359),
.B2(n_1352),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1406),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1399),
.A2(n_1352),
.B1(n_1328),
.B2(n_1450),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1402),
.A2(n_1412),
.B1(n_1405),
.B2(n_1358),
.Y(n_1565)
);

BUFx8_ASAP7_75t_L g1566 ( 
.A(n_1476),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1417),
.A2(n_1337),
.B1(n_1476),
.B2(n_1350),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1401),
.A2(n_1434),
.B1(n_1323),
.B2(n_1445),
.Y(n_1568)
);

OAI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1434),
.A2(n_1343),
.B1(n_1476),
.B2(n_1417),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_SL g1570 ( 
.A1(n_1342),
.A2(n_1487),
.B(n_1484),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1406),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1347),
.A2(n_1422),
.B1(n_1324),
.B2(n_1418),
.Y(n_1572)
);

OAI21xp33_ASAP7_75t_L g1573 ( 
.A1(n_1387),
.A2(n_1366),
.B(n_1397),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1335),
.Y(n_1574)
);

INVx6_ASAP7_75t_L g1575 ( 
.A(n_1347),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1375),
.A2(n_1420),
.B1(n_1353),
.B2(n_1354),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1409),
.B(n_1419),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1428),
.A2(n_1367),
.B1(n_1346),
.B2(n_1398),
.Y(n_1578)
);

CKINVDCx11_ASAP7_75t_R g1579 ( 
.A(n_1413),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1428),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1383),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1389),
.Y(n_1582)
);

INVx6_ASAP7_75t_L g1583 ( 
.A(n_1423),
.Y(n_1583)
);

BUFx2_ASAP7_75t_SL g1584 ( 
.A(n_1423),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1320),
.A2(n_1346),
.B1(n_1321),
.B2(n_1475),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1423),
.A2(n_1368),
.B1(n_1363),
.B2(n_1361),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1338),
.A2(n_1451),
.B1(n_1452),
.B2(n_1488),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1383),
.A2(n_1403),
.B1(n_1368),
.B2(n_1361),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1368),
.A2(n_1361),
.B1(n_1438),
.B2(n_1458),
.Y(n_1589)
);

CKINVDCx6p67_ASAP7_75t_R g1590 ( 
.A(n_1458),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1466),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1319),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1319),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1344),
.Y(n_1594)
);

OAI21xp33_ASAP7_75t_L g1595 ( 
.A1(n_1433),
.A2(n_1459),
.B(n_1454),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1327),
.Y(n_1596)
);

INVx5_ASAP7_75t_L g1597 ( 
.A(n_1449),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1319),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1319),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1327),
.Y(n_1600)
);

BUFx12f_ASAP7_75t_L g1601 ( 
.A(n_1351),
.Y(n_1601)
);

BUFx2_ASAP7_75t_SL g1602 ( 
.A(n_1344),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1433),
.B(n_1454),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1319),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1319),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1471),
.A2(n_1180),
.B1(n_1179),
.B2(n_826),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1433),
.A2(n_1454),
.B1(n_1461),
.B2(n_1459),
.Y(n_1607)
);

CKINVDCx11_ASAP7_75t_R g1608 ( 
.A(n_1344),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1471),
.A2(n_1019),
.B1(n_824),
.B2(n_826),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1491),
.B(n_991),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1336),
.Y(n_1611)
);

INVx4_ASAP7_75t_L g1612 ( 
.A(n_1327),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_SL g1613 ( 
.A1(n_1471),
.A2(n_1378),
.B(n_1433),
.Y(n_1613)
);

CKINVDCx11_ASAP7_75t_R g1614 ( 
.A(n_1344),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1408),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1319),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1471),
.A2(n_1019),
.B1(n_824),
.B2(n_826),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1336),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1473),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1433),
.B(n_1001),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1471),
.A2(n_1019),
.B1(n_824),
.B2(n_826),
.Y(n_1621)
);

BUFx12f_ASAP7_75t_L g1622 ( 
.A(n_1351),
.Y(n_1622)
);

BUFx10_ASAP7_75t_L g1623 ( 
.A(n_1351),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1327),
.Y(n_1624)
);

INVx3_ASAP7_75t_SL g1625 ( 
.A(n_1424),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1330),
.A2(n_824),
.B(n_1333),
.Y(n_1626)
);

CKINVDCx11_ASAP7_75t_R g1627 ( 
.A(n_1344),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1433),
.B(n_1454),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1319),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1471),
.A2(n_1180),
.B1(n_1179),
.B2(n_826),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1433),
.A2(n_1454),
.B1(n_1461),
.B2(n_1459),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1471),
.A2(n_1019),
.B1(n_824),
.B2(n_826),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1471),
.A2(n_1019),
.B1(n_824),
.B2(n_826),
.Y(n_1633)
);

OAI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1378),
.A2(n_1454),
.B1(n_1459),
.B2(n_1433),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1319),
.Y(n_1635)
);

INVx6_ASAP7_75t_L g1636 ( 
.A(n_1408),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1327),
.Y(n_1637)
);

INVx6_ASAP7_75t_L g1638 ( 
.A(n_1408),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1433),
.A2(n_1454),
.B1(n_1461),
.B2(n_1459),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1433),
.A2(n_1454),
.B1(n_1461),
.B2(n_1459),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1473),
.Y(n_1641)
);

INVx8_ASAP7_75t_L g1642 ( 
.A(n_1449),
.Y(n_1642)
);

BUFx12f_ASAP7_75t_L g1643 ( 
.A(n_1351),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1344),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1471),
.A2(n_826),
.B1(n_824),
.B2(n_831),
.Y(n_1645)
);

OAI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1378),
.A2(n_1454),
.B1(n_1459),
.B2(n_1433),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_SL g1647 ( 
.A1(n_1485),
.A2(n_1019),
.B1(n_824),
.B2(n_1179),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1319),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1485),
.A2(n_1019),
.B1(n_824),
.B2(n_1179),
.Y(n_1649)
);

CKINVDCx20_ASAP7_75t_R g1650 ( 
.A(n_1473),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1471),
.A2(n_826),
.B1(n_824),
.B2(n_831),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1471),
.A2(n_1180),
.B1(n_1179),
.B2(n_826),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1494),
.A2(n_1495),
.B1(n_1499),
.B2(n_1613),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1534),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1498),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1634),
.B(n_1646),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1536),
.B(n_1544),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1536),
.B(n_1544),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1540),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1548),
.B(n_1502),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1582),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1591),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1535),
.Y(n_1663)
);

OAI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1561),
.A2(n_1578),
.B(n_1587),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1579),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1537),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1535),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1501),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1498),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1541),
.B(n_1548),
.Y(n_1670)
);

OA21x2_ASAP7_75t_L g1671 ( 
.A1(n_1578),
.A2(n_1573),
.B(n_1570),
.Y(n_1671)
);

BUFx8_ASAP7_75t_L g1672 ( 
.A(n_1515),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1583),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1620),
.B(n_1607),
.Y(n_1674)
);

NAND2x1_ASAP7_75t_L g1675 ( 
.A(n_1565),
.B(n_1559),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1522),
.B(n_1597),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1508),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1506),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1560),
.A2(n_1576),
.B(n_1508),
.Y(n_1679)
);

AO21x2_ASAP7_75t_L g1680 ( 
.A1(n_1585),
.A2(n_1552),
.B(n_1569),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1512),
.Y(n_1681)
);

BUFx3_ASAP7_75t_L g1682 ( 
.A(n_1583),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1590),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1514),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1521),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1525),
.B(n_1533),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1583),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1538),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1522),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1634),
.A2(n_1646),
.B1(n_1630),
.B2(n_1652),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1580),
.Y(n_1691)
);

OA21x2_ASAP7_75t_L g1692 ( 
.A1(n_1581),
.A2(n_1550),
.B(n_1523),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1606),
.A2(n_1531),
.B1(n_1542),
.B2(n_1520),
.Y(n_1693)
);

OAI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1577),
.A2(n_1550),
.B(n_1543),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1547),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1610),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1592),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1523),
.A2(n_1562),
.B(n_1555),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1593),
.B(n_1598),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1599),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1604),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1605),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1555),
.A2(n_1539),
.B(n_1567),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1616),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1629),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1635),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1648),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1584),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1588),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1553),
.B(n_1589),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1552),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1504),
.B(n_1495),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1553),
.B(n_1589),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1586),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1586),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1524),
.B(n_1494),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1585),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1549),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1557),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1498),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1549),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1520),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1511),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1611),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1519),
.A2(n_1564),
.B(n_1510),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1524),
.B(n_1510),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1596),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1618),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1558),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1596),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1569),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1631),
.B(n_1639),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1636),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1566),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1597),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1572),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1636),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1556),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1608),
.Y(n_1739)
);

CKINVDCx16_ASAP7_75t_R g1740 ( 
.A(n_1545),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1572),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1568),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1568),
.Y(n_1743)
);

BUFx6f_ASAP7_75t_L g1744 ( 
.A(n_1597),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1575),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1497),
.B(n_1507),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1497),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1597),
.B(n_1509),
.Y(n_1748)
);

OA21x2_ASAP7_75t_L g1749 ( 
.A1(n_1609),
.A2(n_1632),
.B(n_1633),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1640),
.B(n_1603),
.Y(n_1750)
);

OAI21x1_ASAP7_75t_L g1751 ( 
.A1(n_1509),
.A2(n_1624),
.B(n_1637),
.Y(n_1751)
);

BUFx2_ASAP7_75t_L g1752 ( 
.A(n_1532),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1612),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1532),
.Y(n_1754)
);

INVx4_ASAP7_75t_L g1755 ( 
.A(n_1530),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1624),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1637),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1518),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1518),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1612),
.Y(n_1760)
);

OAI21x1_ASAP7_75t_L g1761 ( 
.A1(n_1626),
.A2(n_1621),
.B(n_1617),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1628),
.B(n_1595),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1638),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1647),
.A2(n_1649),
.B1(n_1632),
.B2(n_1609),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1647),
.B(n_1649),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1517),
.B(n_1516),
.Y(n_1766)
);

AO21x1_ASAP7_75t_L g1767 ( 
.A1(n_1617),
.A2(n_1633),
.B(n_1621),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1600),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1566),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1651),
.A2(n_1645),
.B(n_1642),
.Y(n_1770)
);

OAI21x1_ASAP7_75t_L g1771 ( 
.A1(n_1526),
.A2(n_1527),
.B(n_1642),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1654),
.B(n_1602),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1654),
.B(n_1615),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1701),
.Y(n_1774)
);

OA21x2_ASAP7_75t_L g1775 ( 
.A1(n_1694),
.A2(n_1571),
.B(n_1574),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1675),
.A2(n_1530),
.B(n_1563),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1659),
.B(n_1551),
.Y(n_1777)
);

INVx4_ASAP7_75t_L g1778 ( 
.A(n_1758),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1683),
.B(n_1503),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1653),
.A2(n_1638),
.B1(n_1594),
.B2(n_1644),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1666),
.B(n_1625),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1701),
.Y(n_1782)
);

BUFx3_ASAP7_75t_L g1783 ( 
.A(n_1668),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1690),
.A2(n_1638),
.B1(n_1515),
.B2(n_1650),
.Y(n_1784)
);

OAI21x1_ASAP7_75t_SL g1785 ( 
.A1(n_1690),
.A2(n_1513),
.B(n_1505),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1656),
.A2(n_1653),
.B(n_1761),
.Y(n_1786)
);

AO21x2_ASAP7_75t_L g1787 ( 
.A1(n_1717),
.A2(n_1496),
.B(n_1623),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1739),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1675),
.A2(n_1732),
.B(n_1680),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1683),
.B(n_1546),
.Y(n_1790)
);

OA21x2_ASAP7_75t_L g1791 ( 
.A1(n_1694),
.A2(n_1679),
.B(n_1664),
.Y(n_1791)
);

AOI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1693),
.A2(n_1732),
.B1(n_1765),
.B2(n_1674),
.C(n_1767),
.Y(n_1792)
);

AOI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1765),
.A2(n_1529),
.B1(n_1500),
.B2(n_1619),
.C(n_1641),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1764),
.B(n_1627),
.C(n_1614),
.Y(n_1794)
);

AOI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1767),
.A2(n_1622),
.B1(n_1601),
.B2(n_1643),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1696),
.B(n_1496),
.Y(n_1796)
);

INVxp67_ASAP7_75t_L g1797 ( 
.A(n_1738),
.Y(n_1797)
);

AO21x1_ASAP7_75t_L g1798 ( 
.A1(n_1750),
.A2(n_1713),
.B(n_1710),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1752),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1722),
.B(n_1554),
.Y(n_1800)
);

OAI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1761),
.A2(n_1528),
.B(n_1725),
.Y(n_1801)
);

A2O1A1Ixp33_ASAP7_75t_SL g1802 ( 
.A1(n_1727),
.A2(n_1753),
.B(n_1760),
.C(n_1730),
.Y(n_1802)
);

A2O1A1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1770),
.A2(n_1746),
.B(n_1712),
.C(n_1716),
.Y(n_1803)
);

A2O1A1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1746),
.A2(n_1712),
.B(n_1716),
.C(n_1726),
.Y(n_1804)
);

AO32x2_ASAP7_75t_L g1805 ( 
.A1(n_1655),
.A2(n_1763),
.A3(n_1669),
.B1(n_1733),
.B2(n_1737),
.Y(n_1805)
);

AO32x2_ASAP7_75t_L g1806 ( 
.A1(n_1655),
.A2(n_1763),
.A3(n_1669),
.B1(n_1733),
.B2(n_1737),
.Y(n_1806)
);

A2O1A1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1726),
.A2(n_1703),
.B(n_1725),
.C(n_1743),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1686),
.B(n_1699),
.Y(n_1808)
);

O2A1O1Ixp33_ASAP7_75t_L g1809 ( 
.A1(n_1749),
.A2(n_1722),
.B(n_1742),
.C(n_1743),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1749),
.A2(n_1713),
.B1(n_1710),
.B2(n_1747),
.Y(n_1810)
);

AO22x2_ASAP7_75t_L g1811 ( 
.A1(n_1747),
.A2(n_1715),
.B1(n_1714),
.B2(n_1709),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1683),
.B(n_1665),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1719),
.B(n_1670),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1665),
.B(n_1682),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1711),
.B(n_1762),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_SL g1816 ( 
.A1(n_1749),
.A2(n_1740),
.B1(n_1731),
.B2(n_1742),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1711),
.B(n_1762),
.Y(n_1817)
);

AO21x1_ASAP7_75t_L g1818 ( 
.A1(n_1709),
.A2(n_1670),
.B(n_1698),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1766),
.B(n_1660),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1682),
.B(n_1752),
.Y(n_1820)
);

A2O1A1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1703),
.A2(n_1731),
.B(n_1698),
.C(n_1657),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1729),
.B(n_1720),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_SL g1823 ( 
.A1(n_1749),
.A2(n_1676),
.B(n_1680),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1768),
.B(n_1678),
.Y(n_1824)
);

OA21x2_ASAP7_75t_L g1825 ( 
.A1(n_1679),
.A2(n_1664),
.B(n_1717),
.Y(n_1825)
);

NAND4xp25_ASAP7_75t_L g1826 ( 
.A(n_1657),
.B(n_1658),
.C(n_1677),
.D(n_1715),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1658),
.A2(n_1680),
.B1(n_1692),
.B2(n_1714),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1707),
.B(n_1681),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1677),
.A2(n_1751),
.B(n_1771),
.Y(n_1829)
);

A2O1A1Ixp33_ASAP7_75t_L g1830 ( 
.A1(n_1736),
.A2(n_1741),
.B(n_1718),
.C(n_1721),
.Y(n_1830)
);

OAI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1671),
.A2(n_1692),
.B(n_1736),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1676),
.B(n_1745),
.Y(n_1832)
);

AO32x2_ASAP7_75t_L g1833 ( 
.A1(n_1755),
.A2(n_1692),
.A3(n_1685),
.B1(n_1684),
.B2(n_1688),
.Y(n_1833)
);

O2A1O1Ixp33_ASAP7_75t_L g1834 ( 
.A1(n_1741),
.A2(n_1671),
.B(n_1769),
.C(n_1734),
.Y(n_1834)
);

AOI221xp5_ASAP7_75t_L g1835 ( 
.A1(n_1695),
.A2(n_1697),
.B1(n_1704),
.B2(n_1706),
.C(n_1705),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1695),
.Y(n_1836)
);

BUFx3_ASAP7_75t_L g1837 ( 
.A(n_1734),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1697),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1700),
.Y(n_1839)
);

AO32x2_ASAP7_75t_L g1840 ( 
.A1(n_1755),
.A2(n_1702),
.A3(n_1704),
.B1(n_1705),
.B2(n_1706),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_SL g1841 ( 
.A1(n_1816),
.A2(n_1671),
.B1(n_1744),
.B2(n_1689),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1839),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1815),
.B(n_1663),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1840),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1783),
.B(n_1740),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1789),
.B(n_1671),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1815),
.B(n_1663),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1774),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1782),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1808),
.B(n_1667),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1816),
.A2(n_1735),
.B1(n_1744),
.B2(n_1689),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1799),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1840),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1805),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1819),
.B(n_1677),
.Y(n_1855)
);

INVx2_ASAP7_75t_SL g1856 ( 
.A(n_1812),
.Y(n_1856)
);

NOR2x1_ASAP7_75t_L g1857 ( 
.A(n_1787),
.B(n_1754),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1840),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1828),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1828),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1836),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1838),
.Y(n_1862)
);

NOR2xp67_ASAP7_75t_L g1863 ( 
.A(n_1789),
.B(n_1778),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1797),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1824),
.Y(n_1865)
);

BUFx2_ASAP7_75t_L g1866 ( 
.A(n_1805),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1798),
.A2(n_1673),
.B1(n_1687),
.B2(n_1724),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1820),
.B(n_1756),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1817),
.Y(n_1869)
);

INVxp67_ASAP7_75t_SL g1870 ( 
.A(n_1775),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1829),
.B(n_1708),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1817),
.B(n_1757),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1787),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1826),
.A2(n_1673),
.B1(n_1687),
.B2(n_1724),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1835),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1835),
.B(n_1757),
.Y(n_1876)
);

NOR2x1_ASAP7_75t_L g1877 ( 
.A(n_1801),
.B(n_1727),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1792),
.B(n_1759),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1832),
.B(n_1748),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1792),
.A2(n_1755),
.B1(n_1734),
.B2(n_1769),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1833),
.Y(n_1881)
);

OAI22xp33_ASAP7_75t_SL g1882 ( 
.A1(n_1810),
.A2(n_1723),
.B1(n_1728),
.B2(n_1691),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1833),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1833),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1805),
.B(n_1662),
.Y(n_1885)
);

INVxp67_ASAP7_75t_L g1886 ( 
.A(n_1873),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_SL g1887 ( 
.A(n_1875),
.B(n_1786),
.Y(n_1887)
);

OAI321xp33_ASAP7_75t_L g1888 ( 
.A1(n_1875),
.A2(n_1786),
.A3(n_1826),
.B1(n_1810),
.B2(n_1803),
.C(n_1827),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1854),
.B(n_1772),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1848),
.Y(n_1890)
);

NAND4xp25_ASAP7_75t_L g1891 ( 
.A(n_1878),
.B(n_1794),
.C(n_1793),
.D(n_1780),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1841),
.A2(n_1818),
.B1(n_1827),
.B2(n_1811),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1843),
.B(n_1813),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1848),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1854),
.B(n_1773),
.Y(n_1895)
);

AO21x2_ASAP7_75t_L g1896 ( 
.A1(n_1846),
.A2(n_1831),
.B(n_1821),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1866),
.B(n_1773),
.Y(n_1897)
);

OAI31xp33_ASAP7_75t_L g1898 ( 
.A1(n_1882),
.A2(n_1804),
.A3(n_1807),
.B(n_1794),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1885),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1866),
.B(n_1781),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1844),
.Y(n_1901)
);

AOI221xp5_ASAP7_75t_L g1902 ( 
.A1(n_1882),
.A2(n_1809),
.B1(n_1811),
.B2(n_1834),
.C(n_1784),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1855),
.B(n_1777),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1849),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1844),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1855),
.B(n_1806),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1874),
.A2(n_1831),
.B1(n_1795),
.B2(n_1780),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1881),
.A2(n_1809),
.B1(n_1834),
.B2(n_1784),
.C(n_1823),
.Y(n_1908)
);

OAI221xp5_ASAP7_75t_L g1909 ( 
.A1(n_1867),
.A2(n_1795),
.B1(n_1830),
.B2(n_1793),
.C(n_1800),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1865),
.B(n_1806),
.Y(n_1910)
);

INVxp67_ASAP7_75t_L g1911 ( 
.A(n_1857),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1859),
.B(n_1825),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1849),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1859),
.B(n_1825),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_SL g1915 ( 
.A(n_1880),
.B(n_1800),
.C(n_1776),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1850),
.B(n_1806),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1844),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1853),
.Y(n_1918)
);

AO21x2_ASAP7_75t_L g1919 ( 
.A1(n_1870),
.A2(n_1691),
.B(n_1661),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1871),
.Y(n_1920)
);

INVx4_ASAP7_75t_R g1921 ( 
.A(n_1856),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1860),
.B(n_1869),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1843),
.B(n_1791),
.Y(n_1923)
);

NAND3xp33_ASAP7_75t_L g1924 ( 
.A(n_1876),
.B(n_1791),
.C(n_1672),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_1852),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1853),
.Y(n_1926)
);

INVx5_ASAP7_75t_SL g1927 ( 
.A(n_1871),
.Y(n_1927)
);

OR2x4_ASAP7_75t_L g1928 ( 
.A(n_1845),
.B(n_1822),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1853),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1851),
.A2(n_1864),
.B1(n_1858),
.B2(n_1877),
.Y(n_1930)
);

INVx3_ASAP7_75t_L g1931 ( 
.A(n_1871),
.Y(n_1931)
);

AND2x2_ASAP7_75t_SL g1932 ( 
.A(n_1858),
.B(n_1814),
.Y(n_1932)
);

NAND4xp25_ASAP7_75t_L g1933 ( 
.A(n_1842),
.B(n_1796),
.C(n_1802),
.D(n_1788),
.Y(n_1933)
);

INVx2_ASAP7_75t_SL g1934 ( 
.A(n_1921),
.Y(n_1934)
);

NOR2x1p5_ASAP7_75t_L g1935 ( 
.A(n_1891),
.B(n_1769),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1906),
.B(n_1858),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1893),
.B(n_1847),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1890),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1890),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1916),
.B(n_1863),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1893),
.B(n_1847),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1894),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1910),
.B(n_1884),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1910),
.B(n_1884),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1932),
.B(n_1852),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1932),
.B(n_1872),
.Y(n_1946)
);

NOR2xp67_ASAP7_75t_SL g1947 ( 
.A(n_1888),
.B(n_1837),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1922),
.B(n_1860),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1894),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1920),
.B(n_1871),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1904),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1922),
.B(n_1881),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1932),
.B(n_1872),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1928),
.B(n_1790),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1925),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1928),
.Y(n_1956)
);

NOR2xp67_ASAP7_75t_L g1957 ( 
.A(n_1911),
.B(n_1883),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1899),
.B(n_1842),
.Y(n_1958)
);

BUFx2_ASAP7_75t_L g1959 ( 
.A(n_1928),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1887),
.Y(n_1960)
);

HB1xp67_ASAP7_75t_L g1961 ( 
.A(n_1901),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1912),
.B(n_1861),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1919),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1927),
.B(n_1868),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1901),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1912),
.B(n_1861),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1920),
.B(n_1877),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1927),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1930),
.B(n_1879),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1927),
.B(n_1868),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1920),
.B(n_1879),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1927),
.B(n_1895),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1904),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1913),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1914),
.B(n_1862),
.Y(n_1975)
);

NOR2x1_ASAP7_75t_L g1976 ( 
.A(n_1933),
.B(n_1790),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1919),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1968),
.B(n_1931),
.Y(n_1978)
);

INVx2_ASAP7_75t_SL g1979 ( 
.A(n_1968),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1938),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1938),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1976),
.A2(n_1928),
.B1(n_1909),
.B2(n_1892),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1976),
.B(n_1927),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1937),
.B(n_1923),
.Y(n_1984)
);

BUFx2_ASAP7_75t_L g1985 ( 
.A(n_1956),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1939),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1972),
.B(n_1895),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1937),
.B(n_1941),
.Y(n_1988)
);

NAND2x2_ASAP7_75t_L g1989 ( 
.A(n_1935),
.B(n_1672),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1955),
.B(n_1914),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1940),
.B(n_1931),
.Y(n_1991)
);

INVxp67_ASAP7_75t_SL g1992 ( 
.A(n_1960),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1940),
.B(n_1931),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1972),
.B(n_1897),
.Y(n_1994)
);

INVx3_ASAP7_75t_L g1995 ( 
.A(n_1968),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1963),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1955),
.B(n_1941),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1940),
.B(n_1946),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1948),
.B(n_1905),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1961),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1972),
.B(n_1897),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1958),
.B(n_1923),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1963),
.Y(n_2003)
);

INVx1_ASAP7_75t_SL g2004 ( 
.A(n_1956),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1948),
.B(n_1905),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1946),
.B(n_1953),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1963),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1939),
.Y(n_2008)
);

AND2x4_ASAP7_75t_SL g2009 ( 
.A(n_1968),
.B(n_1900),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1942),
.Y(n_2010)
);

NOR2x1p5_ASAP7_75t_L g2011 ( 
.A(n_1971),
.B(n_1891),
.Y(n_2011)
);

AOI221xp5_ASAP7_75t_L g2012 ( 
.A1(n_1969),
.A2(n_1930),
.B1(n_1888),
.B2(n_1898),
.C(n_1908),
.Y(n_2012)
);

NAND2x1p5_ASAP7_75t_L g2013 ( 
.A(n_1947),
.B(n_1857),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1946),
.B(n_1900),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1942),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1949),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1949),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1958),
.B(n_1917),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1953),
.B(n_1889),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1953),
.B(n_1959),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1959),
.B(n_1889),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1934),
.B(n_1931),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1951),
.B(n_1917),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1934),
.B(n_1903),
.Y(n_2024)
);

NOR2x1p5_ASAP7_75t_L g2025 ( 
.A(n_1971),
.B(n_1915),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1951),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1977),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1973),
.B(n_1917),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_2025),
.B(n_1934),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2025),
.B(n_1936),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_2013),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1988),
.B(n_1997),
.Y(n_2032)
);

AOI221x1_ASAP7_75t_SL g2033 ( 
.A1(n_1982),
.A2(n_1957),
.B1(n_1952),
.B2(n_1933),
.C(n_1954),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_2012),
.B(n_1961),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2006),
.B(n_1936),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_2006),
.B(n_1936),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_SL g2037 ( 
.A1(n_2012),
.A2(n_2011),
.B(n_1982),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2000),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1988),
.B(n_1952),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1997),
.B(n_1962),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2006),
.B(n_1964),
.Y(n_2041)
);

INVxp67_ASAP7_75t_L g2042 ( 
.A(n_1992),
.Y(n_2042)
);

INVx1_ASAP7_75t_SL g2043 ( 
.A(n_2004),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1990),
.B(n_1962),
.Y(n_2044)
);

INVxp67_ASAP7_75t_SL g2045 ( 
.A(n_1992),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2000),
.B(n_1965),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1980),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1980),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_2019),
.B(n_1943),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1983),
.B(n_1960),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2009),
.B(n_1964),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2009),
.B(n_1964),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2011),
.B(n_1965),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_1990),
.B(n_1966),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2009),
.B(n_1970),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1987),
.B(n_1970),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_1984),
.B(n_1966),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1987),
.B(n_1994),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1994),
.B(n_1970),
.Y(n_2059)
);

HB1xp67_ASAP7_75t_L g2060 ( 
.A(n_1981),
.Y(n_2060)
);

NAND2x1_ASAP7_75t_L g2061 ( 
.A(n_1983),
.B(n_1921),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1981),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2001),
.B(n_1971),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_1985),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_1984),
.B(n_1975),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1986),
.B(n_1973),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1986),
.B(n_1974),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2001),
.B(n_1971),
.Y(n_2068)
);

A2O1A1Ixp33_ASAP7_75t_L g2069 ( 
.A1(n_2033),
.A2(n_1898),
.B(n_1947),
.C(n_1935),
.Y(n_2069)
);

AOI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_2030),
.A2(n_1887),
.B1(n_1908),
.B2(n_1902),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2043),
.B(n_2004),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2043),
.B(n_1985),
.Y(n_2072)
);

OAI211xp5_ASAP7_75t_L g2073 ( 
.A1(n_2037),
.A2(n_1995),
.B(n_1979),
.C(n_2020),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2060),
.Y(n_2074)
);

AOI322xp5_ASAP7_75t_L g2075 ( 
.A1(n_2034),
.A2(n_1944),
.A3(n_1943),
.B1(n_1902),
.B2(n_1998),
.C1(n_2014),
.C2(n_2019),
.Y(n_2075)
);

OAI211xp5_ASAP7_75t_L g2076 ( 
.A1(n_2037),
.A2(n_1995),
.B(n_1979),
.C(n_2020),
.Y(n_2076)
);

AOI22xp33_ASAP7_75t_L g2077 ( 
.A1(n_2034),
.A2(n_2013),
.B1(n_1896),
.B2(n_1909),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2060),
.Y(n_2078)
);

AOI321xp33_ASAP7_75t_L g2079 ( 
.A1(n_2045),
.A2(n_1907),
.A3(n_1977),
.B1(n_1998),
.B2(n_2021),
.C(n_2007),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_2030),
.A2(n_1896),
.B1(n_2013),
.B2(n_1924),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2042),
.B(n_2021),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2047),
.Y(n_2082)
);

AOI221xp5_ASAP7_75t_L g2083 ( 
.A1(n_2033),
.A2(n_1977),
.B1(n_2005),
.B2(n_1999),
.C(n_1944),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2047),
.Y(n_2084)
);

AOI221xp5_ASAP7_75t_L g2085 ( 
.A1(n_2045),
.A2(n_2005),
.B1(n_1999),
.B2(n_1943),
.C(n_1944),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2048),
.Y(n_2086)
);

AOI211x1_ASAP7_75t_L g2087 ( 
.A1(n_2050),
.A2(n_2053),
.B(n_2058),
.C(n_2036),
.Y(n_2087)
);

OAI322xp33_ASAP7_75t_L g2088 ( 
.A1(n_2042),
.A2(n_2013),
.A3(n_2002),
.B1(n_1886),
.B2(n_1911),
.C1(n_2023),
.C2(n_2028),
.Y(n_2088)
);

NAND2x1p5_ASAP7_75t_L g2089 ( 
.A(n_2061),
.B(n_1995),
.Y(n_2089)
);

OAI21xp5_ASAP7_75t_L g2090 ( 
.A1(n_2053),
.A2(n_1957),
.B(n_1979),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2035),
.Y(n_2091)
);

INVx1_ASAP7_75t_SL g2092 ( 
.A(n_2032),
.Y(n_2092)
);

OAI221xp5_ASAP7_75t_SL g2093 ( 
.A1(n_2032),
.A2(n_1998),
.B1(n_2014),
.B2(n_1945),
.C(n_1924),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2048),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2062),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2062),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_SL g2097 ( 
.A1(n_2029),
.A2(n_1945),
.B1(n_1995),
.B2(n_1779),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2035),
.A2(n_1896),
.B1(n_1989),
.B2(n_1915),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2082),
.Y(n_2099)
);

O2A1O1Ixp33_ASAP7_75t_SL g2100 ( 
.A1(n_2073),
.A2(n_2064),
.B(n_2061),
.C(n_2038),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2084),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2070),
.A2(n_2077),
.B1(n_2069),
.B2(n_2080),
.Y(n_2102)
);

INVx1_ASAP7_75t_SL g2103 ( 
.A(n_2092),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2086),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_2091),
.Y(n_2105)
);

AOI322xp5_ASAP7_75t_L g2106 ( 
.A1(n_2077),
.A2(n_2036),
.A3(n_2049),
.B1(n_2029),
.B2(n_2031),
.C1(n_2064),
.C2(n_2041),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2094),
.Y(n_2107)
);

NAND2xp33_ASAP7_75t_SL g2108 ( 
.A(n_2071),
.B(n_2058),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2095),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2096),
.Y(n_2110)
);

NOR3xp33_ASAP7_75t_L g2111 ( 
.A(n_2069),
.B(n_2038),
.C(n_2046),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2081),
.B(n_2049),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2074),
.Y(n_2113)
);

OAI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2093),
.A2(n_1989),
.B1(n_2049),
.B2(n_2041),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2078),
.Y(n_2115)
);

AOI221xp5_ASAP7_75t_L g2116 ( 
.A1(n_2088),
.A2(n_2054),
.B1(n_2044),
.B2(n_2031),
.C(n_2040),
.Y(n_2116)
);

INVx1_ASAP7_75t_SL g2117 ( 
.A(n_2072),
.Y(n_2117)
);

OAI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_2093),
.A2(n_2087),
.B1(n_2076),
.B2(n_2098),
.Y(n_2118)
);

NAND3xp33_ASAP7_75t_SL g2119 ( 
.A(n_2079),
.B(n_2052),
.C(n_2051),
.Y(n_2119)
);

INVxp33_ASAP7_75t_L g2120 ( 
.A(n_2089),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2075),
.B(n_2056),
.Y(n_2121)
);

AOI221xp5_ASAP7_75t_SL g2122 ( 
.A1(n_2118),
.A2(n_2083),
.B1(n_2085),
.B2(n_2090),
.C(n_2046),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2105),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2103),
.B(n_2056),
.Y(n_2124)
);

AOI211xp5_ASAP7_75t_L g2125 ( 
.A1(n_2111),
.A2(n_2040),
.B(n_2054),
.C(n_2044),
.Y(n_2125)
);

AOI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_2100),
.A2(n_2089),
.B(n_2067),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_2117),
.B(n_2051),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2113),
.Y(n_2128)
);

OAI21xp33_ASAP7_75t_L g2129 ( 
.A1(n_2111),
.A2(n_2059),
.B(n_2055),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2099),
.Y(n_2130)
);

AOI222xp33_ASAP7_75t_L g2131 ( 
.A1(n_2121),
.A2(n_2119),
.B1(n_2116),
.B2(n_2102),
.C1(n_2114),
.C2(n_2108),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2101),
.Y(n_2132)
);

AOI22xp33_ASAP7_75t_L g2133 ( 
.A1(n_2112),
.A2(n_1896),
.B1(n_2031),
.B2(n_2007),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2104),
.Y(n_2134)
);

NOR2x1_ASAP7_75t_L g2135 ( 
.A(n_2123),
.B(n_2115),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2124),
.B(n_2127),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2124),
.B(n_2106),
.Y(n_2137)
);

NAND4xp25_ASAP7_75t_L g2138 ( 
.A(n_2131),
.B(n_2100),
.C(n_2110),
.D(n_2109),
.Y(n_2138)
);

NAND3xp33_ASAP7_75t_SL g2139 ( 
.A(n_2126),
.B(n_2120),
.C(n_2107),
.Y(n_2139)
);

OAI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_2122),
.A2(n_2120),
.B(n_2097),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_2125),
.B(n_2052),
.Y(n_2141)
);

NOR2x1_ASAP7_75t_L g2142 ( 
.A(n_2123),
.B(n_2055),
.Y(n_2142)
);

NOR3xp33_ASAP7_75t_L g2143 ( 
.A(n_2128),
.B(n_2065),
.C(n_2057),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2129),
.B(n_2059),
.Y(n_2144)
);

INVxp33_ASAP7_75t_L g2145 ( 
.A(n_2128),
.Y(n_2145)
);

NAND4xp25_ASAP7_75t_L g2146 ( 
.A(n_2132),
.B(n_2134),
.C(n_2130),
.D(n_2133),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2134),
.B(n_2039),
.Y(n_2147)
);

OAI211xp5_ASAP7_75t_SL g2148 ( 
.A1(n_2140),
.A2(n_2130),
.B(n_2039),
.C(n_2057),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2143),
.B(n_2063),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2142),
.B(n_2063),
.Y(n_2150)
);

OAI221xp5_ASAP7_75t_L g2151 ( 
.A1(n_2137),
.A2(n_2065),
.B1(n_1989),
.B2(n_2002),
.C(n_2067),
.Y(n_2151)
);

AOI222xp33_ASAP7_75t_L g2152 ( 
.A1(n_2139),
.A2(n_1996),
.B1(n_2007),
.B2(n_2003),
.C1(n_2027),
.C2(n_1926),
.Y(n_2152)
);

OAI211xp5_ASAP7_75t_L g2153 ( 
.A1(n_2138),
.A2(n_2068),
.B(n_2022),
.C(n_2066),
.Y(n_2153)
);

AOI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_2145),
.A2(n_1926),
.B1(n_1918),
.B2(n_1929),
.Y(n_2154)
);

NAND3xp33_ASAP7_75t_SL g2155 ( 
.A(n_2150),
.B(n_2136),
.C(n_2147),
.Y(n_2155)
);

OAI31xp33_ASAP7_75t_L g2156 ( 
.A1(n_2148),
.A2(n_2146),
.A3(n_2141),
.B(n_2144),
.Y(n_2156)
);

OAI221xp5_ASAP7_75t_L g2157 ( 
.A1(n_2151),
.A2(n_2135),
.B1(n_2066),
.B2(n_2023),
.C(n_2028),
.Y(n_2157)
);

OAI21xp5_ASAP7_75t_L g2158 ( 
.A1(n_2149),
.A2(n_2068),
.B(n_1993),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2153),
.Y(n_2159)
);

OAI21xp33_ASAP7_75t_SL g2160 ( 
.A1(n_2152),
.A2(n_1993),
.B(n_1991),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2154),
.B(n_2024),
.Y(n_2161)
);

AOI221xp5_ASAP7_75t_L g2162 ( 
.A1(n_2148),
.A2(n_1996),
.B1(n_2003),
.B2(n_2027),
.C(n_1926),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_2155),
.A2(n_1978),
.B1(n_2022),
.B2(n_1991),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_2159),
.A2(n_2160),
.B1(n_2161),
.B2(n_2157),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2158),
.Y(n_2165)
);

NAND4xp75_ASAP7_75t_L g2166 ( 
.A(n_2156),
.B(n_1991),
.C(n_1993),
.D(n_1672),
.Y(n_2166)
);

NAND4xp75_ASAP7_75t_L g2167 ( 
.A(n_2162),
.B(n_1672),
.C(n_1945),
.D(n_2024),
.Y(n_2167)
);

AOI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2155),
.A2(n_1978),
.B1(n_1929),
.B2(n_1918),
.Y(n_2168)
);

NOR2x1_ASAP7_75t_L g2169 ( 
.A(n_2155),
.B(n_1978),
.Y(n_2169)
);

AOI22xp5_ASAP7_75t_L g2170 ( 
.A1(n_2164),
.A2(n_1978),
.B1(n_2003),
.B2(n_1996),
.Y(n_2170)
);

OAI221xp5_ASAP7_75t_L g2171 ( 
.A1(n_2168),
.A2(n_2027),
.B1(n_2018),
.B2(n_2026),
.C(n_2017),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_2169),
.B(n_1950),
.Y(n_2172)
);

OAI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_2166),
.A2(n_2165),
.B(n_2167),
.Y(n_2173)
);

OAI21xp5_ASAP7_75t_SL g2174 ( 
.A1(n_2163),
.A2(n_1779),
.B(n_1950),
.Y(n_2174)
);

NOR4xp25_ASAP7_75t_L g2175 ( 
.A(n_2173),
.B(n_2171),
.C(n_2174),
.D(n_2170),
.Y(n_2175)
);

AOI22xp33_ASAP7_75t_SL g2176 ( 
.A1(n_2172),
.A2(n_1785),
.B1(n_1929),
.B2(n_1918),
.Y(n_2176)
);

AO22x2_ASAP7_75t_L g2177 ( 
.A1(n_2175),
.A2(n_2026),
.B1(n_2008),
.B2(n_2017),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2177),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2177),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2179),
.A2(n_2176),
.B1(n_2010),
.B2(n_2016),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2178),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2180),
.Y(n_2182)
);

OAI21xp5_ASAP7_75t_L g2183 ( 
.A1(n_2181),
.A2(n_2018),
.B(n_2010),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_SL g2184 ( 
.A(n_2182),
.B(n_2008),
.Y(n_2184)
);

AO21x2_ASAP7_75t_L g2185 ( 
.A1(n_2184),
.A2(n_2183),
.B(n_2016),
.Y(n_2185)
);

XNOR2xp5_ASAP7_75t_L g2186 ( 
.A(n_2185),
.B(n_1814),
.Y(n_2186)
);

AOI221xp5_ASAP7_75t_L g2187 ( 
.A1(n_2186),
.A2(n_2015),
.B1(n_1886),
.B2(n_1950),
.C(n_1967),
.Y(n_2187)
);

AOI211xp5_ASAP7_75t_L g2188 ( 
.A1(n_2187),
.A2(n_2015),
.B(n_1925),
.C(n_1967),
.Y(n_2188)
);


endmodule