module fake_ibex_866_n_7605 (n_904, n_179, n_1086, n_564, n_737, n_120, n_1100, n_999, n_48, n_1037, n_560, n_40, n_1104, n_597, n_622, n_811, n_1098, n_412, n_939, n_689, n_1123, n_536, n_325, n_662, n_781, n_1012, n_598, n_698, n_732, n_973, n_1031, n_1034, n_113, n_1115, n_1113, n_290, n_215, n_477, n_826, n_388, n_221, n_26, n_567, n_827, n_178, n_875, n_497, n_282, n_55, n_679, n_810, n_277, n_723, n_982, n_424, n_541, n_976, n_588, n_683, n_170, n_962, n_555, n_758, n_1042, n_1066, n_663, n_859, n_1043, n_575, n_767, n_454, n_367, n_1118, n_29, n_650, n_1056, n_2, n_320, n_707, n_470, n_1111, n_533, n_593, n_395, n_699, n_262, n_1024, n_181, n_888, n_729, n_1008, n_861, n_368, n_1069, n_483, n_1063, n_753, n_161, n_508, n_625, n_415, n_24, n_239, n_585, n_631, n_971, n_1053, n_1, n_233, n_500, n_1016, n_311, n_563, n_626, n_291, n_371, n_843, n_1027, n_552, n_100, n_220, n_579, n_673, n_110, n_881, n_935, n_829, n_869, n_799, n_1007, n_496, n_331, n_793, n_891, n_1083, n_279, n_981, n_125, n_381, n_658, n_858, n_231, n_1085, n_775, n_608, n_710, n_154, n_251, n_206, n_983, n_460, n_1038, n_1124, n_352, n_343, n_950, n_590, n_965, n_997, n_551, n_436, n_833, n_911, n_784, n_64, n_418, n_724, n_762, n_445, n_348, n_131, n_527, n_540, n_908, n_561, n_545, n_850, n_19, n_715, n_202, n_751, n_614, n_535, n_709, n_237, n_628, n_823, n_1046, n_696, n_704, n_39, n_130, n_792, n_862, n_900, n_1084, n_708, n_63, n_592, n_1089, n_189, n_38, n_380, n_576, n_736, n_895, n_15, n_339, n_84, n_183, n_703, n_20, n_335, n_518, n_640, n_68, n_80, n_865, n_928, n_596, n_693, n_507, n_898, n_624, n_953, n_991, n_37, n_75, n_107, n_482, n_119, n_133, n_356, n_333, n_472, n_595, n_745, n_387, n_91, n_538, n_1058, n_187, n_307, n_135, n_317, n_800, n_952, n_305, n_925, n_682, n_139, n_390, n_481, n_157, n_1090, n_410, n_491, n_980, n_1078, n_448, n_582, n_57, n_149, n_253, n_550, n_828, n_584, n_342, n_602, n_749, n_818, n_532, n_813, n_394, n_163, n_162, n_209, n_401, n_630, n_883, n_502, n_398, n_442, n_890, n_116, n_1035, n_816, n_366, n_534, n_905, n_543, n_944, n_559, n_515, n_954, n_386, n_548, n_95, n_200, n_747, n_766, n_989, n_984, n_1054, n_1065, n_167, n_948, n_396, n_750, n_322, n_743, n_610, n_903, n_773, n_441, n_717, n_529, n_361, n_318, n_855, n_910, n_456, n_728, n_79, n_10, n_641, n_1057, n_152, n_88, n_1029, n_160, n_927, n_433, n_229, n_480, n_657, n_666, n_798, n_603, n_138, n_417, n_192, n_420, n_1079, n_1004, n_840, n_272, n_473, n_684, n_772, n_853, n_164, n_403, n_490, n_785, n_933, n_241, n_414, n_228, n_504, n_190, n_661, n_727, n_198, n_169, n_655, n_791, n_967, n_876, n_644, n_310, n_5, n_122, n_701, n_825, n_916, n_646, n_730, n_344, n_615, n_719, n_72, n_558, n_616, n_674, n_224, n_1075, n_102, n_243, n_992, n_400, n_821, n_1064, n_369, n_62, n_421, n_947, n_392, n_951, n_1080, n_197, n_232, n_104, n_213, n_428, n_172, n_194, n_76, n_294, n_848, n_587, n_438, n_804, n_986, n_118, n_166, n_812, n_882, n_1097, n_713, n_432, n_146, n_247, n_795, n_912, n_1039, n_901, n_376, n_451, n_868, n_411, n_523, n_955, n_283, n_637, n_83, n_499, n_226, n_45, n_405, n_36, n_365, n_528, n_820, n_542, n_721, n_712, n_359, n_1048, n_260, n_573, n_128, n_830, n_943, n_776, n_115, n_106, n_327, n_245, n_32, n_796, n_556, n_150, n_236, n_664, n_788, n_4, n_81, n_921, n_300, n_651, n_618, n_16, n_458, n_690, n_329, n_814, n_6, n_147, n_457, n_93, n_675, n_734, n_121, n_140, n_742, n_759, n_893, n_338, n_332, n_605, n_1018, n_1015, n_570, n_142, n_429, n_539, n_49, n_252, n_839, n_894, n_580, n_255, n_234, n_304, n_488, n_731, n_1099, n_902, n_303, n_1110, n_274, n_671, n_7, n_475, n_520, n_256, n_312, n_466, n_1023, n_836, n_461, n_1105, n_936, n_887, n_831, n_807, n_308, n_354, n_464, n_134, n_270, n_1101, n_1021, n_937, n_970, n_212, n_180, n_292, n_854, n_553, n_375, n_738, n_35, n_845, n_695, n_184, n_676, n_562, n_218, n_316, n_498, n_56, n_643, n_1120, n_996, n_397, n_771, n_101, n_722, n_815, n_613, n_977, n_21, n_379, n_281, n_514, n_219, n_711, n_50, n_897, n_459, n_678, n_680, n_1055, n_416, n_42, n_1014, n_754, n_566, n_607, n_993, n_112, n_806, n_156, n_922, n_957, n_1045, n_86, n_382, n_1010, n_47, n_1122, n_565, n_67, n_633, n_357, n_434, n_941, n_216, n_1088, n_748, n_82, n_204, n_639, n_223, n_909, n_298, n_87, n_757, n_492, n_857, n_171, n_265, n_439, n_103, n_96, n_27, n_647, n_978, n_1096, n_33, n_987, n_756, n_301, n_309, n_513, n_452, n_468, n_768, n_22, n_314, n_1009, n_501, n_778, n_966, n_782, n_254, n_660, n_258, n_196, n_606, n_1030, n_1082, n_1067, n_746, n_340, n_779, n_225, n_884, n_958, n_266, n_74, n_288, n_173, n_185, n_505, n_735, n_822, n_1112, n_467, n_870, n_315, n_31, n_516, n_422, n_503, n_687, n_153, n_817, n_852, n_969, n_1036, n_177, n_511, n_617, n_659, n_509, n_512, n_702, n_867, n_968, n_264, n_151, n_443, n_733, n_1000, n_287, n_246, n_634, n_787, n_453, n_645, n_923, n_574, n_129, n_959, n_694, n_1062, n_132, n_886, n_469, n_90, n_364, n_985, n_426, n_276, n_127, n_249, n_521, n_519, n_52, n_990, n_399, n_763, n_847, n_878, n_547, n_718, n_794, n_665, n_601, n_1059, n_609, n_964, n_273, n_111, n_319, n_321, n_244, n_783, n_809, n_524, n_856, n_926, n_360, n_44, n_94, n_168, n_589, n_60, n_182, n_549, n_280, n_358, n_370, n_688, n_78, n_69, n_714, n_780, n_838, n_960, n_97, n_261, n_355, n_437, n_571, n_510, n_544, n_841, n_700, n_846, n_945, n_837, n_716, n_769, n_636, n_284, n_988, n_143, n_1025, n_885, n_413, n_51, n_835, n_871, n_208, n_402, n_726, n_449, n_594, n_455, n_423, n_669, n_569, n_350, n_790, n_341, n_849, n_73, n_17, n_803, n_210, n_872, n_940, n_175, n_979, n_485, n_92, n_336, n_599, n_1106, n_278, n_230, n_3, n_108, n_440, n_419, n_638, n_65, n_85, n_377, n_145, n_740, n_656, n_478, n_257, n_248, n_789, n_1044, n_877, n_808, n_1001, n_61, n_677, n_450, n_1005, n_144, n_1050, n_672, n_53, n_972, n_1041, n_383, n_1070, n_1109, n_938, n_956, n_30, n_620, n_238, n_1093, n_12, n_864, n_654, n_1121, n_89, n_54, n_1081, n_1061, n_1087, n_158, n_755, n_517, n_546, n_1091, n_8, n_324, n_299, n_374, n_526, n_578, n_896, n_302, n_1092, n_1119, n_109, n_525, n_1076, n_915, n_296, n_583, n_924, n_59, n_46, n_123, n_11, n_572, n_917, n_188, n_347, n_363, n_653, n_201, n_691, n_819, n_946, n_462, n_629, n_961, n_1068, n_275, n_330, n_444, n_802, n_774, n_323, n_1095, n_621, n_407, n_117, n_242, n_447, n_604, n_34, n_293, n_879, n_1028, n_801, n_899, n_851, n_203, n_1032, n_522, n_1017, n_25, n_913, n_866, n_99, n_227, n_431, n_124, n_632, n_425, n_136, n_530, n_554, n_725, n_577, n_66, n_28, n_934, n_77, n_408, n_1103, n_176, n_126, n_471, n_744, n_844, n_919, n_995, n_465, n_1073, n_71, n_685, n_313, n_765, n_619, n_686, n_770, n_148, n_353, n_537, n_385, n_285, n_435, n_141, n_860, n_932, n_1102, n_1071, n_1107, n_705, n_586, n_760, n_191, n_207, n_842, n_268, n_761, n_326, n_777, n_155, n_493, n_222, n_41, n_351, n_0, n_1060, n_476, n_174, n_1033, n_892, n_531, n_235, n_479, n_474, n_557, n_600, n_975, n_649, n_58, n_974, n_1006, n_263, n_834, n_1074, n_963, n_874, n_1116, n_486, n_463, n_697, n_907, n_998, n_752, n_487, n_214, n_345, n_918, n_1022, n_668, n_193, n_739, n_391, n_337, n_1077, n_797, n_931, n_18, n_211, n_306, n_240, n_623, n_949, n_205, n_373, n_1020, n_930, n_114, n_267, n_427, n_741, n_863, n_1013, n_873, n_297, n_764, n_409, n_70, n_289, n_195, n_914, n_384, n_98, n_1047, n_259, n_269, n_349, n_159, n_805, n_929, n_652, n_43, n_14, n_165, n_372, n_13, n_430, n_1011, n_1094, n_994, n_1052, n_9, n_217, n_484, n_489, n_627, n_648, n_1003, n_495, n_137, n_346, n_286, n_611, n_612, n_706, n_1019, n_681, n_378, n_186, n_271, n_942, n_667, n_199, n_1026, n_824, n_334, n_906, n_1040, n_250, n_670, n_786, n_1049, n_446, n_494, n_642, n_591, n_1117, n_692, n_635, n_889, n_506, n_568, n_1114, n_1072, n_406, n_105, n_1002, n_404, n_1108, n_920, n_362, n_23, n_389, n_295, n_581, n_393, n_880, n_1051, n_832, n_720, n_328, n_7605);

input n_904;
input n_179;
input n_1086;
input n_564;
input n_737;
input n_120;
input n_1100;
input n_999;
input n_48;
input n_1037;
input n_560;
input n_40;
input n_1104;
input n_597;
input n_622;
input n_811;
input n_1098;
input n_412;
input n_939;
input n_689;
input n_1123;
input n_536;
input n_325;
input n_662;
input n_781;
input n_1012;
input n_598;
input n_698;
input n_732;
input n_973;
input n_1031;
input n_1034;
input n_113;
input n_1115;
input n_1113;
input n_290;
input n_215;
input n_477;
input n_826;
input n_388;
input n_221;
input n_26;
input n_567;
input n_827;
input n_178;
input n_875;
input n_497;
input n_282;
input n_55;
input n_679;
input n_810;
input n_277;
input n_723;
input n_982;
input n_424;
input n_541;
input n_976;
input n_588;
input n_683;
input n_170;
input n_962;
input n_555;
input n_758;
input n_1042;
input n_1066;
input n_663;
input n_859;
input n_1043;
input n_575;
input n_767;
input n_454;
input n_367;
input n_1118;
input n_29;
input n_650;
input n_1056;
input n_2;
input n_320;
input n_707;
input n_470;
input n_1111;
input n_533;
input n_593;
input n_395;
input n_699;
input n_262;
input n_1024;
input n_181;
input n_888;
input n_729;
input n_1008;
input n_861;
input n_368;
input n_1069;
input n_483;
input n_1063;
input n_753;
input n_161;
input n_508;
input n_625;
input n_415;
input n_24;
input n_239;
input n_585;
input n_631;
input n_971;
input n_1053;
input n_1;
input n_233;
input n_500;
input n_1016;
input n_311;
input n_563;
input n_626;
input n_291;
input n_371;
input n_843;
input n_1027;
input n_552;
input n_100;
input n_220;
input n_579;
input n_673;
input n_110;
input n_881;
input n_935;
input n_829;
input n_869;
input n_799;
input n_1007;
input n_496;
input n_331;
input n_793;
input n_891;
input n_1083;
input n_279;
input n_981;
input n_125;
input n_381;
input n_658;
input n_858;
input n_231;
input n_1085;
input n_775;
input n_608;
input n_710;
input n_154;
input n_251;
input n_206;
input n_983;
input n_460;
input n_1038;
input n_1124;
input n_352;
input n_343;
input n_950;
input n_590;
input n_965;
input n_997;
input n_551;
input n_436;
input n_833;
input n_911;
input n_784;
input n_64;
input n_418;
input n_724;
input n_762;
input n_445;
input n_348;
input n_131;
input n_527;
input n_540;
input n_908;
input n_561;
input n_545;
input n_850;
input n_19;
input n_715;
input n_202;
input n_751;
input n_614;
input n_535;
input n_709;
input n_237;
input n_628;
input n_823;
input n_1046;
input n_696;
input n_704;
input n_39;
input n_130;
input n_792;
input n_862;
input n_900;
input n_1084;
input n_708;
input n_63;
input n_592;
input n_1089;
input n_189;
input n_38;
input n_380;
input n_576;
input n_736;
input n_895;
input n_15;
input n_339;
input n_84;
input n_183;
input n_703;
input n_20;
input n_335;
input n_518;
input n_640;
input n_68;
input n_80;
input n_865;
input n_928;
input n_596;
input n_693;
input n_507;
input n_898;
input n_624;
input n_953;
input n_991;
input n_37;
input n_75;
input n_107;
input n_482;
input n_119;
input n_133;
input n_356;
input n_333;
input n_472;
input n_595;
input n_745;
input n_387;
input n_91;
input n_538;
input n_1058;
input n_187;
input n_307;
input n_135;
input n_317;
input n_800;
input n_952;
input n_305;
input n_925;
input n_682;
input n_139;
input n_390;
input n_481;
input n_157;
input n_1090;
input n_410;
input n_491;
input n_980;
input n_1078;
input n_448;
input n_582;
input n_57;
input n_149;
input n_253;
input n_550;
input n_828;
input n_584;
input n_342;
input n_602;
input n_749;
input n_818;
input n_532;
input n_813;
input n_394;
input n_163;
input n_162;
input n_209;
input n_401;
input n_630;
input n_883;
input n_502;
input n_398;
input n_442;
input n_890;
input n_116;
input n_1035;
input n_816;
input n_366;
input n_534;
input n_905;
input n_543;
input n_944;
input n_559;
input n_515;
input n_954;
input n_386;
input n_548;
input n_95;
input n_200;
input n_747;
input n_766;
input n_989;
input n_984;
input n_1054;
input n_1065;
input n_167;
input n_948;
input n_396;
input n_750;
input n_322;
input n_743;
input n_610;
input n_903;
input n_773;
input n_441;
input n_717;
input n_529;
input n_361;
input n_318;
input n_855;
input n_910;
input n_456;
input n_728;
input n_79;
input n_10;
input n_641;
input n_1057;
input n_152;
input n_88;
input n_1029;
input n_160;
input n_927;
input n_433;
input n_229;
input n_480;
input n_657;
input n_666;
input n_798;
input n_603;
input n_138;
input n_417;
input n_192;
input n_420;
input n_1079;
input n_1004;
input n_840;
input n_272;
input n_473;
input n_684;
input n_772;
input n_853;
input n_164;
input n_403;
input n_490;
input n_785;
input n_933;
input n_241;
input n_414;
input n_228;
input n_504;
input n_190;
input n_661;
input n_727;
input n_198;
input n_169;
input n_655;
input n_791;
input n_967;
input n_876;
input n_644;
input n_310;
input n_5;
input n_122;
input n_701;
input n_825;
input n_916;
input n_646;
input n_730;
input n_344;
input n_615;
input n_719;
input n_72;
input n_558;
input n_616;
input n_674;
input n_224;
input n_1075;
input n_102;
input n_243;
input n_992;
input n_400;
input n_821;
input n_1064;
input n_369;
input n_62;
input n_421;
input n_947;
input n_392;
input n_951;
input n_1080;
input n_197;
input n_232;
input n_104;
input n_213;
input n_428;
input n_172;
input n_194;
input n_76;
input n_294;
input n_848;
input n_587;
input n_438;
input n_804;
input n_986;
input n_118;
input n_166;
input n_812;
input n_882;
input n_1097;
input n_713;
input n_432;
input n_146;
input n_247;
input n_795;
input n_912;
input n_1039;
input n_901;
input n_376;
input n_451;
input n_868;
input n_411;
input n_523;
input n_955;
input n_283;
input n_637;
input n_83;
input n_499;
input n_226;
input n_45;
input n_405;
input n_36;
input n_365;
input n_528;
input n_820;
input n_542;
input n_721;
input n_712;
input n_359;
input n_1048;
input n_260;
input n_573;
input n_128;
input n_830;
input n_943;
input n_776;
input n_115;
input n_106;
input n_327;
input n_245;
input n_32;
input n_796;
input n_556;
input n_150;
input n_236;
input n_664;
input n_788;
input n_4;
input n_81;
input n_921;
input n_300;
input n_651;
input n_618;
input n_16;
input n_458;
input n_690;
input n_329;
input n_814;
input n_6;
input n_147;
input n_457;
input n_93;
input n_675;
input n_734;
input n_121;
input n_140;
input n_742;
input n_759;
input n_893;
input n_338;
input n_332;
input n_605;
input n_1018;
input n_1015;
input n_570;
input n_142;
input n_429;
input n_539;
input n_49;
input n_252;
input n_839;
input n_894;
input n_580;
input n_255;
input n_234;
input n_304;
input n_488;
input n_731;
input n_1099;
input n_902;
input n_303;
input n_1110;
input n_274;
input n_671;
input n_7;
input n_475;
input n_520;
input n_256;
input n_312;
input n_466;
input n_1023;
input n_836;
input n_461;
input n_1105;
input n_936;
input n_887;
input n_831;
input n_807;
input n_308;
input n_354;
input n_464;
input n_134;
input n_270;
input n_1101;
input n_1021;
input n_937;
input n_970;
input n_212;
input n_180;
input n_292;
input n_854;
input n_553;
input n_375;
input n_738;
input n_35;
input n_845;
input n_695;
input n_184;
input n_676;
input n_562;
input n_218;
input n_316;
input n_498;
input n_56;
input n_643;
input n_1120;
input n_996;
input n_397;
input n_771;
input n_101;
input n_722;
input n_815;
input n_613;
input n_977;
input n_21;
input n_379;
input n_281;
input n_514;
input n_219;
input n_711;
input n_50;
input n_897;
input n_459;
input n_678;
input n_680;
input n_1055;
input n_416;
input n_42;
input n_1014;
input n_754;
input n_566;
input n_607;
input n_993;
input n_112;
input n_806;
input n_156;
input n_922;
input n_957;
input n_1045;
input n_86;
input n_382;
input n_1010;
input n_47;
input n_1122;
input n_565;
input n_67;
input n_633;
input n_357;
input n_434;
input n_941;
input n_216;
input n_1088;
input n_748;
input n_82;
input n_204;
input n_639;
input n_223;
input n_909;
input n_298;
input n_87;
input n_757;
input n_492;
input n_857;
input n_171;
input n_265;
input n_439;
input n_103;
input n_96;
input n_27;
input n_647;
input n_978;
input n_1096;
input n_33;
input n_987;
input n_756;
input n_301;
input n_309;
input n_513;
input n_452;
input n_468;
input n_768;
input n_22;
input n_314;
input n_1009;
input n_501;
input n_778;
input n_966;
input n_782;
input n_254;
input n_660;
input n_258;
input n_196;
input n_606;
input n_1030;
input n_1082;
input n_1067;
input n_746;
input n_340;
input n_779;
input n_225;
input n_884;
input n_958;
input n_266;
input n_74;
input n_288;
input n_173;
input n_185;
input n_505;
input n_735;
input n_822;
input n_1112;
input n_467;
input n_870;
input n_315;
input n_31;
input n_516;
input n_422;
input n_503;
input n_687;
input n_153;
input n_817;
input n_852;
input n_969;
input n_1036;
input n_177;
input n_511;
input n_617;
input n_659;
input n_509;
input n_512;
input n_702;
input n_867;
input n_968;
input n_264;
input n_151;
input n_443;
input n_733;
input n_1000;
input n_287;
input n_246;
input n_634;
input n_787;
input n_453;
input n_645;
input n_923;
input n_574;
input n_129;
input n_959;
input n_694;
input n_1062;
input n_132;
input n_886;
input n_469;
input n_90;
input n_364;
input n_985;
input n_426;
input n_276;
input n_127;
input n_249;
input n_521;
input n_519;
input n_52;
input n_990;
input n_399;
input n_763;
input n_847;
input n_878;
input n_547;
input n_718;
input n_794;
input n_665;
input n_601;
input n_1059;
input n_609;
input n_964;
input n_273;
input n_111;
input n_319;
input n_321;
input n_244;
input n_783;
input n_809;
input n_524;
input n_856;
input n_926;
input n_360;
input n_44;
input n_94;
input n_168;
input n_589;
input n_60;
input n_182;
input n_549;
input n_280;
input n_358;
input n_370;
input n_688;
input n_78;
input n_69;
input n_714;
input n_780;
input n_838;
input n_960;
input n_97;
input n_261;
input n_355;
input n_437;
input n_571;
input n_510;
input n_544;
input n_841;
input n_700;
input n_846;
input n_945;
input n_837;
input n_716;
input n_769;
input n_636;
input n_284;
input n_988;
input n_143;
input n_1025;
input n_885;
input n_413;
input n_51;
input n_835;
input n_871;
input n_208;
input n_402;
input n_726;
input n_449;
input n_594;
input n_455;
input n_423;
input n_669;
input n_569;
input n_350;
input n_790;
input n_341;
input n_849;
input n_73;
input n_17;
input n_803;
input n_210;
input n_872;
input n_940;
input n_175;
input n_979;
input n_485;
input n_92;
input n_336;
input n_599;
input n_1106;
input n_278;
input n_230;
input n_3;
input n_108;
input n_440;
input n_419;
input n_638;
input n_65;
input n_85;
input n_377;
input n_145;
input n_740;
input n_656;
input n_478;
input n_257;
input n_248;
input n_789;
input n_1044;
input n_877;
input n_808;
input n_1001;
input n_61;
input n_677;
input n_450;
input n_1005;
input n_144;
input n_1050;
input n_672;
input n_53;
input n_972;
input n_1041;
input n_383;
input n_1070;
input n_1109;
input n_938;
input n_956;
input n_30;
input n_620;
input n_238;
input n_1093;
input n_12;
input n_864;
input n_654;
input n_1121;
input n_89;
input n_54;
input n_1081;
input n_1061;
input n_1087;
input n_158;
input n_755;
input n_517;
input n_546;
input n_1091;
input n_8;
input n_324;
input n_299;
input n_374;
input n_526;
input n_578;
input n_896;
input n_302;
input n_1092;
input n_1119;
input n_109;
input n_525;
input n_1076;
input n_915;
input n_296;
input n_583;
input n_924;
input n_59;
input n_46;
input n_123;
input n_11;
input n_572;
input n_917;
input n_188;
input n_347;
input n_363;
input n_653;
input n_201;
input n_691;
input n_819;
input n_946;
input n_462;
input n_629;
input n_961;
input n_1068;
input n_275;
input n_330;
input n_444;
input n_802;
input n_774;
input n_323;
input n_1095;
input n_621;
input n_407;
input n_117;
input n_242;
input n_447;
input n_604;
input n_34;
input n_293;
input n_879;
input n_1028;
input n_801;
input n_899;
input n_851;
input n_203;
input n_1032;
input n_522;
input n_1017;
input n_25;
input n_913;
input n_866;
input n_99;
input n_227;
input n_431;
input n_124;
input n_632;
input n_425;
input n_136;
input n_530;
input n_554;
input n_725;
input n_577;
input n_66;
input n_28;
input n_934;
input n_77;
input n_408;
input n_1103;
input n_176;
input n_126;
input n_471;
input n_744;
input n_844;
input n_919;
input n_995;
input n_465;
input n_1073;
input n_71;
input n_685;
input n_313;
input n_765;
input n_619;
input n_686;
input n_770;
input n_148;
input n_353;
input n_537;
input n_385;
input n_285;
input n_435;
input n_141;
input n_860;
input n_932;
input n_1102;
input n_1071;
input n_1107;
input n_705;
input n_586;
input n_760;
input n_191;
input n_207;
input n_842;
input n_268;
input n_761;
input n_326;
input n_777;
input n_155;
input n_493;
input n_222;
input n_41;
input n_351;
input n_0;
input n_1060;
input n_476;
input n_174;
input n_1033;
input n_892;
input n_531;
input n_235;
input n_479;
input n_474;
input n_557;
input n_600;
input n_975;
input n_649;
input n_58;
input n_974;
input n_1006;
input n_263;
input n_834;
input n_1074;
input n_963;
input n_874;
input n_1116;
input n_486;
input n_463;
input n_697;
input n_907;
input n_998;
input n_752;
input n_487;
input n_214;
input n_345;
input n_918;
input n_1022;
input n_668;
input n_193;
input n_739;
input n_391;
input n_337;
input n_1077;
input n_797;
input n_931;
input n_18;
input n_211;
input n_306;
input n_240;
input n_623;
input n_949;
input n_205;
input n_373;
input n_1020;
input n_930;
input n_114;
input n_267;
input n_427;
input n_741;
input n_863;
input n_1013;
input n_873;
input n_297;
input n_764;
input n_409;
input n_70;
input n_289;
input n_195;
input n_914;
input n_384;
input n_98;
input n_1047;
input n_259;
input n_269;
input n_349;
input n_159;
input n_805;
input n_929;
input n_652;
input n_43;
input n_14;
input n_165;
input n_372;
input n_13;
input n_430;
input n_1011;
input n_1094;
input n_994;
input n_1052;
input n_9;
input n_217;
input n_484;
input n_489;
input n_627;
input n_648;
input n_1003;
input n_495;
input n_137;
input n_346;
input n_286;
input n_611;
input n_612;
input n_706;
input n_1019;
input n_681;
input n_378;
input n_186;
input n_271;
input n_942;
input n_667;
input n_199;
input n_1026;
input n_824;
input n_334;
input n_906;
input n_1040;
input n_250;
input n_670;
input n_786;
input n_1049;
input n_446;
input n_494;
input n_642;
input n_591;
input n_1117;
input n_692;
input n_635;
input n_889;
input n_506;
input n_568;
input n_1114;
input n_1072;
input n_406;
input n_105;
input n_1002;
input n_404;
input n_1108;
input n_920;
input n_362;
input n_23;
input n_389;
input n_295;
input n_581;
input n_393;
input n_880;
input n_1051;
input n_832;
input n_720;
input n_328;

output n_7605;



endmodule