module fake_jpeg_2068_n_215 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_215);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_9),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_15),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_77),
.Y(n_92)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_70),
.Y(n_89)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_84),
.Y(n_93)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_75),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_60),
.B1(n_83),
.B2(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_69),
.B1(n_58),
.B2(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_69),
.B1(n_59),
.B2(n_73),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_98),
.B1(n_84),
.B2(n_86),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_69),
.B1(n_59),
.B2(n_71),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_102),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_54),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_118),
.B1(n_63),
.B2(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_108),
.Y(n_126)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_64),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_113),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_117),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_55),
.B1(n_58),
.B2(n_76),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_86),
.B1(n_61),
.B2(n_63),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_62),
.B1(n_74),
.B2(n_61),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_123),
.B1(n_128),
.B2(n_139),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_100),
.B1(n_106),
.B2(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_68),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_130),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_67),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_1),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_86),
.B(n_78),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_136),
.B(n_3),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_78),
.B1(n_66),
.B2(n_72),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_1),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_20),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_66),
.B1(n_72),
.B2(n_4),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_152),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_66),
.C(n_25),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_23),
.C(n_49),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_50),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_2),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_147),
.B(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_134),
.B(n_131),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_26),
.B1(n_48),
.B2(n_47),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_162),
.B1(n_42),
.B2(n_37),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_3),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_158),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_163),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_4),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_160),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_124),
.A2(n_19),
.B1(n_46),
.B2(n_43),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_124),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_166),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_171),
.B1(n_153),
.B2(n_162),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_36),
.B(n_35),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_175),
.B(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_34),
.B(n_30),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_190),
.B1(n_167),
.B2(n_185),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_187),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_145),
.B(n_161),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_186),
.A2(n_188),
.B1(n_192),
.B2(n_175),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_161),
.B1(n_142),
.B2(n_163),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_28),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_181),
.C(n_180),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_182),
.A2(n_164),
.B1(n_180),
.B2(n_169),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_170),
.B(n_27),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_197),
.B1(n_199),
.B2(n_178),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_202),
.B(n_204),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_181),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_205),
.C(n_198),
.Y(n_206)
);

XOR2x2_ASAP7_75t_SL g205 ( 
.A(n_193),
.B(n_11),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_207),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_196),
.C(n_12),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_209),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_208),
.C(n_205),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_16),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_11),
.B(n_12),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_13),
.Y(n_215)
);


endmodule