module real_aes_1273_n_335 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_335);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_335;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_635;
wire n_357;
wire n_503;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_865;
wire n_551;
wire n_884;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_550;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_875;
wire n_467;
wire n_951;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_702;
wire n_954;
wire n_912;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_749;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_831;
wire n_487;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_507;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_0), .A2(n_287), .B1(n_490), .B2(n_491), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_1), .A2(n_187), .B1(n_496), .B2(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_2), .A2(n_238), .B1(n_516), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_3), .A2(n_137), .B1(n_455), .B2(n_670), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_4), .A2(n_103), .B1(n_597), .B2(n_598), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_5), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_6), .A2(n_164), .B1(n_632), .B2(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_7), .B(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_8), .A2(n_218), .B1(n_490), .B2(n_491), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_9), .A2(n_158), .B1(n_513), .B2(n_720), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_10), .A2(n_244), .B1(n_371), .B2(n_586), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_11), .A2(n_320), .B1(n_783), .B2(n_784), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_12), .A2(n_172), .B1(n_498), .B2(n_499), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_13), .A2(n_69), .B1(n_380), .B2(n_720), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g753 ( .A1(n_14), .A2(n_72), .B1(n_485), .B2(n_486), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_15), .A2(n_283), .B1(n_462), .B2(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_16), .A2(n_161), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_17), .A2(n_188), .B1(n_483), .B2(n_544), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_18), .A2(n_151), .B1(n_592), .B2(n_659), .Y(n_658) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_19), .A2(n_149), .B1(n_496), .B2(n_551), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_20), .A2(n_306), .B1(n_511), .B2(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_21), .A2(n_119), .B1(n_518), .B2(n_651), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_22), .A2(n_54), .B1(n_419), .B2(n_516), .Y(n_824) );
AO222x2_ASAP7_75t_L g538 ( .A1(n_23), .A2(n_115), .B1(n_203), .B2(n_445), .C1(n_450), .C2(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_24), .A2(n_292), .B1(n_544), .B2(n_545), .Y(n_543) );
INVx1_ASAP7_75t_SL g365 ( .A(n_25), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g915 ( .A(n_25), .B(n_38), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_26), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g948 ( .A1(n_27), .A2(n_145), .B1(n_399), .B2(n_949), .Y(n_948) );
AOI22xp33_ASAP7_75t_SL g453 ( .A1(n_28), .A2(n_109), .B1(n_454), .B2(n_455), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_29), .B(n_673), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_30), .A2(n_254), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22x1_ASAP7_75t_L g760 ( .A1(n_31), .A2(n_166), .B1(n_465), .B2(n_498), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_32), .A2(n_97), .B1(n_544), .B2(n_545), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_33), .A2(n_186), .B1(n_384), .B2(n_391), .Y(n_383) );
OA22x2_ASAP7_75t_L g857 ( .A1(n_34), .A2(n_858), .B1(n_859), .B2(n_888), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_34), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_35), .A2(n_240), .B1(n_524), .B2(n_527), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_36), .A2(n_157), .B1(n_485), .B2(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_37), .A2(n_286), .B1(n_350), .B2(n_680), .Y(n_775) );
AO22x2_ASAP7_75t_L g368 ( .A1(n_38), .A2(n_311), .B1(n_356), .B2(n_369), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_39), .A2(n_144), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_40), .A2(n_181), .B1(n_371), .B2(n_509), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_41), .A2(n_313), .B1(n_511), .B2(n_513), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_42), .A2(n_49), .B1(n_516), .B2(n_610), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_43), .A2(n_285), .B1(n_371), .B2(n_509), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_44), .A2(n_154), .B1(n_430), .B2(n_622), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_45), .A2(n_245), .B1(n_350), .B2(n_468), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_46), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g366 ( .A(n_47), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_48), .A2(n_270), .B1(n_495), .B2(n_499), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_50), .A2(n_268), .B1(n_498), .B2(n_550), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_51), .A2(n_275), .B1(n_350), .B2(n_805), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_52), .A2(n_309), .B1(n_396), .B2(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_53), .A2(n_263), .B1(n_635), .B2(n_636), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_55), .A2(n_211), .B1(n_605), .B2(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_56), .A2(n_305), .B1(n_683), .B2(n_779), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_57), .A2(n_182), .B1(n_513), .B2(n_683), .Y(n_682) );
AO22x2_ASAP7_75t_L g359 ( .A1(n_58), .A2(n_163), .B1(n_356), .B2(n_360), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_59), .A2(n_271), .B1(n_371), .B2(n_592), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_60), .A2(n_114), .B1(n_499), .B2(n_847), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_61), .A2(n_202), .B1(n_391), .B2(n_462), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_62), .A2(n_90), .B1(n_448), .B2(n_451), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_63), .A2(n_134), .B1(n_485), .B2(n_486), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_64), .A2(n_280), .B1(n_375), .B2(n_465), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_65), .A2(n_138), .B1(n_499), .B2(n_550), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_66), .A2(n_170), .B1(n_350), .B2(n_680), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_67), .A2(n_127), .B1(n_465), .B2(n_470), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_68), .A2(n_93), .B1(n_490), .B2(n_491), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_70), .A2(n_169), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_71), .A2(n_250), .B1(n_550), .B2(n_551), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_73), .A2(n_214), .B1(n_450), .B2(n_451), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g881 ( .A1(n_74), .A2(n_312), .B1(n_882), .B2(n_883), .C(n_884), .Y(n_881) );
AOI222xp33_ASAP7_75t_L g528 ( .A1(n_75), .A2(n_120), .B1(n_198), .B2(n_429), .C1(n_529), .C2(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_76), .B(n_529), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_77), .A2(n_201), .B1(n_509), .B2(n_636), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_78), .A2(n_326), .B1(n_430), .B2(n_605), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g901 ( .A1(n_79), .A2(n_265), .B1(n_783), .B2(n_855), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_80), .A2(n_242), .B1(n_527), .B2(n_947), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_81), .A2(n_110), .B1(n_685), .B2(n_686), .Y(n_684) );
AO222x2_ASAP7_75t_L g568 ( .A1(n_82), .A2(n_180), .B1(n_317), .B2(n_445), .C1(n_483), .C2(n_486), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_83), .A2(n_104), .B1(n_588), .B2(n_589), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_84), .A2(n_199), .B1(n_482), .B2(n_483), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_85), .A2(n_200), .B1(n_622), .B2(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g862 ( .A(n_86), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_87), .A2(n_220), .B1(n_450), .B2(n_451), .Y(n_571) );
AOI222xp33_ASAP7_75t_L g902 ( .A1(n_88), .A2(n_147), .B1(n_299), .B2(n_430), .C1(n_530), .C2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_89), .A2(n_129), .B1(n_486), .B2(n_542), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_91), .A2(n_291), .B1(n_396), .B2(n_468), .Y(n_467) );
AO22x2_ASAP7_75t_L g355 ( .A1(n_92), .A2(n_248), .B1(n_356), .B2(n_357), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_94), .A2(n_262), .B1(n_612), .B2(n_651), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_95), .Y(n_871) );
OAI22x1_ASAP7_75t_L g821 ( .A1(n_96), .A2(n_822), .B1(n_837), .B2(n_838), .Y(n_821) );
CKINVDCx16_ASAP7_75t_R g838 ( .A(n_96), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_98), .A2(n_125), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_99), .A2(n_330), .B1(n_396), .B2(n_399), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_100), .A2(n_230), .B1(n_597), .B2(n_598), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_101), .A2(n_193), .B1(n_468), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_102), .A2(n_207), .B1(n_455), .B2(n_670), .Y(n_781) );
INVx1_ASAP7_75t_L g904 ( .A(n_105), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_106), .A2(n_304), .B1(n_491), .B2(n_733), .Y(n_732) );
OA22x2_ASAP7_75t_L g692 ( .A1(n_107), .A2(n_693), .B1(n_694), .B2(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_107), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_108), .A2(n_175), .B1(n_496), .B2(n_638), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_111), .A2(n_143), .B1(n_522), .B2(n_718), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_112), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_113), .A2(n_234), .B1(n_430), .B2(n_605), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_116), .A2(n_141), .B1(n_518), .B2(n_613), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_117), .A2(n_126), .B1(n_550), .B2(n_551), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_118), .A2(n_289), .B1(n_455), .B2(n_670), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_121), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_122), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_123), .A2(n_206), .B1(n_605), .B2(n_699), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_124), .B(n_606), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_128), .A2(n_189), .B1(n_468), .B2(n_831), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_130), .A2(n_331), .B1(n_680), .B2(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_131), .B(n_529), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_132), .A2(n_251), .B1(n_393), .B2(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_133), .A2(n_322), .B1(n_457), .B2(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_135), .B(n_603), .Y(n_649) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_136), .A2(n_279), .B1(n_462), .B2(n_463), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_139), .A2(n_253), .B1(n_371), .B2(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g806 ( .A1(n_140), .A2(n_264), .B1(n_391), .B2(n_462), .Y(n_806) );
INVx1_ASAP7_75t_L g790 ( .A(n_142), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_146), .A2(n_231), .B1(n_412), .B2(n_519), .Y(n_868) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_148), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_150), .A2(n_300), .B1(n_465), .B2(n_635), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_152), .A2(n_332), .B1(n_429), .B2(n_433), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_153), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_155), .A2(n_178), .B1(n_455), .B2(n_516), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_156), .A2(n_223), .B1(n_516), .B2(n_610), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_159), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_160), .A2(n_272), .B1(n_592), .B2(n_594), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_162), .A2(n_216), .B1(n_411), .B2(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g914 ( .A(n_163), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_165), .A2(n_197), .B1(n_498), .B2(n_499), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_167), .A2(n_224), .B1(n_490), .B2(n_491), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_168), .Y(n_879) );
XNOR2xp5_ASAP7_75t_L g744 ( .A(n_171), .B(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_173), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_174), .A2(n_314), .B1(n_419), .B2(n_516), .Y(n_625) );
INVx1_ASAP7_75t_L g601 ( .A(n_176), .Y(n_601) );
AOI22xp33_ASAP7_75t_SL g570 ( .A1(n_177), .A2(n_278), .B1(n_542), .B2(n_544), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_179), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_183), .A2(n_241), .B1(n_349), .B2(n_370), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_184), .A2(n_274), .B1(n_375), .B2(n_378), .Y(n_374) );
OA22x2_ASAP7_75t_L g770 ( .A1(n_185), .A2(n_771), .B1(n_772), .B2(n_787), .Y(n_770) );
INVxp67_ASAP7_75t_L g787 ( .A(n_185), .Y(n_787) );
INVx2_ASAP7_75t_L g927 ( .A(n_190), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_191), .A2(n_325), .B1(n_495), .B2(n_496), .Y(n_553) );
OA22x2_ASAP7_75t_L g663 ( .A1(n_192), .A2(n_664), .B1(n_687), .B2(n_688), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_192), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_194), .A2(n_235), .B1(n_597), .B2(n_882), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_195), .A2(n_208), .B1(n_471), .B2(n_683), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_196), .A2(n_217), .B1(n_454), .B2(n_455), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_204), .A2(n_243), .B1(n_527), .B2(n_632), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_205), .Y(n_886) );
CKINVDCx16_ASAP7_75t_R g738 ( .A(n_209), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_210), .A2(n_581), .B1(n_582), .B2(n_614), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_210), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_212), .A2(n_565), .B1(n_566), .B2(n_579), .Y(n_564) );
INVx1_ASAP7_75t_L g579 ( .A(n_212), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_213), .A2(n_298), .B1(n_457), .B2(n_458), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_215), .A2(n_935), .B1(n_956), .B2(n_957), .Y(n_955) );
CKINVDCx20_ASAP7_75t_R g957 ( .A(n_215), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_219), .A2(n_294), .B1(n_450), .B2(n_539), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_221), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_222), .A2(n_261), .B1(n_419), .B2(n_516), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_225), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_226), .A2(n_232), .B1(n_430), .B2(n_605), .Y(n_940) );
AOI22xp33_ASAP7_75t_SL g541 ( .A1(n_227), .A2(n_246), .B1(n_486), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_228), .A2(n_334), .B1(n_496), .B2(n_638), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_229), .A2(n_259), .B1(n_430), .B2(n_622), .Y(n_621) );
AOI222xp33_ASAP7_75t_L g929 ( .A1(n_233), .A2(n_930), .B1(n_953), .B2(n_955), .C1(n_958), .C2(n_959), .Y(n_929) );
XNOR2x1_ASAP7_75t_L g934 ( .A(n_233), .B(n_935), .Y(n_934) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_236), .A2(n_310), .B1(n_635), .B2(n_636), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_237), .A2(n_307), .B1(n_463), .B2(n_632), .Y(n_850) );
OA22x2_ASAP7_75t_L g343 ( .A1(n_239), .A2(n_344), .B1(n_345), .B2(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_239), .Y(n_344) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_247), .A2(n_288), .B1(n_399), .B2(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g912 ( .A(n_248), .B(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g928 ( .A(n_249), .Y(n_928) );
AOI222xp33_ASAP7_75t_L g835 ( .A1(n_252), .A2(n_260), .B1(n_295), .B2(n_445), .C1(n_539), .C2(n_836), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_255), .A2(n_297), .B1(n_495), .B2(n_496), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_256), .B(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_257), .A2(n_333), .B1(n_462), .B2(n_463), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_258), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_266), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_267), .A2(n_281), .B1(n_463), .B2(n_777), .Y(n_776) );
INVx3_ASAP7_75t_L g356 ( .A(n_269), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_273), .A2(n_282), .B1(n_495), .B2(n_496), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_276), .A2(n_321), .B1(n_412), .B2(n_784), .Y(n_797) );
OAI22x1_ASAP7_75t_L g646 ( .A1(n_277), .A2(n_647), .B1(n_660), .B2(n_661), .Y(n_646) );
INVx1_ASAP7_75t_L g661 ( .A(n_277), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_284), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_290), .A2(n_316), .B1(n_419), .B2(n_424), .Y(n_418) );
XNOR2x1_ASAP7_75t_L g842 ( .A(n_293), .B(n_843), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_296), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_301), .Y(n_709) );
INVx1_ASAP7_75t_L g440 ( .A(n_302), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_303), .A2(n_329), .B1(n_414), .B2(n_518), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_308), .A2(n_319), .B1(n_455), .B2(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g909 ( .A(n_315), .Y(n_909) );
NAND2xp5_ASAP7_75t_SL g926 ( .A(n_315), .B(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g910 ( .A(n_318), .Y(n_910) );
AND2x2_ASAP7_75t_R g958 ( .A(n_318), .B(n_909), .Y(n_958) );
OA22x2_ASAP7_75t_L g504 ( .A1(n_323), .A2(n_505), .B1(n_506), .B2(n_532), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_323), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_324), .B(n_926), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_327), .B(n_445), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_328), .B(n_529), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_916), .B(n_919), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_814), .B(n_906), .Y(n_336) );
INVx1_ASAP7_75t_L g917 ( .A(n_337), .Y(n_917) );
XNOR2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_641), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_558), .B2(n_559), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_501), .B1(n_556), .B2(n_557), .Y(n_340) );
INVx3_ASAP7_75t_L g557 ( .A(n_341), .Y(n_557) );
OA22x2_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_436), .B2(n_437), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NOR3x1_ASAP7_75t_SL g346 ( .A(n_347), .B(n_382), .C(n_402), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_374), .Y(n_347) );
BUFx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx3_ASAP7_75t_SL g470 ( .A(n_351), .Y(n_470) );
INVx2_ASAP7_75t_SL g522 ( .A(n_351), .Y(n_522) );
INVx4_ASAP7_75t_L g593 ( .A(n_351), .Y(n_593) );
INVx2_ASAP7_75t_L g635 ( .A(n_351), .Y(n_635) );
INVx8_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_361), .Y(n_352) );
AND2x4_ASAP7_75t_L g376 ( .A(n_353), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g398 ( .A(n_353), .B(n_390), .Y(n_398) );
AND2x2_ASAP7_75t_L g408 ( .A(n_353), .B(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g445 ( .A(n_353), .B(n_409), .Y(n_445) );
AND2x2_ASAP7_75t_L g495 ( .A(n_353), .B(n_377), .Y(n_495) );
AND2x6_ASAP7_75t_L g498 ( .A(n_353), .B(n_390), .Y(n_498) );
AND2x2_ASAP7_75t_L g550 ( .A(n_353), .B(n_361), .Y(n_550) );
AND2x2_ASAP7_75t_L g638 ( .A(n_353), .B(n_377), .Y(n_638) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_358), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g373 ( .A(n_355), .B(n_358), .Y(n_373) );
AND2x2_ASAP7_75t_L g381 ( .A(n_355), .B(n_359), .Y(n_381) );
INVx1_ASAP7_75t_L g389 ( .A(n_355), .Y(n_389) );
INVx2_ASAP7_75t_L g357 ( .A(n_356), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_356), .Y(n_360) );
OAI22x1_ASAP7_75t_L g363 ( .A1(n_356), .A2(n_364), .B1(n_365), .B2(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_356), .Y(n_364) );
INVx1_ASAP7_75t_L g369 ( .A(n_356), .Y(n_369) );
INVxp67_ASAP7_75t_L g417 ( .A(n_358), .Y(n_417) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g388 ( .A(n_359), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g372 ( .A(n_361), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g380 ( .A(n_361), .B(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g401 ( .A(n_361), .B(n_388), .Y(n_401) );
AND2x4_ASAP7_75t_L g496 ( .A(n_361), .B(n_381), .Y(n_496) );
AND2x6_ASAP7_75t_L g499 ( .A(n_361), .B(n_388), .Y(n_499) );
AND2x2_ASAP7_75t_L g551 ( .A(n_361), .B(n_373), .Y(n_551) );
AND2x4_ASAP7_75t_L g361 ( .A(n_362), .B(n_367), .Y(n_361) );
AND2x2_ASAP7_75t_L g390 ( .A(n_362), .B(n_368), .Y(n_390) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g377 ( .A(n_363), .B(n_367), .Y(n_377) );
AND2x2_ASAP7_75t_L g409 ( .A(n_363), .B(n_368), .Y(n_409) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_363), .Y(n_432) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
BUFx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_372), .Y(n_465) );
INVx2_ASAP7_75t_L g595 ( .A(n_372), .Y(n_595) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_372), .Y(n_636) );
AND2x4_ASAP7_75t_L g413 ( .A(n_373), .B(n_390), .Y(n_413) );
AND2x2_ASAP7_75t_L g435 ( .A(n_373), .B(n_377), .Y(n_435) );
AND2x4_ASAP7_75t_L g450 ( .A(n_373), .B(n_377), .Y(n_450) );
AND2x2_ASAP7_75t_L g485 ( .A(n_373), .B(n_390), .Y(n_485) );
AND2x2_ASAP7_75t_L g542 ( .A(n_373), .B(n_390), .Y(n_542) );
BUFx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx6_ASAP7_75t_L g512 ( .A(n_376), .Y(n_512) );
BUFx3_ASAP7_75t_L g720 ( .A(n_376), .Y(n_720) );
AND2x2_ASAP7_75t_L g427 ( .A(n_377), .B(n_388), .Y(n_427) );
AND2x4_ASAP7_75t_L g544 ( .A(n_377), .B(n_388), .Y(n_544) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_SL g779 ( .A(n_379), .Y(n_779) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g471 ( .A(n_380), .Y(n_471) );
BUFx3_ASAP7_75t_L g513 ( .A(n_380), .Y(n_513) );
BUFx2_ASAP7_75t_SL g598 ( .A(n_380), .Y(n_598) );
BUFx2_ASAP7_75t_SL g882 ( .A(n_380), .Y(n_882) );
AND2x4_ASAP7_75t_L g393 ( .A(n_381), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g431 ( .A(n_381), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_381), .B(n_432), .Y(n_451) );
AND2x4_ASAP7_75t_L g491 ( .A(n_381), .B(n_394), .Y(n_491) );
AND2x2_ASAP7_75t_SL g539 ( .A(n_381), .B(n_432), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_395), .Y(n_382) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g526 ( .A(n_386), .Y(n_526) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_387), .Y(n_462) );
BUFx3_ASAP7_75t_L g632 ( .A(n_387), .Y(n_632) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
AND2x2_ASAP7_75t_SL g490 ( .A(n_388), .B(n_390), .Y(n_490) );
AND2x2_ASAP7_75t_L g733 ( .A(n_388), .B(n_390), .Y(n_733) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_389), .Y(n_423) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g527 ( .A(n_392), .Y(n_527) );
INVx2_ASAP7_75t_L g589 ( .A(n_392), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g870 ( .A1(n_392), .A2(n_871), .B1(n_872), .B2(n_875), .Y(n_870) );
INVx5_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g463 ( .A(n_393), .Y(n_463) );
BUFx3_ASAP7_75t_L g715 ( .A(n_393), .Y(n_715) );
BUFx2_ASAP7_75t_L g829 ( .A(n_393), .Y(n_829) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g509 ( .A(n_397), .Y(n_509) );
INVx2_ASAP7_75t_SL g586 ( .A(n_397), .Y(n_586) );
INVx2_ASAP7_75t_L g685 ( .A(n_397), .Y(n_685) );
INVx2_ASAP7_75t_SL g949 ( .A(n_397), .Y(n_949) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g713 ( .A(n_398), .Y(n_713) );
BUFx2_ASAP7_75t_L g831 ( .A(n_398), .Y(n_831) );
INVx2_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g468 ( .A(n_400), .Y(n_468) );
INVx2_ASAP7_75t_SL g630 ( .A(n_400), .Y(n_630) );
INVx2_ASAP7_75t_L g659 ( .A(n_400), .Y(n_659) );
INVx2_ASAP7_75t_L g680 ( .A(n_400), .Y(n_680) );
INVx1_ASAP7_75t_SL g805 ( .A(n_400), .Y(n_805) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_400), .Y(n_887) );
INVx8_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND4xp25_ASAP7_75t_SL g402 ( .A(n_403), .B(n_410), .C(n_418), .D(n_428), .Y(n_402) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_406), .Y(n_603) );
INVx3_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx4_ASAP7_75t_SL g478 ( .A(n_407), .Y(n_478) );
INVx3_ASAP7_75t_L g529 ( .A(n_407), .Y(n_529) );
INVx3_ASAP7_75t_L g673 ( .A(n_407), .Y(n_673) );
INVx4_ASAP7_75t_SL g903 ( .A(n_407), .Y(n_903) );
INVx6_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g416 ( .A(n_409), .B(n_417), .Y(n_416) );
AND2x4_ASAP7_75t_L g421 ( .A(n_409), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g483 ( .A(n_409), .B(n_422), .Y(n_483) );
AND2x2_ASAP7_75t_L g486 ( .A(n_409), .B(n_417), .Y(n_486) );
AND2x2_ASAP7_75t_L g545 ( .A(n_409), .B(n_422), .Y(n_545) );
AND2x2_ASAP7_75t_L g826 ( .A(n_409), .B(n_417), .Y(n_826) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx4f_ASAP7_75t_SL g612 ( .A(n_412), .Y(n_612) );
INVx1_ASAP7_75t_L g708 ( .A(n_412), .Y(n_708) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx2_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
BUFx3_ASAP7_75t_L g518 ( .A(n_413), .Y(n_518) );
BUFx2_ASAP7_75t_L g783 ( .A(n_413), .Y(n_783) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g458 ( .A(n_415), .Y(n_458) );
INVx2_ASAP7_75t_L g519 ( .A(n_415), .Y(n_519) );
INVx2_ASAP7_75t_SL g613 ( .A(n_415), .Y(n_613) );
INVx2_ASAP7_75t_SL g651 ( .A(n_415), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_415), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g784 ( .A(n_415), .Y(n_784) );
INVx2_ASAP7_75t_L g855 ( .A(n_415), .Y(n_855) );
INVx6_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_SL g455 ( .A(n_421), .Y(n_455) );
BUFx4f_ASAP7_75t_L g610 ( .A(n_421), .Y(n_610) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx4_ASAP7_75t_L g482 ( .A(n_426), .Y(n_482) );
INVx2_ASAP7_75t_L g670 ( .A(n_426), .Y(n_670) );
INVx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_427), .Y(n_454) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_427), .Y(n_516) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx12f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g607 ( .A(n_431), .Y(n_607) );
INVx1_ASAP7_75t_L g863 ( .A(n_433), .Y(n_863) );
BUFx6f_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g531 ( .A(n_435), .Y(n_531) );
BUFx5_ASAP7_75t_L g605 ( .A(n_435), .Y(n_605) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B1(n_472), .B2(n_473), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
XNOR2x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
NAND2x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_459), .Y(n_441) );
NOR2xp67_ASAP7_75t_L g442 ( .A(n_443), .B(n_452), .Y(n_442) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_446), .B(n_447), .Y(n_443) );
OAI222xp33_ASAP7_75t_L g747 ( .A1(n_444), .A2(n_449), .B1(n_748), .B2(n_749), .C1(n_750), .C2(n_751), .Y(n_747) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_450), .Y(n_836) );
INVxp67_ASAP7_75t_L g751 ( .A(n_451), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g703 ( .A(n_454), .Y(n_703) );
INVxp67_ASAP7_75t_L g705 ( .A(n_455), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_466), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_464), .Y(n_460) );
INVx2_ASAP7_75t_L g880 ( .A(n_465), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
XOR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_500), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_475), .B(n_487), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .Y(n_476) );
INVx1_ASAP7_75t_SL g799 ( .A(n_478), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_484), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_493), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_492), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_497), .Y(n_493) );
INVx1_ASAP7_75t_L g848 ( .A(n_498), .Y(n_848) );
INVx1_ASAP7_75t_L g556 ( .A(n_501), .Y(n_556) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OAI22xp5_ASAP7_75t_SL g502 ( .A1(n_503), .A2(n_504), .B1(n_533), .B2(n_555), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_SL g532 ( .A(n_506), .Y(n_532) );
NAND4xp75_ASAP7_75t_L g506 ( .A(n_507), .B(n_514), .C(n_520), .D(n_528), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g597 ( .A(n_512), .Y(n_597) );
INVx2_ASAP7_75t_L g683 ( .A(n_512), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_512), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_884) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .Y(n_514) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g588 ( .A(n_525), .Y(n_588) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g777 ( .A(n_526), .Y(n_777) );
INVx1_ASAP7_75t_L g874 ( .A(n_526), .Y(n_874) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g622 ( .A(n_531), .Y(n_622) );
INVx1_ASAP7_75t_L g555 ( .A(n_533), .Y(n_555) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
XNOR2x1_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_546), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_552), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_615), .B1(n_616), .B2(n_640), .Y(n_560) );
INVx3_ASAP7_75t_L g640 ( .A(n_561), .Y(n_640) );
XNOR2x1_ASAP7_75t_L g561 ( .A(n_562), .B(n_580), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OA22x2_ASAP7_75t_L g840 ( .A1(n_563), .A2(n_564), .B1(n_841), .B2(n_842), .Y(n_840) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_567), .B(n_572), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_SL g614 ( .A(n_582), .Y(n_614) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_599), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_590), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_596), .Y(n_590) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g878 ( .A(n_593), .Y(n_878) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g686 ( .A(n_595), .Y(n_686) );
INVx1_ASAP7_75t_L g718 ( .A(n_595), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_608), .Y(n_599) );
OAI21xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B(n_604), .Y(n_600) );
INVx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx3_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g668 ( .A(n_607), .Y(n_668) );
INVx2_ASAP7_75t_L g699 ( .A(n_607), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVxp67_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
XOR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_639), .Y(n_617) );
NAND2x1p5_ASAP7_75t_L g618 ( .A(n_619), .B(n_627), .Y(n_618) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_620), .B(n_624), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_628), .B(n_633), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_637), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_765), .B1(n_766), .B2(n_813), .Y(n_641) );
INVx1_ASAP7_75t_L g813 ( .A(n_642), .Y(n_813) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_690), .B(n_762), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g764 ( .A(n_644), .Y(n_764) );
AO22x2_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_662), .B2(n_663), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g660 ( .A(n_647), .Y(n_660) );
OR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_654), .Y(n_647) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .C(n_652), .D(n_653), .Y(n_648) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .C(n_657), .D(n_658), .Y(n_654) );
AO22x2_ASAP7_75t_SL g788 ( .A1(n_662), .A2(n_663), .B1(n_789), .B2(n_811), .Y(n_788) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_676), .Y(n_664) );
NOR3xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_671), .C(n_674), .Y(n_665) );
NOR4xp25_ASAP7_75t_L g688 ( .A(n_666), .B(n_677), .C(n_681), .D(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVxp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_672), .B(n_675), .Y(n_689) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_681), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_690), .B(n_763), .Y(n_762) );
XNOR2x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_741), .Y(n_690) );
AO22x2_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_721), .B1(n_739), .B2(n_740), .Y(n_691) );
INVx1_ASAP7_75t_L g739 ( .A(n_692), .Y(n_739) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_710), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_701), .C(n_706), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_716), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
BUFx3_ASAP7_75t_L g883 ( .A(n_713), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
INVx1_ASAP7_75t_L g740 ( .A(n_721), .Y(n_740) );
XOR2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_738), .Y(n_721) );
NAND2x1p5_ASAP7_75t_L g722 ( .A(n_723), .B(n_730), .Y(n_722) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
NOR2x1_ASAP7_75t_L g730 ( .A(n_731), .B(n_735), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2x1p5_ASAP7_75t_L g745 ( .A(n_746), .B(n_755), .Y(n_745) );
NOR2x1_ASAP7_75t_L g746 ( .A(n_747), .B(n_752), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
NOR2x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVxp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OA21x2_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_788), .B(n_812), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_768), .B(n_788), .Y(n_812) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
NOR2x1_ASAP7_75t_L g772 ( .A(n_773), .B(n_780), .Y(n_772) );
NAND4xp25_ASAP7_75t_SL g773 ( .A(n_774), .B(n_775), .C(n_776), .D(n_778), .Y(n_773) );
NAND4xp25_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .C(n_785), .D(n_786), .Y(n_780) );
INVx2_ASAP7_75t_L g811 ( .A(n_789), .Y(n_811) );
OAI21x1_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B(n_810), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_790), .B(n_793), .Y(n_810) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_802), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_798), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
OAI21xp33_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B(n_801), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_799), .A2(n_862), .B1(n_863), .B2(n_864), .C(n_865), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_807), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_806), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
INVx1_ASAP7_75t_L g918 ( .A(n_814), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B1(n_890), .B2(n_905), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
AO22x1_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_818), .B1(n_857), .B2(n_889), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
AO22x2_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_820), .B1(n_839), .B2(n_840), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NAND4xp25_ASAP7_75t_SL g822 ( .A(n_823), .B(n_827), .C(n_832), .D(n_835), .Y(n_822) );
AND4x1_ASAP7_75t_L g837 ( .A(n_823), .B(n_827), .C(n_832), .D(n_835), .Y(n_837) );
AND2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
AND2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_830), .Y(n_827) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_SL g841 ( .A(n_842), .Y(n_841) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_844), .B(n_851), .Y(n_843) );
NAND4xp25_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .C(n_849), .D(n_850), .Y(n_844) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NAND4xp25_ASAP7_75t_SL g851 ( .A(n_852), .B(n_853), .C(n_854), .D(n_856), .Y(n_851) );
INVx1_ASAP7_75t_L g889 ( .A(n_857), .Y(n_889) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
AND3x2_ASAP7_75t_L g859 ( .A(n_860), .B(n_869), .C(n_881), .Y(n_859) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_866), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_870), .B(n_876), .Y(n_869) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g947 ( .A(n_874), .Y(n_947) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_876) );
INVx1_ASAP7_75t_L g905 ( .A(n_890), .Y(n_905) );
INVx3_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
XOR2x2_ASAP7_75t_L g891 ( .A(n_892), .B(n_904), .Y(n_891) );
NAND4xp75_ASAP7_75t_L g892 ( .A(n_893), .B(n_896), .C(n_899), .D(n_902), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
AND2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
AND2x2_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
INVx1_ASAP7_75t_L g938 ( .A(n_903), .Y(n_938) );
INVx1_ASAP7_75t_SL g906 ( .A(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_908), .B(n_911), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_908), .B(n_912), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_910), .Y(n_908) );
INVx1_ASAP7_75t_L g924 ( .A(n_910), .Y(n_924) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
OAI21xp5_ASAP7_75t_L g919 ( .A1(n_920), .A2(n_928), .B(n_929), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
BUFx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AND2x2_ASAP7_75t_SL g922 ( .A(n_923), .B(n_925), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
OR2x2_ASAP7_75t_L g960 ( .A(n_924), .B(n_925), .Y(n_960) );
INVx1_ASAP7_75t_SL g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVxp67_ASAP7_75t_SL g956 ( .A(n_935), .Y(n_956) );
AND2x4_ASAP7_75t_L g935 ( .A(n_936), .B(n_944), .Y(n_935) );
NOR2xp67_ASAP7_75t_L g936 ( .A(n_937), .B(n_941), .Y(n_936) );
OAI21xp5_ASAP7_75t_SL g937 ( .A1(n_938), .A2(n_939), .B(n_940), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_942), .B(n_943), .Y(n_941) );
NOR2x1_ASAP7_75t_L g944 ( .A(n_945), .B(n_950), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_946), .B(n_948), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_951), .B(n_952), .Y(n_950) );
CKINVDCx6p67_ASAP7_75t_R g953 ( .A(n_954), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_960), .Y(n_959) );
endmodule