module fake_jpeg_19911_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_3),
.B(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_18),
.B(n_37),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_0),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_49),
.B(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_1),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_75),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_89),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_2),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_48),
.B1(n_54),
.B2(n_55),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_83),
.B1(n_47),
.B2(n_56),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_41),
.B1(n_50),
.B2(n_38),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_10),
.B(n_12),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_1),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_96),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_94),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_44),
.B(n_5),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_98),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_4),
.B(n_7),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_13),
.B1(n_14),
.B2(n_19),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_106),
.B(n_93),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_24),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_109),
.Y(n_112)
);

AOI221xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_101),
.B1(n_100),
.B2(n_91),
.C(n_32),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_111),
.B1(n_110),
.B2(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_102),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_108),
.B1(n_105),
.B2(n_31),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_25),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_116),
.A2(n_30),
.B(n_35),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g119 ( 
.A(n_118),
.Y(n_119)
);


endmodule