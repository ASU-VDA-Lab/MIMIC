module fake_netlist_1_4055_n_33 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_7;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g7 ( .A(n_3), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_0), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_0), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_5), .Y(n_12) );
AOI22xp33_ASAP7_75t_L g13 ( .A1(n_8), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_13) );
O2A1O1Ixp33_ASAP7_75t_L g14 ( .A1(n_8), .A2(n_1), .B(n_2), .C(n_3), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_11), .B(n_1), .Y(n_15) );
A2O1A1Ixp33_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_4), .B(n_6), .C(n_9), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_7), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_17), .B(n_7), .Y(n_19) );
NOR2x1p5_ASAP7_75t_L g20 ( .A(n_15), .B(n_12), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_15), .B(n_6), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_18), .B(n_15), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
INVx2_ASAP7_75t_SL g24 ( .A(n_20), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
BUFx3_ASAP7_75t_L g26 ( .A(n_22), .Y(n_26) );
OAI211xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_16), .B(n_14), .C(n_13), .Y(n_27) );
AOI322xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_18), .A3(n_19), .B1(n_22), .B2(n_23), .C1(n_24), .C2(n_25), .Y(n_28) );
OAI211xp5_ASAP7_75t_SL g29 ( .A1(n_28), .A2(n_24), .B(n_25), .C(n_19), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_27), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
XNOR2xp5_ASAP7_75t_L g32 ( .A(n_29), .B(n_26), .Y(n_32) );
AOI222xp33_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_25), .B1(n_26), .B2(n_31), .C1(n_29), .C2(n_30), .Y(n_33) );
endmodule