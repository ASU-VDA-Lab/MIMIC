module fake_jpeg_625_n_119 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_5),
.B(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_0),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_50),
.Y(n_55)
);

OR2x4_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_0),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_37),
.B1(n_35),
.B2(n_40),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_56),
.B1(n_43),
.B2(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_49),
.B1(n_47),
.B2(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_59),
.B1(n_41),
.B2(n_2),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_34),
.B1(n_42),
.B2(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_1),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_33),
.B1(n_39),
.B2(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_70),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_41),
.B1(n_15),
.B2(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_66),
.B(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_3),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_3),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_41),
.C(n_18),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_55),
.C(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_68),
.C(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_4),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_5),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_62),
.B1(n_81),
.B2(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_92),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_67),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_32),
.B(n_27),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_93),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_95),
.C(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_54),
.B(n_7),
.C(n_8),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_7),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_19),
.C(n_30),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_6),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_99),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_6),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_103),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_94),
.B(n_85),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_104),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_25),
.C(n_23),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_10),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_104),
.B1(n_96),
.B2(n_11),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_9),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_112),
.C(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_113),
.B(n_106),
.Y(n_115)
);

NOR5xp2_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_109),
.C(n_114),
.D(n_22),
.E(n_13),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_109),
.C(n_11),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_12),
.Y(n_119)
);


endmodule