module fake_jpeg_18894_n_170 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_10),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_18),
.B(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_81),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_0),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NAND2x1_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_1),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_83),
.Y(n_98)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_52),
.B1(n_63),
.B2(n_55),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_70),
.B1(n_66),
.B2(n_60),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_64),
.B1(n_54),
.B2(n_65),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_70),
.B1(n_56),
.B2(n_69),
.Y(n_109)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_68),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_98),
.A2(n_83),
.B(n_59),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_97),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_106),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_109),
.B(n_111),
.C(n_74),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_73),
.B(n_68),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_58),
.B(n_57),
.C(n_4),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_74),
.B(n_75),
.C(n_76),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_91),
.B1(n_92),
.B2(n_67),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_120),
.B1(n_100),
.B2(n_5),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_125),
.B(n_7),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_72),
.B1(n_62),
.B2(n_61),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_123),
.B(n_6),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_101),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_1),
.B(n_2),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_127),
.A2(n_128),
.B(n_133),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_111),
.B(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_135),
.B1(n_138),
.B2(n_9),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_4),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_26),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_6),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_7),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_9),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_122),
.B1(n_115),
.B2(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_32),
.A3(n_44),
.B1(n_11),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_145),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_37),
.C(n_43),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_47),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_10),
.B(n_20),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_154),
.B(n_155),
.CI(n_140),
.CON(n_156),
.SN(n_156)
);

INVxp33_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_159),
.C(n_153),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_156),
.C(n_148),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_152),
.B1(n_156),
.B2(n_147),
.Y(n_167)
);

OAI321xp33_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_155),
.A3(n_144),
.B1(n_36),
.B2(n_39),
.C(n_25),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_30),
.B(n_40),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_42),
.Y(n_170)
);


endmodule