module fake_jpeg_31792_n_181 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_181);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_14),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_75),
.Y(n_83)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

NAND2x1_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_81),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_57),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_86),
.CI(n_62),
.CON(n_111),
.SN(n_111)
);

OR2x4_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_93),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_69),
.B1(n_44),
.B2(n_47),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_62),
.B1(n_60),
.B2(n_65),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_50),
.B(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_101),
.Y(n_119)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

BUFx24_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_47),
.B1(n_63),
.B2(n_64),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_108),
.B1(n_0),
.B2(n_2),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx5_ASAP7_75t_SL g104 ( 
.A(n_82),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_117),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_70),
.B1(n_52),
.B2(n_51),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_116),
.B1(n_10),
.B2(n_11),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_60),
.C(n_46),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_10),
.Y(n_136)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_114),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_56),
.Y(n_114)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_0),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_59),
.B1(n_53),
.B2(n_49),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_48),
.B1(n_45),
.B2(n_55),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_17),
.B(n_20),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_132),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_131),
.B1(n_41),
.B2(n_18),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_103),
.B(n_111),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_7),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_8),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_134),
.B(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_8),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_141),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_139),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_15),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_124),
.C(n_120),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_124),
.C(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_155),
.B1(n_125),
.B2(n_124),
.Y(n_159)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_158),
.A2(n_21),
.B(n_23),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_161),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_146),
.B(n_143),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_167),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_158),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_168),
.B(n_164),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_163),
.C(n_172),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_171),
.B1(n_153),
.B2(n_157),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_148),
.C(n_162),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_162),
.C(n_165),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_160),
.C(n_147),
.Y(n_179)
);

OAI322xp33_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_156),
.A3(n_170),
.B1(n_28),
.B2(n_29),
.C1(n_31),
.C2(n_33),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_156),
.Y(n_181)
);


endmodule