module fake_ariane_2456_n_1789 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1789);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1789;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_105),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_45),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_72),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_77),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_76),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_73),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_108),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_3),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_149),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_32),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_36),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_32),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_43),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_39),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_51),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_33),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_94),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_154),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_41),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_66),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_93),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_147),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_38),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_33),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_61),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_37),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_20),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_39),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_34),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_20),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_129),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_84),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_113),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_136),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_143),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_13),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_28),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_15),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_134),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_101),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_25),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_107),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_42),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_79),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_58),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_144),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_56),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_92),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_110),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_151),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_155),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_96),
.Y(n_220)
);

BUFx8_ASAP7_75t_SL g221 ( 
.A(n_98),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_45),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_21),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_25),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_121),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_26),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_140),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_54),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_82),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_37),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_43),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_91),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_13),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_99),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_12),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_97),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_6),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_17),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_44),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_127),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_74),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_153),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_95),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_69),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_106),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_36),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_24),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_68),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_90),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_131),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_123),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_9),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_78),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_46),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_81),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_150),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_156),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_89),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_6),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_86),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_48),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_9),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_17),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_18),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_4),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_19),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_104),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_130),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_124),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_65),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_1),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_18),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_49),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_30),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_16),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_55),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_103),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_115),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_27),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_5),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_29),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_83),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_70),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_87),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_31),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_64),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_138),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_5),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_60),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_132),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_50),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_53),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_44),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_128),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_11),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_1),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_8),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_117),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_114),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_137),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_8),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_4),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_126),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_63),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_10),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_71),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_48),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_40),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_38),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_41),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_221),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_173),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_267),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_160),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_160),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_179),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_161),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_161),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_165),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_157),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_200),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_165),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_173),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_214),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_166),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_166),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_171),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_242),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_171),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_179),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_181),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_222),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_237),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_181),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_186),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_292),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_186),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_187),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_187),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_222),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_237),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_201),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_201),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_210),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_182),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_210),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_182),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_158),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_216),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_307),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_311),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_307),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_216),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_192),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_159),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_175),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_220),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_263),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_220),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_225),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_176),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_177),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_178),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_167),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_185),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_225),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_189),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_311),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_311),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_227),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_227),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_196),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_194),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_298),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_196),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_304),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_236),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_236),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_246),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_311),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_246),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_257),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_219),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_195),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_280),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_205),
.Y(n_390)
);

CKINVDCx8_ASAP7_75t_R g391 ( 
.A(n_313),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_250),
.Y(n_392)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_342),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_358),
.B(n_306),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_384),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_355),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_317),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_319),
.B(n_162),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_319),
.B(n_229),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_362),
.A2(n_312),
.B1(n_233),
.B2(n_254),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_320),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_314),
.B(n_228),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_321),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_324),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_324),
.B(n_257),
.Y(n_411)
);

NOR2x1_ASAP7_75t_L g412 ( 
.A(n_328),
.B(n_164),
.Y(n_412)
);

NOR2x1_ASAP7_75t_L g413 ( 
.A(n_328),
.B(n_164),
.Y(n_413)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_329),
.A2(n_278),
.B(n_258),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_330),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_332),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_334),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_378),
.A2(n_380),
.B1(n_339),
.B2(n_322),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g422 ( 
.A(n_334),
.B(n_162),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_337),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_338),
.B(n_258),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_340),
.B(n_190),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_323),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_340),
.A2(n_305),
.B(n_278),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_318),
.B(n_228),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_327),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_343),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_331),
.Y(n_436)
);

CKINVDCx6p67_ASAP7_75t_R g437 ( 
.A(n_368),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_346),
.B(n_190),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_347),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_333),
.B(n_228),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_347),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_348),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_365),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_350),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_353),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_357),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_342),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_357),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_361),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_335),
.B(n_215),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_361),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_363),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_363),
.B(n_311),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_387),
.B(n_215),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_452),
.B(n_342),
.Y(n_460)
);

NOR2x1p5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_446),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_398),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_352),
.Y(n_463)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_398),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_398),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_452),
.B(n_367),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_398),
.B(n_370),
.C(n_364),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_389),
.B(n_369),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_398),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_407),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_407),
.A2(n_325),
.B1(n_386),
.B2(n_385),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_393),
.B(n_371),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_400),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_400),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_393),
.B(n_325),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_428),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_455),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_400),
.Y(n_480)
);

AOI21x1_ASAP7_75t_L g481 ( 
.A1(n_414),
.A2(n_429),
.B(n_425),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_L g483 ( 
.A(n_400),
.B(n_377),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_393),
.B(n_364),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_393),
.B(n_370),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_405),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_403),
.B(n_374),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_405),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_405),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_403),
.B(n_359),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_SL g492 ( 
.A(n_438),
.B(n_388),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_396),
.B(n_374),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_375),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_455),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_408),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_430),
.B(n_336),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_430),
.B(n_315),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_444),
.B(n_375),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_408),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_416),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_434),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_427),
.B(n_344),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_444),
.B(n_381),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_416),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_416),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_444),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_416),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_416),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_416),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_432),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_432),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_432),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_432),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_432),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_432),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_417),
.B(n_381),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_435),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_435),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_435),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_435),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_435),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_435),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_450),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_442),
.B(n_354),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_427),
.A2(n_386),
.B1(n_385),
.B2(n_383),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_450),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_442),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_450),
.Y(n_535)
);

CKINVDCx6p67_ASAP7_75t_R g536 ( 
.A(n_437),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_450),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_417),
.B(n_382),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_417),
.B(n_382),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_427),
.B(n_383),
.Y(n_540)
);

NOR3xp33_ASAP7_75t_L g541 ( 
.A(n_438),
.B(n_193),
.C(n_356),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_450),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_459),
.A2(n_360),
.B1(n_366),
.B2(n_223),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_427),
.B(n_326),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_L g545 ( 
.A(n_450),
.B(n_163),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_436),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_457),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_457),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_439),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_457),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_459),
.B(n_349),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_457),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_457),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_439),
.B(n_417),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_457),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_397),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_439),
.A2(n_268),
.B1(n_203),
.B2(n_204),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_439),
.A2(n_268),
.B1(n_203),
.B2(n_204),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_391),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_418),
.B(n_351),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_397),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_390),
.B(n_376),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_418),
.B(n_379),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_418),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_437),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_418),
.B(n_170),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_390),
.B(n_392),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_433),
.A2(n_310),
.B1(n_202),
.B2(n_208),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_392),
.A2(n_266),
.B1(n_224),
.B2(n_303),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_433),
.B(n_180),
.Y(n_570)
);

INVx4_ASAP7_75t_SL g571 ( 
.A(n_402),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_404),
.A2(n_275),
.B1(n_235),
.B2(n_299),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_433),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_411),
.B(n_211),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_433),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_401),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_454),
.Y(n_577)
);

BUFx8_ASAP7_75t_SL g578 ( 
.A(n_391),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_454),
.B(n_239),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_454),
.B(n_240),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_454),
.B(n_305),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_401),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_391),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_401),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_399),
.B(n_289),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_399),
.B(n_272),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_411),
.B(n_211),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_409),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_458),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_406),
.B(n_241),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_406),
.B(n_256),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_409),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_409),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_410),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_410),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_412),
.A2(n_309),
.B1(n_281),
.B2(n_232),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_410),
.Y(n_597)
);

AO21x2_ASAP7_75t_L g598 ( 
.A1(n_414),
.A2(n_259),
.B(n_217),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_458),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_415),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_415),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_415),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_426),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_426),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_426),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_395),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_419),
.B(n_284),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_419),
.B(n_284),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_448),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_412),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_573),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_490),
.B(n_420),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_567),
.A2(n_441),
.B1(n_420),
.B2(n_453),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_573),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_562),
.B(n_423),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_599),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_544),
.B(n_395),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_601),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_470),
.B(n_423),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_577),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_544),
.B(n_424),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_463),
.B(n_424),
.Y(n_622)
);

NOR3xp33_ASAP7_75t_L g623 ( 
.A(n_569),
.B(n_425),
.C(n_404),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_549),
.B(n_431),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_564),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_554),
.B(n_458),
.Y(n_626)
);

NAND3xp33_ASAP7_75t_L g627 ( 
.A(n_468),
.B(n_440),
.C(n_431),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_470),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_479),
.B(n_440),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_601),
.Y(n_630)
);

NAND2x1_ASAP7_75t_L g631 ( 
.A(n_516),
.B(n_441),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_601),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_564),
.B(n_443),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_564),
.B(n_443),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_513),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_549),
.B(n_445),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_564),
.B(n_445),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_544),
.B(n_447),
.Y(n_638)
);

NOR3xp33_ASAP7_75t_L g639 ( 
.A(n_531),
.B(n_449),
.C(n_447),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_508),
.B(n_453),
.C(n_451),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_479),
.B(n_497),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_L g642 ( 
.A(n_504),
.B(n_449),
.C(n_451),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_484),
.A2(n_429),
.B(n_414),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_575),
.B(n_448),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_534),
.Y(n_645)
);

INVxp33_ASAP7_75t_L g646 ( 
.A(n_578),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_508),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_575),
.Y(n_648)
);

OAI221xp5_ASAP7_75t_L g649 ( 
.A1(n_471),
.A2(n_248),
.B1(n_283),
.B2(n_282),
.C(n_281),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_601),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_497),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_534),
.B(n_448),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_513),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_554),
.A2(n_413),
.B1(n_456),
.B2(n_422),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_487),
.B(n_456),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_540),
.B(n_456),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_546),
.B(n_413),
.C(n_277),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_599),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_575),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_540),
.B(n_458),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_513),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_461),
.B(n_232),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_R g663 ( 
.A(n_559),
.B(n_394),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_601),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_575),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_576),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_584),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_560),
.B(n_402),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_584),
.Y(n_669)
);

INVxp67_ASAP7_75t_SL g670 ( 
.A(n_589),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_563),
.B(n_402),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_477),
.B(n_261),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_588),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_588),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_585),
.B(n_402),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_509),
.B(n_402),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_576),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_603),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_546),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_544),
.B(n_248),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_492),
.B(n_293),
.C(n_264),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_509),
.B(n_402),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_485),
.B(n_429),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_559),
.B(n_274),
.Y(n_684)
);

O2A1O1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_523),
.A2(n_283),
.B(n_309),
.C(n_295),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_610),
.B(n_276),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_610),
.B(n_402),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_460),
.B(n_402),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_503),
.A2(n_422),
.B1(n_197),
.B2(n_252),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_543),
.B(n_287),
.C(n_297),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_532),
.B(n_422),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_576),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_574),
.B(n_422),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_551),
.B(n_290),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_473),
.B(n_516),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_SL g696 ( 
.A1(n_572),
.A2(n_295),
.B1(n_273),
.B2(n_265),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_574),
.B(n_422),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_SL g698 ( 
.A1(n_606),
.A2(n_421),
.B1(n_572),
.B2(n_583),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_603),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_583),
.B(n_215),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_466),
.B(n_474),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_589),
.B(n_249),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_582),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_483),
.A2(n_422),
.B1(n_183),
.B2(n_184),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_599),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_587),
.B(n_422),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_604),
.Y(n_707)
);

NOR2x1p5_ASAP7_75t_L g708 ( 
.A(n_536),
.B(n_587),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_478),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_473),
.B(n_198),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_493),
.A2(n_249),
.B1(n_273),
.B2(n_265),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_590),
.B(n_282),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_604),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_566),
.B(n_422),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_461),
.B(n_570),
.Y(n_715)
);

BUFx6f_ASAP7_75t_SL g716 ( 
.A(n_478),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_582),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_582),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_557),
.A2(n_253),
.B1(n_198),
.B2(n_259),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_600),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_599),
.A2(n_168),
.B1(n_169),
.B2(n_301),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_505),
.B(n_510),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_558),
.A2(n_605),
.B1(n_597),
.B2(n_594),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_496),
.B(n_394),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_592),
.A2(n_253),
.B1(n_217),
.B2(n_234),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_600),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_538),
.B(n_394),
.Y(n_727)
);

O2A1O1Ixp5_ASAP7_75t_L g728 ( 
.A1(n_579),
.A2(n_234),
.B(n_394),
.C(n_251),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_539),
.B(n_172),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_565),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_473),
.B(n_302),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_600),
.B(n_586),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_600),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_473),
.B(n_516),
.Y(n_734)
);

BUFx4f_ASAP7_75t_L g735 ( 
.A(n_536),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_473),
.B(n_302),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_607),
.B(n_174),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_556),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_565),
.B(n_0),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_580),
.A2(n_247),
.B1(n_191),
.B2(n_199),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_592),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_571),
.B(n_0),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_478),
.B(n_421),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_606),
.B(n_2),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_478),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_476),
.B(n_188),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_571),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_608),
.B(n_593),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_568),
.B(n_2),
.Y(n_749)
);

O2A1O1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_581),
.A2(n_591),
.B(n_602),
.C(n_609),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_593),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_541),
.B(n_206),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_556),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_596),
.B(n_3),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_561),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_609),
.B(n_207),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_594),
.B(n_209),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_595),
.B(n_7),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_602),
.B(n_212),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_595),
.B(n_7),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_516),
.B(n_213),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_597),
.B(n_218),
.Y(n_762)
);

OR2x2_ASAP7_75t_SL g763 ( 
.A(n_467),
.B(n_302),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_502),
.B(n_302),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_502),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_561),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_476),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_472),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_476),
.B(n_529),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_472),
.Y(n_770)
);

AND2x6_ASAP7_75t_L g771 ( 
.A(n_502),
.B(n_506),
.Y(n_771)
);

BUFx12f_ASAP7_75t_SL g772 ( 
.A(n_571),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_464),
.B(n_226),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_476),
.B(n_11),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_464),
.B(n_270),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_482),
.A2(n_271),
.B1(n_231),
.B2(n_300),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_L g777 ( 
.A(n_529),
.B(n_230),
.C(n_238),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_529),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_462),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_482),
.A2(n_279),
.B1(n_244),
.B2(n_296),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_464),
.B(n_308),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_647),
.B(n_529),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_612),
.A2(n_488),
.B1(n_489),
.B2(n_553),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_747),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_611),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_612),
.B(n_488),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_623),
.A2(n_754),
.B1(n_698),
.B2(n_649),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_617),
.B(n_506),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_747),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_666),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_679),
.B(n_506),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_614),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_705),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_677),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_735),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_622),
.B(n_489),
.Y(n_796)
);

AOI21x1_ASAP7_75t_L g797 ( 
.A1(n_683),
.A2(n_481),
.B(n_520),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_615),
.B(n_491),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_619),
.B(n_491),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_739),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_623),
.A2(n_522),
.B1(n_462),
.B2(n_555),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_735),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_692),
.Y(n_803)
);

NOR2xp67_ASAP7_75t_L g804 ( 
.A(n_730),
.B(n_514),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_739),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_616),
.B(n_464),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_745),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_651),
.B(n_494),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_620),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_SL g810 ( 
.A(n_640),
.B(n_634),
.C(n_633),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_719),
.A2(n_524),
.B1(n_465),
.B2(n_555),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_742),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_663),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_769),
.A2(n_519),
.B(n_553),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_667),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_616),
.B(n_464),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_R g817 ( 
.A(n_772),
.B(n_481),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_743),
.B(n_514),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_703),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_705),
.Y(n_820)
);

AND2x6_ASAP7_75t_L g821 ( 
.A(n_742),
.B(n_514),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_717),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_670),
.A2(n_641),
.B1(n_626),
.B2(n_686),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_718),
.Y(n_824)
);

NAND2x1p5_ASAP7_75t_L g825 ( 
.A(n_635),
.B(n_464),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_635),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_670),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_626),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_702),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_653),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_708),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_626),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_741),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_658),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_619),
.B(n_494),
.Y(n_835)
);

NAND3xp33_ASAP7_75t_SL g836 ( 
.A(n_749),
.B(n_269),
.C(n_255),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_651),
.B(n_645),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_751),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_621),
.B(n_571),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_641),
.A2(n_520),
.B1(n_495),
.B2(n_498),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_626),
.Y(n_841)
);

AND2x2_ASAP7_75t_SL g842 ( 
.A(n_719),
.B(n_515),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_669),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_673),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_730),
.B(n_515),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_663),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_674),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_678),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_645),
.B(n_495),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_SL g850 ( 
.A1(n_696),
.A2(n_260),
.B1(n_243),
.B2(n_262),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_628),
.B(n_498),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_699),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_638),
.B(n_515),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_658),
.B(n_511),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_652),
.B(n_499),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_765),
.B(n_511),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_656),
.A2(n_499),
.B(n_500),
.C(n_507),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_766),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_707),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_720),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_765),
.B(n_511),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_733),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_701),
.B(n_500),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_652),
.B(n_507),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_662),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_738),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_713),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_R g868 ( 
.A(n_716),
.B(n_512),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_626),
.B(n_512),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_702),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_765),
.B(n_511),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_690),
.A2(n_598),
.B1(n_245),
.B2(n_294),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_686),
.A2(n_526),
.B1(n_517),
.B2(n_519),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_672),
.B(n_517),
.Y(n_874)
);

AND2x2_ASAP7_75t_SL g875 ( 
.A(n_725),
.B(n_518),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_765),
.B(n_701),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_767),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_771),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_672),
.B(n_526),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_711),
.A2(n_680),
.B1(n_676),
.B2(n_682),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_767),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_778),
.B(n_613),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_753),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_755),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_778),
.B(n_675),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_SL g886 ( 
.A1(n_744),
.A2(n_291),
.B1(n_288),
.B2(n_286),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_625),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_771),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_648),
.Y(n_889)
);

OR2x6_ASAP7_75t_L g890 ( 
.A(n_709),
.B(n_518),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_642),
.B(n_465),
.Y(n_891)
);

BUFx8_ASAP7_75t_L g892 ( 
.A(n_646),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_659),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_627),
.B(n_527),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_SL g895 ( 
.A1(n_694),
.A2(n_598),
.B1(n_285),
.B2(n_550),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_771),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_665),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_726),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_660),
.B(n_527),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_655),
.B(n_528),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_653),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_693),
.B(n_697),
.Y(n_902)
);

BUFx4f_ASAP7_75t_L g903 ( 
.A(n_771),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_779),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_771),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_642),
.B(n_469),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_768),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_639),
.B(n_469),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_661),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_764),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_618),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_706),
.B(n_511),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_694),
.B(n_528),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_631),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_770),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_624),
.B(n_511),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_R g917 ( 
.A(n_715),
.B(n_537),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_630),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_636),
.B(n_530),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_722),
.B(n_537),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_644),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_632),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_650),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_644),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_664),
.B(n_661),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_714),
.B(n_525),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_712),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_633),
.Y(n_928)
);

INVx5_ASAP7_75t_L g929 ( 
.A(n_764),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_684),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_637),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_639),
.A2(n_525),
.B1(n_552),
.B2(n_550),
.Y(n_932)
);

INVx5_ASAP7_75t_L g933 ( 
.A(n_764),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_758),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_760),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_637),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_712),
.B(n_530),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_748),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_629),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_724),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_723),
.B(n_533),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_681),
.B(n_524),
.Y(n_942)
);

NOR3xp33_ASAP7_75t_SL g943 ( 
.A(n_657),
.B(n_12),
.C(n_14),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_727),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_700),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_763),
.Y(n_946)
);

BUFx4f_ASAP7_75t_L g947 ( 
.A(n_764),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_764),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_732),
.Y(n_949)
);

NAND2x1p5_ASAP7_75t_L g950 ( 
.A(n_695),
.B(n_522),
.Y(n_950)
);

OR2x6_ASAP7_75t_L g951 ( 
.A(n_752),
.B(n_521),
.Y(n_951)
);

NOR2x1p5_ASAP7_75t_L g952 ( 
.A(n_737),
.B(n_729),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_L g953 ( 
.A(n_711),
.B(n_545),
.C(n_480),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_723),
.B(n_533),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_654),
.B(n_535),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_689),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_695),
.Y(n_957)
);

INVx5_ASAP7_75t_L g958 ( 
.A(n_734),
.Y(n_958)
);

BUFx12f_ASAP7_75t_L g959 ( 
.A(n_777),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_721),
.B(n_535),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_691),
.B(n_521),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_687),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_668),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_750),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_774),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_774),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_688),
.B(n_501),
.Y(n_967)
);

BUFx8_ASAP7_75t_L g968 ( 
.A(n_777),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_671),
.Y(n_969)
);

XOR2x2_ASAP7_75t_L g970 ( 
.A(n_850),
.B(n_740),
.Y(n_970)
);

AOI21x1_ASAP7_75t_L g971 ( 
.A1(n_965),
.A2(n_683),
.B(n_710),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_868),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_868),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_898),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_786),
.A2(n_643),
.B(n_734),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_827),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_829),
.B(n_776),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_823),
.B(n_780),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_827),
.Y(n_979)
);

INVx6_ASAP7_75t_L g980 ( 
.A(n_795),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_870),
.B(n_756),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_813),
.B(n_757),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_927),
.B(n_759),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_837),
.B(n_725),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_784),
.Y(n_985)
);

OR2x6_ASAP7_75t_SL g986 ( 
.A(n_945),
.B(n_762),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_966),
.A2(n_746),
.B(n_761),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_837),
.B(n_685),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_784),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_865),
.B(n_552),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_863),
.A2(n_728),
.B(n_542),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_874),
.A2(n_775),
.B(n_773),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_785),
.Y(n_993)
);

NAND2x1p5_ASAP7_75t_L g994 ( 
.A(n_828),
.B(n_781),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_SL g995 ( 
.A(n_795),
.B(n_547),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_SL g996 ( 
.A1(n_796),
.A2(n_548),
.B(n_480),
.C(n_486),
.Y(n_996)
);

OAI21xp33_ASAP7_75t_SL g997 ( 
.A1(n_830),
.A2(n_781),
.B(n_710),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_800),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_846),
.B(n_704),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_787),
.A2(n_542),
.B1(n_475),
.B2(n_486),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_788),
.B(n_475),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_879),
.A2(n_547),
.B(n_548),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_797),
.A2(n_501),
.B(n_731),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_901),
.A2(n_736),
.B1(n_731),
.B2(n_308),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_802),
.Y(n_1005)
);

OR2x6_ASAP7_75t_SL g1006 ( 
.A(n_968),
.B(n_14),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_882),
.A2(n_736),
.B(n_598),
.C(n_19),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_828),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_787),
.B(n_15),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_885),
.A2(n_308),
.B(n_302),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_812),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_SL g1012 ( 
.A(n_896),
.B(n_308),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_832),
.B(n_841),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_882),
.A2(n_16),
.B(n_21),
.C(n_22),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_885),
.A2(n_308),
.B(n_23),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_796),
.A2(n_22),
.B(n_23),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_832),
.B(n_24),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_807),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_836),
.B(n_26),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_909),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_938),
.B(n_30),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_792),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_938),
.B(n_31),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_892),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_818),
.B(n_34),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_841),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_909),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_812),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_863),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_805),
.B(n_930),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_903),
.B(n_47),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_807),
.Y(n_1032)
);

BUFx12f_ASAP7_75t_L g1033 ( 
.A(n_892),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_809),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_968),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_903),
.B(n_49),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_940),
.B(n_50),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_898),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_939),
.B(n_52),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_849),
.B(n_944),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_849),
.B(n_57),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_866),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_946),
.B(n_59),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_839),
.B(n_913),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_799),
.A2(n_62),
.B(n_67),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_886),
.A2(n_959),
.B1(n_821),
.B2(n_913),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_907),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_831),
.B(n_152),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_SL g1049 ( 
.A(n_887),
.B(n_80),
.C(n_85),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_839),
.B(n_109),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_SL g1051 ( 
.A(n_889),
.B(n_111),
.C(n_118),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_798),
.A2(n_120),
.B(n_133),
.C(n_139),
.Y(n_1052)
);

AOI21x1_ASAP7_75t_L g1053 ( 
.A1(n_964),
.A2(n_141),
.B(n_146),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_810),
.A2(n_894),
.B(n_808),
.C(n_934),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_835),
.A2(n_920),
.B(n_864),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_959),
.A2(n_821),
.B1(n_853),
.B2(n_808),
.Y(n_1056)
);

NAND3xp33_ASAP7_75t_SL g1057 ( 
.A(n_943),
.B(n_810),
.C(n_872),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_878),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_880),
.A2(n_815),
.B1(n_847),
.B2(n_867),
.Y(n_1059)
);

INVxp67_ASAP7_75t_SL g1060 ( 
.A(n_878),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_853),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_915),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_876),
.B(n_877),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_894),
.A2(n_935),
.B(n_934),
.C(n_851),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_SL g1065 ( 
.A(n_896),
.B(n_905),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_905),
.B(n_888),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_SL g1067 ( 
.A(n_893),
.B(n_897),
.C(n_783),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_883),
.A2(n_884),
.B1(n_858),
.B2(n_880),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_876),
.B(n_877),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_883),
.Y(n_1070)
);

AO21x1_ASAP7_75t_L g1071 ( 
.A1(n_916),
.A2(n_925),
.B(n_912),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_804),
.B(n_935),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_845),
.B(n_943),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_851),
.A2(n_873),
.B(n_857),
.C(n_952),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_884),
.A2(n_858),
.B1(n_949),
.B2(n_833),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_834),
.B(n_791),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_881),
.B(n_949),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_899),
.A2(n_855),
.B(n_852),
.C(n_848),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_821),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_881),
.B(n_843),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_821),
.B(n_890),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_844),
.B(n_859),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_833),
.A2(n_838),
.B1(n_842),
.B2(n_904),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_902),
.A2(n_967),
.B(n_900),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_956),
.A2(n_906),
.B(n_936),
.C(n_928),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_888),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_838),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_790),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_890),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_902),
.A2(n_967),
.B(n_912),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_931),
.B(n_842),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_911),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_921),
.A2(n_924),
.B(n_916),
.C(n_919),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_890),
.B(n_782),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_790),
.Y(n_1095)
);

OAI22x1_ASAP7_75t_L g1096 ( 
.A1(n_942),
.A2(n_908),
.B1(n_891),
.B2(n_906),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_794),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_951),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_789),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_926),
.A2(n_814),
.B(n_919),
.Y(n_1100)
);

OAI22x1_ASAP7_75t_L g1101 ( 
.A1(n_942),
.A2(n_908),
.B1(n_891),
.B2(n_906),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_834),
.B(n_957),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_794),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_957),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_926),
.A2(n_816),
.B(n_854),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_951),
.B(n_860),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_957),
.B(n_911),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_950),
.A2(n_963),
.B(n_955),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_951),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_789),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_950),
.A2(n_963),
.B(n_954),
.Y(n_1111)
);

INVx3_ASAP7_75t_SL g1112 ( 
.A(n_957),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_840),
.A2(n_793),
.B1(n_820),
.B2(n_826),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_SL g1114 ( 
.A(n_948),
.B(n_947),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_937),
.B(n_862),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1100),
.A2(n_925),
.B(n_856),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1100),
.A2(n_871),
.B(n_861),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1040),
.B(n_875),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_979),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1011),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1055),
.A2(n_1041),
.B(n_975),
.Y(n_1121)
);

AOI31xp67_ASAP7_75t_L g1122 ( 
.A1(n_978),
.A2(n_871),
.A3(n_856),
.B(n_861),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1111),
.A2(n_962),
.B(n_941),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_983),
.A2(n_895),
.B(n_953),
.C(n_960),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1009),
.A2(n_869),
.B1(n_875),
.B2(n_793),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_998),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_977),
.B(n_918),
.Y(n_1127)
);

NAND2x1p5_ASAP7_75t_L g1128 ( 
.A(n_1081),
.B(n_820),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_SL g1129 ( 
.A(n_1114),
.B(n_948),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1108),
.A2(n_962),
.B(n_801),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1003),
.A2(n_801),
.B(n_854),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1054),
.B(n_1059),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_975),
.A2(n_932),
.B(n_961),
.Y(n_1133)
);

AO21x2_ASAP7_75t_L g1134 ( 
.A1(n_1055),
.A2(n_1090),
.B(n_1084),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_993),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1077),
.B(n_862),
.Y(n_1136)
);

OA21x2_ASAP7_75t_L g1137 ( 
.A1(n_1090),
.A2(n_922),
.B(n_923),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1028),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1084),
.A2(n_816),
.B(n_806),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1064),
.A2(n_961),
.B(n_860),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1022),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_976),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1010),
.A2(n_806),
.B(n_803),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_1033),
.Y(n_1144)
);

AOI221xp5_ASAP7_75t_L g1145 ( 
.A1(n_1019),
.A2(n_1057),
.B1(n_1029),
.B2(n_1014),
.C(n_1027),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1044),
.B(n_958),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1074),
.A2(n_826),
.B(n_914),
.C(n_969),
.Y(n_1147)
);

CKINVDCx6p67_ASAP7_75t_R g1148 ( 
.A(n_1035),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_984),
.B(n_958),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1032),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_SL g1151 ( 
.A1(n_1078),
.A2(n_819),
.B(n_822),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1068),
.B(n_958),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_976),
.B(n_904),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1078),
.A2(n_958),
.B(n_947),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1018),
.B(n_824),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_1082),
.B(n_918),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1091),
.B(n_918),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_SL g1158 ( 
.A1(n_1060),
.A2(n_969),
.B(n_918),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_987),
.A2(n_825),
.B(n_817),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1007),
.A2(n_811),
.B(n_914),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1060),
.B(n_911),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_981),
.B(n_911),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_988),
.B(n_817),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1002),
.A2(n_811),
.B(n_917),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1046),
.A2(n_910),
.B1(n_929),
.B2(n_933),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_972),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1002),
.A2(n_917),
.B(n_910),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1042),
.B(n_933),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_970),
.B(n_933),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1034),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1025),
.A2(n_1067),
.B(n_1007),
.C(n_1014),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1105),
.A2(n_910),
.B(n_929),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1047),
.B(n_910),
.Y(n_1173)
);

AOI221xp5_ASAP7_75t_L g1174 ( 
.A1(n_1057),
.A2(n_929),
.B1(n_933),
.B2(n_1020),
.C(n_1016),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_987),
.A2(n_929),
.B(n_1105),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1093),
.A2(n_1053),
.B(n_992),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1062),
.Y(n_1177)
);

AOI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1096),
.A2(n_1101),
.B(n_1093),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_1067),
.B(n_1016),
.C(n_1051),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_992),
.A2(n_1065),
.B(n_1113),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_996),
.A2(n_1045),
.B(n_991),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1085),
.A2(n_1015),
.B(n_1115),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_SL g1183 ( 
.A1(n_1081),
.A2(n_1066),
.B(n_1017),
.Y(n_1183)
);

AOI21x1_ASAP7_75t_SL g1184 ( 
.A1(n_1037),
.A2(n_1094),
.B(n_1073),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1045),
.A2(n_997),
.B(n_1079),
.Y(n_1185)
);

BUFx4f_ASAP7_75t_L g1186 ( 
.A(n_973),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1083),
.A2(n_994),
.B(n_1004),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_L g1188 ( 
.A(n_1005),
.B(n_1030),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_994),
.A2(n_1052),
.B(n_1069),
.Y(n_1189)
);

AOI221x1_ASAP7_75t_L g1190 ( 
.A1(n_1063),
.A2(n_1021),
.B1(n_1023),
.B2(n_1039),
.C(n_1017),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1031),
.A2(n_1036),
.B(n_982),
.C(n_999),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1052),
.A2(n_974),
.B(n_1038),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1070),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1061),
.B(n_1005),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1008),
.B(n_1026),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1087),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1088),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1095),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1049),
.A2(n_1051),
.B(n_1075),
.Y(n_1199)
);

O2A1O1Ixp5_ASAP7_75t_L g1200 ( 
.A1(n_1076),
.A2(n_1072),
.B(n_1086),
.C(n_1102),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1080),
.A2(n_1079),
.B(n_1012),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1097),
.A2(n_1103),
.A3(n_1107),
.B(n_990),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1049),
.A2(n_1000),
.B(n_1106),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1008),
.A2(n_1026),
.B(n_1099),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_SL g1205 ( 
.A(n_995),
.B(n_1098),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1066),
.A2(n_1110),
.B(n_1099),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1056),
.A2(n_986),
.B1(n_1048),
.B2(n_1089),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1013),
.A2(n_1050),
.B(n_985),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_985),
.A2(n_989),
.B(n_1001),
.Y(n_1209)
);

O2A1O1Ixp5_ASAP7_75t_L g1210 ( 
.A1(n_1086),
.A2(n_1094),
.B(n_1110),
.C(n_989),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1109),
.A2(n_1104),
.B(n_1043),
.C(n_1058),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_1058),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1092),
.A2(n_1112),
.B(n_1058),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1112),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_980),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1092),
.B(n_980),
.Y(n_1216)
);

INVxp67_ASAP7_75t_L g1217 ( 
.A(n_1048),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1006),
.B(n_1048),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_980),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1017),
.B(n_812),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_L g1221 ( 
.A1(n_975),
.A2(n_971),
.B(n_1100),
.Y(n_1221)
);

O2A1O1Ixp5_ASAP7_75t_L g1222 ( 
.A1(n_978),
.A2(n_882),
.B(n_1074),
.C(n_987),
.Y(n_1222)
);

OA22x2_ASAP7_75t_L g1223 ( 
.A1(n_1009),
.A2(n_698),
.B1(n_572),
.B2(n_1046),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_979),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1071),
.A2(n_1100),
.A3(n_1055),
.B(n_1096),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1054),
.A2(n_463),
.B(n_870),
.C(n_829),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1100),
.A2(n_1111),
.B(n_1108),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1009),
.A2(n_546),
.B1(n_508),
.B2(n_559),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1111),
.A2(n_975),
.B(n_1100),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1100),
.A2(n_1111),
.B(n_1108),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1054),
.A2(n_975),
.B(n_1084),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_979),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1054),
.A2(n_463),
.B(n_870),
.C(n_829),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1055),
.A2(n_1041),
.B(n_975),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1040),
.B(n_1054),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1054),
.A2(n_975),
.B(n_1084),
.Y(n_1236)
);

AO21x1_ASAP7_75t_L g1237 ( 
.A1(n_978),
.A2(n_1078),
.B(n_1041),
.Y(n_1237)
);

AOI21xp33_ASAP7_75t_L g1238 ( 
.A1(n_1014),
.A2(n_978),
.B(n_787),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1055),
.A2(n_1078),
.B(n_786),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1100),
.A2(n_1111),
.B(n_1108),
.Y(n_1240)
);

AO21x2_ASAP7_75t_L g1241 ( 
.A1(n_1100),
.A2(n_1055),
.B(n_1090),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_977),
.B(n_647),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1040),
.B(n_1054),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1100),
.A2(n_1111),
.B(n_1108),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1100),
.A2(n_1111),
.B(n_1108),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1055),
.A2(n_1078),
.B(n_786),
.Y(n_1246)
);

NOR2xp67_ASAP7_75t_L g1247 ( 
.A(n_1005),
.B(n_795),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1040),
.B(n_1054),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_983),
.A2(n_612),
.B(n_927),
.C(n_1025),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1055),
.A2(n_1041),
.B(n_975),
.Y(n_1250)
);

NAND2x1_ASAP7_75t_L g1251 ( 
.A(n_1066),
.B(n_1086),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1111),
.A2(n_975),
.B(n_1100),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1054),
.A2(n_975),
.B(n_1084),
.Y(n_1253)
);

NAND2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1081),
.B(n_812),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1100),
.A2(n_1111),
.B(n_1108),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1009),
.B(n_617),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1100),
.A2(n_1111),
.B(n_1108),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1058),
.Y(n_1258)
);

BUFx10_ASAP7_75t_L g1259 ( 
.A(n_1024),
.Y(n_1259)
);

OAI221xp5_ASAP7_75t_L g1260 ( 
.A1(n_1249),
.A2(n_1145),
.B1(n_1238),
.B2(n_1171),
.C(n_1228),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1142),
.B(n_1119),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1214),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1224),
.B(n_1232),
.Y(n_1263)
);

AO21x2_ASAP7_75t_L g1264 ( 
.A1(n_1181),
.A2(n_1237),
.B(n_1239),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1258),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1221),
.A2(n_1230),
.B(n_1227),
.Y(n_1266)
);

OR2x6_ASAP7_75t_L g1267 ( 
.A(n_1183),
.B(n_1158),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1242),
.B(n_1166),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1135),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1121),
.A2(n_1250),
.B(n_1234),
.Y(n_1270)
);

AOI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1175),
.A2(n_1246),
.B(n_1154),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1120),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1238),
.A2(n_1145),
.B(n_1233),
.C(n_1226),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1126),
.B(n_1118),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1141),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1223),
.A2(n_1163),
.B1(n_1132),
.B2(n_1256),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1121),
.A2(n_1234),
.B(n_1250),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1223),
.A2(n_1163),
.B1(n_1132),
.B2(n_1248),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1240),
.A2(n_1245),
.B(n_1257),
.Y(n_1279)
);

AOI221xp5_ASAP7_75t_L g1280 ( 
.A1(n_1124),
.A2(n_1235),
.B1(n_1243),
.B2(n_1248),
.C(n_1179),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1150),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_SL g1282 ( 
.A1(n_1235),
.A2(n_1243),
.B(n_1251),
.C(n_1174),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1220),
.B(n_1212),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1170),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1144),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1177),
.Y(n_1286)
);

AO32x2_ASAP7_75t_L g1287 ( 
.A1(n_1207),
.A2(n_1165),
.A3(n_1231),
.B1(n_1236),
.B2(n_1253),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1220),
.B(n_1212),
.Y(n_1288)
);

BUFx5_ASAP7_75t_L g1289 ( 
.A(n_1196),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1162),
.B(n_1138),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1118),
.A2(n_1207),
.B1(n_1220),
.B2(n_1127),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1217),
.B(n_1186),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1148),
.Y(n_1293)
);

NAND2x1p5_ASAP7_75t_L g1294 ( 
.A(n_1212),
.B(n_1213),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_1126),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1186),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1222),
.A2(n_1180),
.B(n_1147),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1244),
.A2(n_1255),
.B(n_1175),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1197),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1149),
.B(n_1157),
.Y(n_1300)
);

OA21x2_ASAP7_75t_L g1301 ( 
.A1(n_1176),
.A2(n_1231),
.B(n_1253),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1198),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1185),
.A2(n_1123),
.B(n_1143),
.Y(n_1303)
);

NOR2x1_ASAP7_75t_SL g1304 ( 
.A(n_1146),
.B(n_1156),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1155),
.B(n_1153),
.Y(n_1305)
);

AOI21xp33_ASAP7_75t_L g1306 ( 
.A1(n_1199),
.A2(n_1174),
.B(n_1160),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1193),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1130),
.A2(n_1117),
.B(n_1116),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1259),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1218),
.B(n_1259),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1136),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1136),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1160),
.A2(n_1151),
.B(n_1152),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1236),
.A2(n_1133),
.B(n_1131),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1152),
.A2(n_1178),
.B(n_1149),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1258),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1133),
.A2(n_1190),
.B(n_1164),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_SL g1318 ( 
.A1(n_1206),
.A2(n_1191),
.B(n_1159),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1125),
.A2(n_1199),
.B1(n_1203),
.B2(n_1254),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1157),
.Y(n_1320)
);

AO21x2_ASAP7_75t_L g1321 ( 
.A1(n_1178),
.A2(n_1192),
.B(n_1187),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1139),
.A2(n_1172),
.B(n_1167),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1169),
.B(n_1161),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_1161),
.Y(n_1324)
);

BUFx2_ASAP7_75t_R g1325 ( 
.A(n_1216),
.Y(n_1325)
);

AOI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1205),
.A2(n_1203),
.B1(n_1146),
.B2(n_1129),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1194),
.B(n_1215),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1189),
.A2(n_1201),
.B(n_1140),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1254),
.B(n_1173),
.Y(n_1329)
);

INVx8_ASAP7_75t_L g1330 ( 
.A(n_1212),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1215),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1200),
.A2(n_1201),
.B(n_1140),
.C(n_1211),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1206),
.A2(n_1188),
.B1(n_1128),
.B2(n_1195),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1194),
.B(n_1258),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1209),
.A2(n_1195),
.B(n_1208),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1202),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1128),
.A2(n_1247),
.B1(n_1219),
.B2(n_1182),
.Y(n_1337)
);

AO21x2_ASAP7_75t_L g1338 ( 
.A1(n_1241),
.A2(n_1168),
.B(n_1134),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1165),
.A2(n_1252),
.B(n_1229),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1202),
.Y(n_1340)
);

INVx8_ASAP7_75t_L g1341 ( 
.A(n_1215),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1184),
.A2(n_1252),
.B(n_1229),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1204),
.A2(n_1137),
.B(n_1182),
.Y(n_1343)
);

BUFx4f_ASAP7_75t_L g1344 ( 
.A(n_1205),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1122),
.A2(n_1210),
.B(n_1129),
.Y(n_1345)
);

O2A1O1Ixp33_ASAP7_75t_SL g1346 ( 
.A1(n_1225),
.A2(n_1249),
.B(n_1171),
.C(n_1054),
.Y(n_1346)
);

AO31x2_ASAP7_75t_L g1347 ( 
.A1(n_1225),
.A2(n_1237),
.A3(n_1181),
.B(n_1239),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1223),
.A2(n_1009),
.B1(n_787),
.B2(n_1145),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_1126),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1256),
.B(n_1242),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1142),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1186),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1249),
.A2(n_1238),
.B(n_1222),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1135),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1223),
.A2(n_698),
.B1(n_787),
.B2(n_421),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1221),
.A2(n_1230),
.B(n_1227),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1228),
.A2(n_698),
.B1(n_543),
.B2(n_1242),
.Y(n_1357)
);

AOI222xp33_ASAP7_75t_L g1358 ( 
.A1(n_1256),
.A2(n_1009),
.B1(n_698),
.B2(n_787),
.C1(n_970),
.C2(n_404),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1135),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1221),
.A2(n_1230),
.B(n_1227),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1118),
.B(n_1235),
.Y(n_1361)
);

BUFx2_ASAP7_75t_SL g1362 ( 
.A(n_1144),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1221),
.A2(n_1230),
.B(n_1227),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1142),
.B(n_1119),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1221),
.A2(n_1230),
.B(n_1227),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1181),
.A2(n_1237),
.B(n_1239),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1135),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1135),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1228),
.A2(n_698),
.B1(n_543),
.B2(n_1242),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1249),
.B(n_1145),
.C(n_1171),
.Y(n_1370)
);

OAI21xp33_ASAP7_75t_L g1371 ( 
.A1(n_1249),
.A2(n_1171),
.B(n_1145),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1249),
.A2(n_1238),
.B(n_1171),
.C(n_1145),
.Y(n_1372)
);

INVx5_ASAP7_75t_L g1373 ( 
.A(n_1220),
.Y(n_1373)
);

OAI211xp5_ASAP7_75t_L g1374 ( 
.A1(n_1249),
.A2(n_1145),
.B(n_1019),
.C(n_1228),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1221),
.A2(n_1230),
.B(n_1227),
.Y(n_1375)
);

AOI21xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1249),
.A2(n_1233),
.B(n_1226),
.Y(n_1376)
);

AOI21xp33_ASAP7_75t_L g1377 ( 
.A1(n_1238),
.A2(n_1171),
.B(n_1223),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1181),
.A2(n_1237),
.B(n_1239),
.Y(n_1378)
);

INVx3_ASAP7_75t_SL g1379 ( 
.A(n_1148),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1142),
.Y(n_1380)
);

NAND2x1p5_ASAP7_75t_L g1381 ( 
.A(n_1212),
.B(n_812),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1281),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1350),
.B(n_1290),
.Y(n_1383)
);

NOR2xp67_ASAP7_75t_R g1384 ( 
.A(n_1309),
.B(n_1296),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1370),
.A2(n_1260),
.B1(n_1372),
.B2(n_1348),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1324),
.B(n_1320),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1287),
.B(n_1269),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1274),
.B(n_1323),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1275),
.Y(n_1389)
);

AOI21x1_ASAP7_75t_SL g1390 ( 
.A1(n_1351),
.A2(n_1380),
.B(n_1272),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1371),
.A2(n_1348),
.B(n_1370),
.C(n_1377),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1278),
.B(n_1295),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1278),
.B(n_1295),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1297),
.A2(n_1342),
.B(n_1303),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1349),
.B(n_1280),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1362),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1260),
.A2(n_1371),
.B1(n_1374),
.B2(n_1273),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1361),
.B(n_1276),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1357),
.B(n_1369),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1297),
.A2(n_1343),
.B(n_1317),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1305),
.B(n_1261),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1327),
.B(n_1364),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1263),
.B(n_1300),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1361),
.B(n_1276),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1357),
.A2(n_1369),
.B1(n_1355),
.B2(n_1344),
.Y(n_1405)
);

CKINVDCx11_ASAP7_75t_R g1406 ( 
.A(n_1293),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1376),
.A2(n_1377),
.B(n_1353),
.C(n_1346),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1262),
.B(n_1284),
.Y(n_1408)
);

NAND4xp25_ASAP7_75t_L g1409 ( 
.A(n_1376),
.B(n_1358),
.C(n_1353),
.D(n_1268),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1311),
.B(n_1312),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1373),
.B(n_1267),
.Y(n_1411)
);

INVx3_ASAP7_75t_SL g1412 ( 
.A(n_1379),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1300),
.B(n_1286),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1287),
.B(n_1354),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1359),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1344),
.B(n_1326),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1367),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1368),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1317),
.A2(n_1356),
.B(n_1365),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1373),
.B(n_1267),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1291),
.A2(n_1306),
.B1(n_1326),
.B2(n_1352),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1291),
.B(n_1334),
.Y(n_1422)
);

CKINVDCx6p67_ASAP7_75t_R g1423 ( 
.A(n_1285),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1299),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1265),
.B(n_1316),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1302),
.B(n_1329),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1307),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1292),
.B(n_1287),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1331),
.B(n_1310),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1338),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1306),
.A2(n_1319),
.B1(n_1332),
.B2(n_1373),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1304),
.B(n_1325),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1325),
.B(n_1288),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1358),
.A2(n_1282),
.B(n_1318),
.C(n_1319),
.Y(n_1434)
);

CKINVDCx11_ASAP7_75t_R g1435 ( 
.A(n_1341),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1283),
.B(n_1289),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1341),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1264),
.A2(n_1366),
.B(n_1378),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1267),
.A2(n_1337),
.B(n_1333),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1333),
.A2(n_1381),
.B1(n_1345),
.B2(n_1301),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1345),
.A2(n_1337),
.B(n_1264),
.C(n_1378),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1266),
.A2(n_1363),
.B(n_1360),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1366),
.A2(n_1277),
.B(n_1270),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1313),
.B(n_1315),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1336),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1381),
.A2(n_1301),
.B1(n_1314),
.B2(n_1328),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1338),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1328),
.A2(n_1294),
.B1(n_1330),
.B2(n_1335),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1340),
.B(n_1321),
.Y(n_1449)
);

OAI21xp33_ASAP7_75t_L g1450 ( 
.A1(n_1271),
.A2(n_1339),
.B(n_1308),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1321),
.B(n_1322),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1347),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1335),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1270),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1298),
.A2(n_1279),
.B1(n_1375),
.B2(n_1370),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1287),
.B(n_1269),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1338),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1281),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1269),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1350),
.B(n_1290),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1350),
.B(n_1290),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1278),
.B(n_1295),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_SL g1463 ( 
.A1(n_1372),
.A2(n_1171),
.B(n_1267),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1278),
.B(n_1295),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1290),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1350),
.B(n_1290),
.Y(n_1466)
);

A2O1A1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1371),
.A2(n_1348),
.B(n_1370),
.C(n_1238),
.Y(n_1467)
);

AOI21x1_ASAP7_75t_SL g1468 ( 
.A1(n_1351),
.A2(n_1243),
.B(n_1235),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1269),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_SL g1470 ( 
.A1(n_1357),
.A2(n_1369),
.B1(n_1260),
.B2(n_1355),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1370),
.A2(n_1260),
.B1(n_1372),
.B2(n_1249),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1451),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1443),
.A2(n_1438),
.B(n_1450),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1424),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1386),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1436),
.B(n_1451),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1389),
.Y(n_1477)
);

AO21x2_ASAP7_75t_L g1478 ( 
.A1(n_1453),
.A2(n_1454),
.B(n_1430),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1415),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1387),
.B(n_1414),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1409),
.B(n_1397),
.Y(n_1481)
);

BUFx2_ASAP7_75t_SL g1482 ( 
.A(n_1382),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1387),
.B(n_1414),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1417),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1439),
.B(n_1411),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1456),
.B(n_1400),
.Y(n_1486)
);

AO21x2_ASAP7_75t_L g1487 ( 
.A1(n_1430),
.A2(n_1447),
.B(n_1457),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1456),
.B(n_1413),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1428),
.B(n_1403),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1394),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1418),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1439),
.B(n_1411),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1386),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1394),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1444),
.A2(n_1441),
.B(n_1446),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1400),
.B(n_1452),
.Y(n_1496)
);

AND2x4_ASAP7_75t_SL g1497 ( 
.A(n_1420),
.B(n_1386),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1394),
.Y(n_1498)
);

AO21x2_ASAP7_75t_L g1499 ( 
.A1(n_1431),
.A2(n_1399),
.B(n_1421),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1471),
.B(n_1385),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1400),
.Y(n_1501)
);

AO21x2_ASAP7_75t_L g1502 ( 
.A1(n_1449),
.A2(n_1391),
.B(n_1399),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1419),
.B(n_1459),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1401),
.B(n_1398),
.Y(n_1504)
);

OR2x6_ASAP7_75t_L g1505 ( 
.A(n_1420),
.B(n_1434),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1449),
.A2(n_1455),
.B(n_1404),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1467),
.A2(n_1391),
.B(n_1407),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1469),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1445),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1419),
.Y(n_1510)
);

AOI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1448),
.A2(n_1440),
.B(n_1442),
.Y(n_1511)
);

OAI21xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1463),
.A2(n_1416),
.B(n_1405),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1410),
.B(n_1462),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1392),
.B(n_1464),
.Y(n_1514)
);

AOI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1470),
.A2(n_1467),
.B1(n_1463),
.B2(n_1395),
.C(n_1393),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1427),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1408),
.B(n_1402),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1442),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1406),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1388),
.B(n_1465),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1483),
.B(n_1426),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1486),
.B(n_1442),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1500),
.A2(n_1383),
.B1(n_1466),
.B2(n_1461),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1503),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1486),
.B(n_1460),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1508),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1472),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1480),
.B(n_1425),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1480),
.B(n_1422),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1480),
.B(n_1429),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1503),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1496),
.B(n_1382),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1509),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1509),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1488),
.B(n_1458),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1518),
.Y(n_1536)
);

INVx4_ASAP7_75t_L g1537 ( 
.A(n_1485),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1478),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1496),
.B(n_1432),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1508),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1500),
.B(n_1423),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1513),
.B(n_1384),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1481),
.A2(n_1433),
.B1(n_1406),
.B2(n_1423),
.Y(n_1543)
);

AO21x2_ASAP7_75t_L g1544 ( 
.A1(n_1501),
.A2(n_1468),
.B(n_1390),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1474),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1478),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1496),
.B(n_1412),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1507),
.A2(n_1396),
.B(n_1437),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1472),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1535),
.Y(n_1550)
);

CKINVDCx16_ASAP7_75t_R g1551 ( 
.A(n_1547),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1543),
.A2(n_1507),
.B1(n_1515),
.B2(n_1481),
.Y(n_1552)
);

NOR4xp25_ASAP7_75t_SL g1553 ( 
.A(n_1527),
.B(n_1519),
.C(n_1510),
.D(n_1396),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1533),
.Y(n_1554)
);

OAI33xp33_ASAP7_75t_L g1555 ( 
.A1(n_1523),
.A2(n_1513),
.A3(n_1514),
.B1(n_1520),
.B2(n_1504),
.B3(n_1484),
.Y(n_1555)
);

AO21x2_ASAP7_75t_L g1556 ( 
.A1(n_1538),
.A2(n_1511),
.B(n_1495),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1533),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1538),
.A2(n_1511),
.B(n_1495),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1533),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1525),
.B(n_1476),
.Y(n_1560)
);

OAI221xp5_ASAP7_75t_L g1561 ( 
.A1(n_1542),
.A2(n_1512),
.B1(n_1515),
.B2(n_1514),
.C(n_1506),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1525),
.B(n_1476),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1547),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1541),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1542),
.B(n_1512),
.C(n_1506),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1523),
.A2(n_1499),
.B1(n_1502),
.B2(n_1505),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1535),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1534),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1534),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1545),
.Y(n_1570)
);

AOI221xp5_ASAP7_75t_SL g1571 ( 
.A1(n_1547),
.A2(n_1517),
.B1(n_1482),
.B2(n_1484),
.C(n_1477),
.Y(n_1571)
);

AOI211xp5_ASAP7_75t_L g1572 ( 
.A1(n_1548),
.A2(n_1510),
.B(n_1501),
.C(n_1514),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1530),
.B(n_1497),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_R g1574 ( 
.A(n_1543),
.B(n_1412),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1545),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1548),
.A2(n_1505),
.B1(n_1493),
.B2(n_1475),
.Y(n_1576)
);

NAND2xp33_ASAP7_75t_SL g1577 ( 
.A(n_1530),
.B(n_1499),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_R g1578 ( 
.A(n_1539),
.B(n_1506),
.Y(n_1578)
);

AOI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1522),
.A2(n_1499),
.B1(n_1502),
.B2(n_1510),
.C(n_1495),
.Y(n_1579)
);

OAI211xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1526),
.A2(n_1490),
.B(n_1494),
.C(n_1498),
.Y(n_1580)
);

AOI222xp33_ASAP7_75t_L g1581 ( 
.A1(n_1522),
.A2(n_1489),
.B1(n_1520),
.B2(n_1516),
.C1(n_1502),
.C2(n_1491),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1521),
.B(n_1489),
.Y(n_1582)
);

OAI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1535),
.A2(n_1505),
.B1(n_1492),
.B2(n_1485),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1539),
.A2(n_1502),
.B1(n_1495),
.B2(n_1506),
.Y(n_1584)
);

AOI221xp5_ASAP7_75t_L g1585 ( 
.A1(n_1522),
.A2(n_1495),
.B1(n_1516),
.B2(n_1479),
.C(n_1491),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1532),
.B(n_1482),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1545),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_R g1588 ( 
.A(n_1532),
.B(n_1435),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1537),
.B(n_1485),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1554),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1557),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1559),
.Y(n_1592)
);

OA21x2_ASAP7_75t_L g1593 ( 
.A1(n_1579),
.A2(n_1585),
.B(n_1538),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1568),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1563),
.B(n_1549),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1569),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1563),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1560),
.B(n_1531),
.Y(n_1598)
);

NOR2x1p5_ASAP7_75t_L g1599 ( 
.A(n_1565),
.B(n_1537),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1551),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1570),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1575),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1562),
.B(n_1531),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1581),
.B(n_1526),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1587),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1556),
.Y(n_1606)
);

AO21x2_ASAP7_75t_L g1607 ( 
.A1(n_1558),
.A2(n_1546),
.B(n_1487),
.Y(n_1607)
);

NAND3xp33_ASAP7_75t_L g1608 ( 
.A(n_1552),
.B(n_1506),
.C(n_1540),
.Y(n_1608)
);

NAND3xp33_ASAP7_75t_L g1609 ( 
.A(n_1584),
.B(n_1540),
.C(n_1473),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1582),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1550),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1558),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1572),
.B(n_1525),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1573),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1567),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1561),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1589),
.Y(n_1617)
);

NOR2x1_ASAP7_75t_L g1618 ( 
.A(n_1580),
.B(n_1544),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1573),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1571),
.A2(n_1546),
.B(n_1536),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1578),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1600),
.B(n_1553),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1616),
.B(n_1530),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1611),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1600),
.B(n_1586),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1600),
.B(n_1613),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1616),
.B(n_1524),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1600),
.B(n_1586),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1590),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1604),
.B(n_1610),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1604),
.B(n_1577),
.Y(n_1631)
);

NAND5xp2_ASAP7_75t_SL g1632 ( 
.A(n_1613),
.B(n_1566),
.C(n_1574),
.D(n_1532),
.E(n_1588),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1620),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1620),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1590),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1591),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1599),
.B(n_1597),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1613),
.B(n_1528),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1614),
.B(n_1597),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1621),
.A2(n_1584),
.B1(n_1566),
.B2(n_1555),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1591),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1614),
.B(n_1597),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1607),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1614),
.B(n_1597),
.Y(n_1644)
);

OAI21xp33_ASAP7_75t_L g1645 ( 
.A1(n_1608),
.A2(n_1580),
.B(n_1576),
.Y(n_1645)
);

NOR2x1_ASAP7_75t_L g1646 ( 
.A(n_1608),
.B(n_1564),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1610),
.B(n_1611),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1615),
.B(n_1524),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1599),
.B(n_1529),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1619),
.B(n_1528),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1592),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1619),
.B(n_1598),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1592),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1609),
.B(n_1555),
.C(n_1583),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1593),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1620),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1605),
.B(n_1593),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1594),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1649),
.B(n_1620),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1647),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1624),
.B(n_1620),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1623),
.B(n_1596),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1647),
.Y(n_1663)
);

NAND2x1_ASAP7_75t_L g1664 ( 
.A(n_1649),
.B(n_1595),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1654),
.B(n_1605),
.Y(n_1665)
);

AND2x4_ASAP7_75t_SL g1666 ( 
.A(n_1625),
.B(n_1595),
.Y(n_1666)
);

OAI21xp33_ASAP7_75t_L g1667 ( 
.A1(n_1646),
.A2(n_1645),
.B(n_1640),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1627),
.B(n_1596),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1630),
.B(n_1601),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1630),
.B(n_1601),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1650),
.B(n_1605),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1650),
.B(n_1598),
.Y(n_1672)
);

NOR2x1p5_ASAP7_75t_L g1673 ( 
.A(n_1626),
.B(n_1609),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1652),
.B(n_1598),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1649),
.B(n_1595),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1652),
.B(n_1603),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1658),
.Y(n_1677)
);

AOI32xp33_ASAP7_75t_L g1678 ( 
.A1(n_1646),
.A2(n_1618),
.A3(n_1539),
.B1(n_1583),
.B2(n_1617),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1634),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1629),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1634),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1634),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1637),
.B(n_1618),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1657),
.B(n_1603),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1626),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1629),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1649),
.B(n_1638),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1648),
.B(n_1602),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1656),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1637),
.B(n_1595),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1638),
.B(n_1595),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1685),
.B(n_1655),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1682),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1667),
.A2(n_1631),
.B1(n_1656),
.B2(n_1645),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1665),
.Y(n_1695)
);

OAI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1661),
.A2(n_1631),
.B1(n_1634),
.B2(n_1633),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1660),
.B(n_1625),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1682),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1677),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1669),
.B(n_1635),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1687),
.B(n_1666),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1687),
.B(n_1639),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1682),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1666),
.B(n_1639),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1689),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1673),
.B(n_1642),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1689),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1680),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1670),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1663),
.B(n_1628),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1690),
.B(n_1642),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1690),
.B(n_1644),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1686),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1690),
.B(n_1644),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1688),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1662),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1705),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1705),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1704),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1695),
.B(n_1684),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1693),
.Y(n_1721)
);

OAI22xp33_ASAP7_75t_SL g1722 ( 
.A1(n_1694),
.A2(n_1633),
.B1(n_1664),
.B2(n_1683),
.Y(n_1722)
);

OAI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1694),
.A2(n_1633),
.B1(n_1593),
.B2(n_1681),
.Y(n_1723)
);

OAI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1692),
.A2(n_1678),
.B(n_1659),
.C(n_1679),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1696),
.A2(n_1683),
.B(n_1659),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1707),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1707),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1693),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1709),
.A2(n_1676),
.B1(n_1674),
.B2(n_1632),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1706),
.A2(n_1632),
.B(n_1683),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1700),
.Y(n_1731)
);

NAND4xp75_ASAP7_75t_L g1732 ( 
.A(n_1706),
.B(n_1593),
.C(n_1622),
.D(n_1679),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1697),
.B(n_1672),
.Y(n_1733)
);

AOI21xp33_ASAP7_75t_L g1734 ( 
.A1(n_1708),
.A2(n_1713),
.B(n_1698),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1700),
.Y(n_1735)
);

NAND2x1p5_ASAP7_75t_L g1736 ( 
.A(n_1719),
.B(n_1704),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1717),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1718),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1720),
.B(n_1716),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1731),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1723),
.B(n_1716),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1726),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1720),
.B(n_1710),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1732),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1735),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1727),
.Y(n_1746)
);

NAND4xp25_ASAP7_75t_L g1747 ( 
.A(n_1743),
.B(n_1730),
.C(n_1729),
.D(n_1734),
.Y(n_1747)
);

AOI32xp33_ASAP7_75t_L g1748 ( 
.A1(n_1741),
.A2(n_1723),
.A3(n_1739),
.B1(n_1746),
.B2(n_1745),
.Y(n_1748)
);

OAI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1744),
.A2(n_1724),
.B(n_1702),
.Y(n_1749)
);

INVxp67_ASAP7_75t_SL g1750 ( 
.A(n_1736),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_SL g1751 ( 
.A(n_1740),
.B(n_1701),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1737),
.Y(n_1752)
);

AOI21xp33_ASAP7_75t_L g1753 ( 
.A1(n_1741),
.A2(n_1722),
.B(n_1725),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1738),
.A2(n_1727),
.B(n_1699),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1742),
.A2(n_1728),
.B(n_1721),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1744),
.A2(n_1701),
.B(n_1712),
.Y(n_1756)
);

O2A1O1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1753),
.A2(n_1713),
.B(n_1708),
.C(n_1733),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1750),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1752),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_SL g1760 ( 
.A1(n_1748),
.A2(n_1693),
.B(n_1698),
.C(n_1703),
.Y(n_1760)
);

AOI222xp33_ASAP7_75t_L g1761 ( 
.A1(n_1749),
.A2(n_1715),
.B1(n_1681),
.B2(n_1643),
.C1(n_1612),
.C2(n_1606),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1758),
.B(n_1715),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1759),
.Y(n_1763)
);

NOR2x1_ASAP7_75t_L g1764 ( 
.A(n_1760),
.B(n_1747),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1757),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1761),
.B(n_1751),
.Y(n_1766)
);

NOR2x1_ASAP7_75t_L g1767 ( 
.A(n_1760),
.B(n_1754),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1767),
.B(n_1756),
.Y(n_1768)
);

OAI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1766),
.A2(n_1698),
.B1(n_1703),
.B2(n_1755),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1764),
.B(n_1702),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1763),
.B(n_1711),
.Y(n_1771)
);

OA22x2_ASAP7_75t_L g1772 ( 
.A1(n_1765),
.A2(n_1714),
.B1(n_1711),
.B2(n_1712),
.Y(n_1772)
);

NAND4xp75_ASAP7_75t_L g1773 ( 
.A(n_1768),
.B(n_1714),
.C(n_1762),
.D(n_1622),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1770),
.B(n_1769),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1771),
.B(n_1671),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1773),
.A2(n_1774),
.B(n_1772),
.Y(n_1776)
);

INVx4_ASAP7_75t_L g1777 ( 
.A(n_1776),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1777),
.B(n_1775),
.Y(n_1778)
);

XNOR2xp5_ASAP7_75t_L g1779 ( 
.A(n_1777),
.B(n_1693),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1778),
.Y(n_1780)
);

XNOR2x1_ASAP7_75t_L g1781 ( 
.A(n_1779),
.B(n_1637),
.Y(n_1781)
);

OAI22x1_ASAP7_75t_L g1782 ( 
.A1(n_1780),
.A2(n_1637),
.B1(n_1675),
.B2(n_1628),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1781),
.Y(n_1783)
);

NOR2x1_ASAP7_75t_L g1784 ( 
.A(n_1783),
.B(n_1675),
.Y(n_1784)
);

OAI21xp33_ASAP7_75t_L g1785 ( 
.A1(n_1784),
.A2(n_1782),
.B(n_1691),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1785),
.B(n_1668),
.Y(n_1786)
);

AO221x2_ASAP7_75t_L g1787 ( 
.A1(n_1786),
.A2(n_1636),
.B1(n_1635),
.B2(n_1641),
.C(n_1651),
.Y(n_1787)
);

AOI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1787),
.A2(n_1643),
.B1(n_1691),
.B2(n_1612),
.C(n_1606),
.Y(n_1788)
);

OAI31xp33_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1653),
.A3(n_1651),
.B(n_1641),
.Y(n_1789)
);


endmodule