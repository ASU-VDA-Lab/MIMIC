module fake_jpeg_6189_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_19),
.B(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_17),
.C(n_13),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_26),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_17),
.B(n_20),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_16),
.B(n_14),
.Y(n_47)
);

AND2x6_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_20),
.Y(n_37)
);

AND2x6_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_33),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_22),
.B(n_2),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_36),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_16),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_54),
.B1(n_55),
.B2(n_43),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_56),
.C(n_44),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_34),
.B1(n_32),
.B2(n_27),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_29),
.B1(n_35),
.B2(n_21),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_42),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_53),
.B1(n_14),
.B2(n_2),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_59),
.B(n_3),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_61),
.Y(n_63)
);

AOI322xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_46),
.A3(n_49),
.B1(n_40),
.B2(n_48),
.C1(n_21),
.C2(n_29),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_56),
.C(n_52),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_65),
.B(n_7),
.Y(n_67)
);

AOI31xp67_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_1),
.A3(n_3),
.B(n_4),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_63),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_69),
.A2(n_62),
.B(n_60),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_68),
.B(n_7),
.Y(n_71)
);


endmodule