module fake_jpeg_29193_n_158 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_2),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_5),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_11),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_0),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_69),
.Y(n_79)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_2),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_3),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_57),
.Y(n_75)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_88),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_51),
.B1(n_54),
.B2(n_60),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_62),
.B1(n_5),
.B2(n_7),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_63),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_51),
.B1(n_54),
.B2(n_49),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_83),
.B1(n_61),
.B2(n_58),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_65),
.B1(n_52),
.B2(n_48),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_52),
.C(n_50),
.Y(n_88)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_98),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_62),
.B(n_55),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_4),
.B(n_7),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_99),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_62),
.B1(n_10),
.B2(n_8),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_81),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_86),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_104),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_117)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_4),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_23),
.B(n_24),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_116),
.B1(n_109),
.B2(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_14),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_22),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_125),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_16),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_17),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

BUFx2_ASAP7_75t_SL g142 ( 
.A(n_126),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_132),
.B1(n_140),
.B2(n_33),
.C(n_34),
.Y(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_138),
.B(n_30),
.C(n_31),
.D(n_32),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_36),
.B(n_38),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_25),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_125),
.C(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_26),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_145),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_146),
.A2(n_147),
.B(n_133),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_142),
.Y(n_148)
);

HAxp5_ASAP7_75t_SL g151 ( 
.A(n_148),
.B(n_142),
.CON(n_151),
.SN(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_139),
.C(n_128),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_152),
.B(n_137),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_143),
.B1(n_129),
.B2(n_141),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_126),
.A3(n_136),
.B1(n_127),
.B2(n_149),
.C1(n_124),
.C2(n_106),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_41),
.B(n_42),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_43),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_44),
.Y(n_158)
);


endmodule