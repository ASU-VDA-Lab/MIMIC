module fake_jpeg_22629_n_184 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_35),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx6p67_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_28),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_52),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_50),
.B1(n_19),
.B2(n_16),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_18),
.B1(n_21),
.B2(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_26),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_27),
.B(n_20),
.C(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_59),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_30),
.B1(n_21),
.B2(n_18),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_71),
.B1(n_72),
.B2(n_42),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_26),
.B1(n_24),
.B2(n_23),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_66),
.B(n_69),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_24),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_70),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_23),
.B1(n_20),
.B2(n_19),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_15),
.B1(n_28),
.B2(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_79),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_61),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_49),
.B1(n_53),
.B2(n_46),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_84),
.B1(n_92),
.B2(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_88),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_46),
.B1(n_51),
.B2(n_47),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_51),
.B1(n_47),
.B2(n_38),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_70),
.B1(n_68),
.B2(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_44),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_48),
.C(n_45),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_60),
.B(n_65),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_109),
.B(n_81),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_98),
.B1(n_105),
.B2(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_99),
.B(n_106),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_45),
.B1(n_57),
.B2(n_15),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_78),
.C(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_75),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_57),
.B1(n_15),
.B2(n_28),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_83),
.B1(n_90),
.B2(n_13),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_58),
.B(n_2),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_77),
.B(n_85),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_1),
.B(n_2),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_116),
.B(n_120),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_80),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_118),
.B(n_97),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_78),
.B1(n_92),
.B2(n_84),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_115),
.B1(n_117),
.B2(n_3),
.Y(n_136)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_120),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_82),
.B1(n_75),
.B2(n_83),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_98),
.B1(n_94),
.B2(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_3),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_106),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_128),
.C(n_132),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

AOI221xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_101),
.B1(n_109),
.B2(n_99),
.C(n_104),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_111),
.A3(n_118),
.B1(n_116),
.B2(n_122),
.C1(n_125),
.C2(n_114),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_104),
.B(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_135),
.B(n_123),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_139),
.B1(n_119),
.B2(n_124),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_117),
.Y(n_145)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_142),
.A2(n_146),
.B1(n_133),
.B2(n_137),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_145),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_132),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_135),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_115),
.C(n_13),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_138),
.C(n_127),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_151),
.B(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_159),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_157),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_149),
.B(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_147),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_166),
.B(n_5),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_156),
.C(n_153),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_150),
.C(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_4),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_171),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_7),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_172),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_5),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_6),
.Y(n_172)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

AOI21x1_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_171),
.B(n_165),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_179),
.C(n_8),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_7),
.B(n_8),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_175),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_181),
.B(n_9),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_10),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_11),
.Y(n_184)
);


endmodule