module real_jpeg_17738_n_5 (n_4, n_0, n_1, n_2, n_3, n_5);

input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_5;

wire n_17;
wire n_12;
wire n_8;
wire n_18;
wire n_10;
wire n_11;
wire n_14;
wire n_15;
wire n_6;
wire n_7;
wire n_16;
wire n_13;
wire n_9;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_9),
.Y(n_8)
);

OR2x4_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_9),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_16),
.Y(n_15)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_16),
.Y(n_17)
);

INVx13_ASAP7_75t_SL g5 ( 
.A(n_6),
.Y(n_5)
);

AOI22xp5_ASAP7_75t_SL g6 ( 
.A1(n_7),
.A2(n_12),
.B1(n_13),
.B2(n_18),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_10),
.Y(n_7)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NAND3xp33_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_15),
.C(n_17),
.Y(n_13)
);


endmodule