module fake_aes_10323_n_627 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_627);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_627;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_73), .Y(n_74) );
BUFx6f_ASAP7_75t_L g75 ( .A(n_34), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_51), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_5), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_71), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_35), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_23), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_68), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_29), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_38), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_37), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_33), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_57), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_25), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_66), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_27), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_41), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_70), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_62), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_72), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_59), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_69), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_14), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_31), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_26), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_53), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_64), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_2), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_46), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_3), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_8), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_58), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_16), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_43), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_50), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_18), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_36), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_39), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_1), .Y(n_114) );
INVxp33_ASAP7_75t_SL g115 ( .A(n_60), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_65), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_55), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_13), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_110), .Y(n_120) );
NOR2x1_ASAP7_75t_L g121 ( .A(n_110), .B(n_0), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_74), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_76), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_80), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_99), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_91), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_93), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
CKINVDCx11_ASAP7_75t_R g130 ( .A(n_79), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_77), .B(n_0), .Y(n_131) );
BUFx3_ASAP7_75t_L g132 ( .A(n_99), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_77), .B(n_1), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_93), .B(n_2), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_82), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
BUFx8_ASAP7_75t_L g139 ( .A(n_75), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_75), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_88), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_88), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_75), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_96), .B(n_3), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_89), .B(n_22), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_96), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_89), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g150 ( .A1(n_104), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_92), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_95), .B(n_28), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_95), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_97), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_97), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_75), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_107), .B(n_7), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_124), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_124), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_127), .B(n_94), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_127), .B(n_94), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_119), .B(n_85), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_124), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
INVxp67_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g167 ( .A1(n_128), .A2(n_107), .B1(n_111), .B2(n_105), .Y(n_167) );
BUFx4f_ASAP7_75t_L g168 ( .A(n_147), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_119), .B(n_103), .Y(n_170) );
INVx8_ASAP7_75t_L g171 ( .A(n_147), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_122), .B(n_101), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_124), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_125), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_125), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_148), .B(n_111), .Y(n_182) );
BUFx4f_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
OR2x2_ASAP7_75t_L g184 ( .A(n_148), .B(n_114), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_125), .B(n_102), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_129), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_129), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_129), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_122), .B(n_118), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_129), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_123), .B(n_117), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_123), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_151), .A2(n_87), .B1(n_115), .B2(n_100), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
BUFx10_ASAP7_75t_L g198 ( .A(n_147), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_134), .B(n_81), .Y(n_199) );
INVxp67_ASAP7_75t_L g200 ( .A(n_134), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_136), .B(n_113), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_132), .Y(n_202) );
NOR2x1p5_ASAP7_75t_L g203 ( .A(n_130), .B(n_84), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_139), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_137), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
OAI22xp33_ASAP7_75t_SL g207 ( .A1(n_151), .A2(n_116), .B1(n_98), .B2(n_109), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_139), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_136), .B(n_116), .Y(n_209) );
INVxp67_ASAP7_75t_SL g210 ( .A(n_137), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_138), .B(n_108), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_137), .B(n_100), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_163), .B(n_138), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_191), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_200), .B(n_142), .Y(n_215) );
NAND2xp33_ASAP7_75t_SL g216 ( .A(n_187), .B(n_140), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_191), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_184), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_191), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_205), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_205), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_185), .B(n_157), .Y(n_222) );
CKINVDCx8_ASAP7_75t_R g223 ( .A(n_169), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_182), .B(n_121), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_205), .Y(n_225) );
OR2x6_ASAP7_75t_L g226 ( .A(n_171), .B(n_150), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_185), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_166), .A2(n_150), .B1(n_155), .B2(n_142), .Y(n_228) );
NOR2xp33_ASAP7_75t_SL g229 ( .A(n_187), .B(n_152), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_208), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_212), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_182), .A2(n_147), .B1(n_152), .B2(n_140), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_159), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_184), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_195), .B(n_144), .Y(n_235) );
INVx1_ASAP7_75t_SL g236 ( .A(n_169), .Y(n_236) );
NAND2x1p5_ASAP7_75t_L g237 ( .A(n_187), .B(n_149), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_159), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_182), .B(n_144), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_196), .A2(n_162), .B1(n_161), .B2(n_182), .Y(n_240) );
AND3x1_ASAP7_75t_L g241 ( .A(n_196), .B(n_157), .C(n_131), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_208), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_212), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_170), .B(n_155), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_210), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_160), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_160), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_164), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_171), .Y(n_249) );
INVxp67_ASAP7_75t_SL g250 ( .A(n_164), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_172), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_167), .A2(n_153), .B1(n_143), .B2(n_152), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_192), .A2(n_153), .B1(n_143), .B2(n_152), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_194), .B(n_154), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_173), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_199), .B(n_211), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_192), .B(n_154), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_209), .B(n_154), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_212), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_173), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_186), .A2(n_152), .B1(n_147), .B2(n_154), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_209), .B(n_149), .Y(n_262) );
BUFx4f_ASAP7_75t_SL g263 ( .A(n_201), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_174), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_174), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_179), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_171), .A2(n_131), .B1(n_146), .B2(n_133), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_207), .A2(n_152), .B1(n_147), .B2(n_146), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_179), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_180), .A2(n_152), .B(n_149), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_238), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_224), .B(n_186), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_218), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_233), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_227), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_223), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_238), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_246), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_SL g279 ( .A1(n_270), .A2(n_193), .B(n_188), .C(n_190), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_246), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_240), .A2(n_207), .B1(n_204), .B2(n_212), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_247), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_247), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_234), .B(n_213), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_264), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_264), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_231), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_224), .B(n_186), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_224), .B(n_186), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_241), .A2(n_204), .B1(n_203), .B2(n_190), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_237), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_236), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_231), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_257), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_251), .A2(n_203), .B1(n_180), .B2(n_188), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_237), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_266), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_231), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_239), .A2(n_133), .B(n_193), .C(n_149), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_223), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_266), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_237), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_243), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_233), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_243), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_269), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_263), .B(n_183), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_226), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_269), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_235), .B(n_171), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_248), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_267), .A2(n_183), .B1(n_168), .B2(n_171), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_230), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_243), .B(n_121), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_244), .B(n_168), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_313), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_273), .A2(n_226), .B1(n_259), .B2(n_228), .Y(n_317) );
OR2x6_ASAP7_75t_L g318 ( .A(n_296), .B(n_259), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_284), .A2(n_258), .B1(n_262), .B2(n_256), .C(n_120), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_273), .A2(n_226), .B1(n_259), .B2(n_245), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_292), .Y(n_321) );
O2A1O1Ixp33_ASAP7_75t_SL g322 ( .A1(n_271), .A2(n_278), .B(n_277), .C(n_280), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_313), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_L g324 ( .A1(n_284), .A2(n_299), .B(n_282), .C(n_297), .Y(n_324) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_281), .A2(n_226), .B1(n_268), .B2(n_252), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_296), .B(n_221), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_292), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_SL g328 ( .A1(n_271), .A2(n_254), .B(n_253), .C(n_242), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_277), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_274), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g331 ( .A1(n_308), .A2(n_215), .B1(n_137), .B2(n_229), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_274), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_276), .B(n_227), .Y(n_333) );
AOI332xp33_ASAP7_75t_L g334 ( .A1(n_290), .A2(n_120), .A3(n_109), .B1(n_102), .B2(n_98), .B3(n_112), .C1(n_78), .C2(n_232), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_272), .A2(n_216), .B1(n_221), .B2(n_225), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_278), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_280), .Y(n_337) );
AOI22xp33_ASAP7_75t_SL g338 ( .A1(n_276), .A2(n_120), .B1(n_152), .B2(n_250), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_304), .Y(n_339) );
OA21x2_ASAP7_75t_L g340 ( .A1(n_282), .A2(n_261), .B(n_112), .Y(n_340) );
OAI211xp5_ASAP7_75t_L g341 ( .A1(n_295), .A2(n_120), .B(n_222), .C(n_225), .Y(n_341) );
OA21x2_ASAP7_75t_L g342 ( .A1(n_283), .A2(n_78), .B(n_219), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_283), .Y(n_343) );
OAI222xp33_ASAP7_75t_L g344 ( .A1(n_325), .A2(n_300), .B1(n_302), .B2(n_294), .C1(n_286), .C2(n_297), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_325), .A2(n_291), .B1(n_302), .B2(n_286), .Y(n_345) );
CKINVDCx6p67_ASAP7_75t_R g346 ( .A(n_321), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_319), .A2(n_327), .B1(n_321), .B2(n_317), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_329), .B(n_272), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_331), .A2(n_285), .B1(n_306), .B2(n_301), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_327), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_329), .Y(n_351) );
NOR2x1_ASAP7_75t_SL g352 ( .A(n_318), .B(n_285), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_330), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_319), .A2(n_300), .B1(n_314), .B2(n_272), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_336), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_326), .Y(n_356) );
NAND4xp25_ASAP7_75t_L g357 ( .A(n_320), .B(n_314), .C(n_288), .D(n_272), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_318), .A2(n_301), .B1(n_306), .B2(n_309), .Y(n_358) );
AO21x2_ASAP7_75t_L g359 ( .A1(n_328), .A2(n_279), .B(n_309), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_331), .A2(n_314), .B1(n_289), .B2(n_288), .Y(n_360) );
NOR2xp67_ASAP7_75t_L g361 ( .A(n_316), .B(n_304), .Y(n_361) );
OR2x6_ASAP7_75t_L g362 ( .A(n_318), .B(n_326), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_318), .A2(n_312), .B1(n_310), .B2(n_275), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_336), .B(n_289), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_318), .A2(n_311), .B1(n_288), .B2(n_289), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_337), .B(n_289), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_318), .A2(n_311), .B1(n_315), .B2(n_275), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_316), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_337), .B(n_307), .Y(n_369) );
NAND2xp33_ASAP7_75t_R g370 ( .A(n_362), .B(n_342), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_353), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_362), .Y(n_372) );
OAI31xp33_ASAP7_75t_L g373 ( .A1(n_344), .A2(n_341), .A3(n_324), .B(n_343), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_353), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_353), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_351), .B(n_343), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_351), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_355), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_347), .A2(n_324), .B1(n_322), .B2(n_341), .C(n_333), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_355), .B(n_330), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_349), .A2(n_339), .B(n_330), .Y(n_381) );
OAI21xp5_ASAP7_75t_SL g382 ( .A1(n_357), .A2(n_338), .B(n_335), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_352), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g385 ( .A1(n_354), .A2(n_338), .B1(n_303), .B2(n_305), .C(n_287), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_350), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_349), .A2(n_326), .B1(n_298), .B2(n_287), .C(n_293), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_362), .B(n_332), .Y(n_388) );
NAND4xp25_ASAP7_75t_L g389 ( .A(n_357), .B(n_132), .C(n_126), .D(n_334), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_362), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_359), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_352), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_346), .Y(n_393) );
OAI31xp33_ASAP7_75t_L g394 ( .A1(n_365), .A2(n_315), .A3(n_326), .B(n_216), .Y(n_394) );
OA21x2_ASAP7_75t_L g395 ( .A1(n_360), .A2(n_339), .B(n_332), .Y(n_395) );
NAND3xp33_ASAP7_75t_L g396 ( .A(n_365), .B(n_342), .C(n_340), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_346), .A2(n_334), .B1(n_339), .B2(n_332), .Y(n_397) );
AOI21xp5_ASAP7_75t_SL g398 ( .A1(n_367), .A2(n_342), .B(n_340), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_348), .B(n_342), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_356), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_358), .A2(n_323), .B1(n_316), .B2(n_342), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_348), .B(n_287), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_377), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_397), .A2(n_345), .B1(n_367), .B2(n_356), .Y(n_404) );
BUFx2_ASAP7_75t_SL g405 ( .A(n_383), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_377), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_382), .A2(n_363), .B1(n_369), .B2(n_361), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_377), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_378), .B(n_368), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_371), .Y(n_411) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_375), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_393), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_382), .A2(n_366), .B1(n_364), .B2(n_361), .C(n_106), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_386), .B(n_364), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_378), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_392), .B(n_368), .Y(n_418) );
OAI31xp33_ASAP7_75t_L g419 ( .A1(n_389), .A2(n_366), .A3(n_368), .B(n_323), .Y(n_419) );
NAND4xp25_ASAP7_75t_L g420 ( .A(n_373), .B(n_132), .C(n_126), .D(n_368), .Y(n_420) );
AO21x2_ASAP7_75t_L g421 ( .A1(n_396), .A2(n_359), .B(n_219), .Y(n_421) );
OAI31xp33_ASAP7_75t_L g422 ( .A1(n_389), .A2(n_323), .A3(n_316), .B(n_293), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_399), .B(n_323), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_371), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_379), .A2(n_126), .B1(n_75), .B2(n_305), .C(n_298), .Y(n_425) );
OAI211xp5_ASAP7_75t_SL g426 ( .A1(n_373), .A2(n_165), .B(n_175), .C(n_176), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_371), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_394), .B(n_139), .C(n_145), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_399), .B(n_340), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_374), .B(n_340), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_374), .Y(n_431) );
AOI33xp33_ASAP7_75t_L g432 ( .A1(n_392), .A2(n_175), .A3(n_176), .B1(n_177), .B2(n_178), .B3(n_181), .Y(n_432) );
INVx4_ASAP7_75t_L g433 ( .A(n_375), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_374), .B(n_340), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_375), .Y(n_435) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_375), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_380), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_376), .A2(n_126), .B1(n_305), .B2(n_298), .C(n_293), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_394), .A2(n_359), .B1(n_313), .B2(n_183), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_388), .B(n_8), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_400), .Y(n_441) );
NOR3xp33_ASAP7_75t_L g442 ( .A(n_385), .B(n_221), .C(n_90), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_388), .B(n_9), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_390), .Y(n_444) );
AOI21xp33_ASAP7_75t_L g445 ( .A1(n_370), .A2(n_313), .B(n_202), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_391), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_398), .A2(n_168), .B(n_313), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_372), .B(n_9), .Y(n_448) );
OAI33xp33_ASAP7_75t_L g449 ( .A1(n_401), .A2(n_10), .A3(n_11), .B1(n_12), .B2(n_14), .B3(n_15), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g450 ( .A(n_408), .B(n_390), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_403), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_423), .B(n_384), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_423), .B(n_384), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_442), .B(n_145), .C(n_396), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_429), .B(n_372), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_408), .B(n_390), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_418), .B(n_400), .Y(n_458) );
NOR3xp33_ASAP7_75t_L g459 ( .A(n_449), .B(n_387), .C(n_402), .Y(n_459) );
AO21x1_ASAP7_75t_L g460 ( .A1(n_407), .A2(n_381), .B(n_391), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_429), .B(n_406), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_406), .B(n_395), .Y(n_462) );
AOI322xp5_ASAP7_75t_L g463 ( .A1(n_448), .A2(n_400), .A3(n_11), .B1(n_15), .B2(n_16), .C1(n_17), .C2(n_18), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_409), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_417), .B(n_395), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_417), .B(n_395), .Y(n_466) );
NAND2x1_ASAP7_75t_L g467 ( .A(n_433), .B(n_418), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_413), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_418), .B(n_391), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_424), .B(n_398), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_416), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_440), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_411), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_424), .B(n_10), .Y(n_474) );
INVx1_ASAP7_75t_SL g475 ( .A(n_414), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_437), .B(n_17), .Y(n_476) );
NAND2xp33_ASAP7_75t_SL g477 ( .A(n_444), .B(n_230), .Y(n_477) );
AND3x1_ASAP7_75t_L g478 ( .A(n_419), .B(n_19), .C(n_20), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_437), .B(n_265), .Y(n_479) );
OAI211xp5_ASAP7_75t_SL g480 ( .A1(n_415), .A2(n_165), .B(n_178), .C(n_181), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_411), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_428), .A2(n_217), .B1(n_220), .B2(n_214), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_427), .B(n_177), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_422), .B(n_158), .C(n_206), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_427), .B(n_21), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_404), .A2(n_214), .B1(n_217), .B2(n_220), .Y(n_487) );
OAI33xp33_ASAP7_75t_L g488 ( .A1(n_410), .A2(n_197), .A3(n_189), .B1(n_255), .B2(n_248), .B3(n_265), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_410), .Y(n_489) );
AOI211x1_ASAP7_75t_L g490 ( .A1(n_448), .A2(n_24), .B(n_30), .C(n_32), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_443), .B(n_260), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_443), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_431), .B(n_40), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_431), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_435), .B(n_42), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_405), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_433), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_405), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_446), .Y(n_499) );
AOI21xp33_ASAP7_75t_SL g500 ( .A1(n_441), .A2(n_44), .B(n_45), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_444), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_441), .B(n_202), .Y(n_502) );
INVx2_ASAP7_75t_SL g503 ( .A(n_433), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_471), .B(n_412), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_501), .B(n_436), .Y(n_505) );
AND2x4_ASAP7_75t_SL g506 ( .A(n_498), .B(n_435), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_453), .B(n_434), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_451), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_452), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_468), .Y(n_510) );
AOI322xp5_ASAP7_75t_L g511 ( .A1(n_472), .A2(n_439), .A3(n_425), .B1(n_434), .B2(n_430), .C1(n_446), .C2(n_445), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_494), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_464), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_453), .B(n_430), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_476), .A2(n_420), .B(n_426), .C(n_447), .Y(n_515) );
AOI21xp33_ASAP7_75t_L g516 ( .A1(n_474), .A2(n_421), .B(n_438), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_461), .B(n_421), .Y(n_517) );
NAND4xp75_ASAP7_75t_SL g518 ( .A(n_478), .B(n_432), .C(n_48), .D(n_49), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_499), .Y(n_519) );
AOI221x1_ASAP7_75t_SL g520 ( .A1(n_492), .A2(n_421), .B1(n_197), .B2(n_189), .C(n_56), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_455), .A2(n_242), .B(n_230), .Y(n_521) );
AND2x4_ASAP7_75t_SL g522 ( .A(n_497), .B(n_260), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_464), .Y(n_523) );
NOR2xp67_ASAP7_75t_L g524 ( .A(n_497), .B(n_47), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_489), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_461), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_483), .B(n_52), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_456), .B(n_54), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_475), .B(n_61), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_474), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_473), .Y(n_531) );
INVx3_ASAP7_75t_L g532 ( .A(n_467), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_454), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_456), .B(n_63), .Y(n_534) );
INVx3_ASAP7_75t_L g535 ( .A(n_497), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_485), .A2(n_255), .B(n_249), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_477), .A2(n_67), .B(n_249), .C(n_206), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_481), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_503), .B(n_158), .Y(n_539) );
INVx4_ASAP7_75t_L g540 ( .A(n_503), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_458), .B(n_206), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_457), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_496), .B(n_158), .Y(n_543) );
OAI31xp33_ASAP7_75t_L g544 ( .A1(n_477), .A2(n_158), .A3(n_206), .B(n_198), .Y(n_544) );
NOR3xp33_ASAP7_75t_L g545 ( .A(n_488), .B(n_158), .C(n_206), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_481), .B(n_198), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_450), .B(n_198), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_462), .B(n_198), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_465), .Y(n_549) );
AOI211x1_ASAP7_75t_L g550 ( .A1(n_520), .A2(n_460), .B(n_491), .C(n_463), .Y(n_550) );
NOR2x1_ASAP7_75t_L g551 ( .A(n_540), .B(n_493), .Y(n_551) );
HB1xp67_ASAP7_75t_SL g552 ( .A(n_540), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_526), .B(n_470), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_540), .A2(n_459), .B1(n_457), .B2(n_460), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_510), .Y(n_555) );
XNOR2xp5_ASAP7_75t_L g556 ( .A(n_533), .B(n_458), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_531), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_532), .B(n_457), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_532), .B(n_450), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_535), .B(n_458), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_508), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g562 ( .A1(n_537), .A2(n_500), .B(n_479), .C(n_480), .Y(n_562) );
NOR2xp67_ASAP7_75t_L g563 ( .A(n_535), .B(n_470), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_507), .B(n_514), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_509), .Y(n_565) );
NAND4xp75_ASAP7_75t_L g566 ( .A(n_524), .B(n_490), .C(n_486), .D(n_493), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_512), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_545), .B(n_502), .C(n_482), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_522), .A2(n_487), .B1(n_502), .B2(n_469), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_525), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_542), .B(n_505), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_504), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_531), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_513), .Y(n_574) );
OA211x2_ASAP7_75t_L g575 ( .A1(n_536), .A2(n_486), .B(n_469), .C(n_495), .Y(n_575) );
XOR2xp5_ASAP7_75t_SL g576 ( .A(n_528), .B(n_465), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_523), .Y(n_577) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_518), .B(n_484), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_529), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_538), .Y(n_580) );
INVxp67_ASAP7_75t_L g581 ( .A(n_535), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_530), .A2(n_466), .B1(n_495), .B2(n_484), .Y(n_582) );
OAI21xp5_ASAP7_75t_SL g583 ( .A1(n_522), .A2(n_466), .B(n_506), .Y(n_583) );
XNOR2x1_ASAP7_75t_L g584 ( .A(n_518), .B(n_534), .Y(n_584) );
OA22x2_ASAP7_75t_L g585 ( .A1(n_506), .A2(n_527), .B1(n_519), .B2(n_521), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_517), .B(n_511), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_545), .B(n_516), .C(n_537), .Y(n_587) );
OAI211xp5_ASAP7_75t_SL g588 ( .A1(n_515), .A2(n_543), .B(n_544), .C(n_539), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_541), .B(n_515), .Y(n_589) );
AO21x1_ASAP7_75t_L g590 ( .A1(n_548), .A2(n_547), .B(n_546), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_549), .Y(n_591) );
INVxp67_ASAP7_75t_L g592 ( .A(n_531), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_510), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_526), .B(n_475), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_545), .A2(n_537), .B(n_536), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_526), .B(n_549), .Y(n_596) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_587), .B(n_583), .Y(n_597) );
AOI211xp5_ASAP7_75t_SL g598 ( .A1(n_595), .A2(n_586), .B(n_554), .C(n_569), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_576), .A2(n_559), .B(n_595), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_589), .A2(n_585), .B1(n_579), .B2(n_572), .Y(n_600) );
NAND3xp33_ASAP7_75t_SL g601 ( .A(n_562), .B(n_559), .C(n_590), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_588), .A2(n_591), .B(n_573), .C(n_557), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_576), .A2(n_585), .B(n_558), .Y(n_603) );
AOI321xp33_ASAP7_75t_L g604 ( .A1(n_594), .A2(n_558), .A3(n_578), .B1(n_560), .B2(n_551), .C(n_582), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_552), .A2(n_575), .B1(n_584), .B2(n_563), .Y(n_605) );
AOI211xp5_ASAP7_75t_SL g606 ( .A1(n_588), .A2(n_581), .B(n_592), .C(n_557), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_560), .B(n_571), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_573), .Y(n_608) );
INVx2_ASAP7_75t_SL g609 ( .A(n_607), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_599), .A2(n_592), .B(n_568), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_601), .A2(n_596), .B(n_556), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_597), .B(n_564), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_605), .B(n_564), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_598), .A2(n_566), .B(n_593), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_603), .A2(n_555), .B(n_570), .Y(n_615) );
OAI211xp5_ASAP7_75t_L g616 ( .A1(n_614), .A2(n_600), .B(n_604), .C(n_606), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_612), .A2(n_608), .B1(n_561), .B2(n_565), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_615), .A2(n_602), .B(n_567), .Y(n_618) );
OAI22xp33_ASAP7_75t_SL g619 ( .A1(n_610), .A2(n_553), .B1(n_574), .B2(n_577), .Y(n_619) );
XNOR2xp5_ASAP7_75t_L g620 ( .A(n_616), .B(n_611), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_617), .Y(n_621) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_620), .B(n_619), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_620), .Y(n_623) );
AND3x4_ASAP7_75t_L g624 ( .A(n_622), .B(n_621), .C(n_618), .Y(n_624) );
XNOR2xp5_ASAP7_75t_L g625 ( .A(n_624), .B(n_623), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_625), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_626), .A2(n_609), .B1(n_613), .B2(n_550), .C(n_580), .Y(n_627) );
endmodule