module fake_netlist_6_1142_n_1188 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1188);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1188;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_760;
wire n_680;
wire n_741;
wire n_465;
wire n_1027;
wire n_1008;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_1033;
wire n_1052;
wire n_671;
wire n_726;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_1164;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_955;
wire n_337;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1101;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_1139;
wire n_198;
wire n_300;
wire n_718;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_742;
wire n_532;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_1119;
wire n_344;
wire n_946;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_1163;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_838;
wire n_302;
wire n_499;
wire n_380;
wire n_294;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_1176;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_1181;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_236;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_1183;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_216;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_608;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_811;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_689;
wire n_354;
wire n_231;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_550;
wire n_487;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_1107;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_474;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_1167;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_1153;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_1185;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_1175;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1154;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1023;
wire n_1013;
wire n_1076;
wire n_1118;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_855;
wire n_283;

INVx1_ASAP7_75t_L g179 ( 
.A(n_12),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_68),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_103),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_88),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_55),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_70),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_108),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_42),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_126),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_91),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_25),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_10),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_95),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_54),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_43),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_129),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_45),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_63),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_111),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_76),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_44),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_115),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_52),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_20),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_151),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_69),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_0),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_2),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_3),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_166),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_64),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_177),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_4),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_82),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_4),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_49),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_137),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_77),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_11),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_48),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_20),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_207),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_182),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_184),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_185),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_189),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_190),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_192),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_208),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_195),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_196),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_198),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_199),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_204),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_205),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_206),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_209),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_215),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_245),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_247),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_237),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_238),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_256),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_255),
.Y(n_283)
);

BUFx8_ASAP7_75t_SL g284 ( 
.A(n_257),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_194),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_260),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_244),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_248),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_262),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_263),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_264),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_251),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_237),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_239),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_245),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_239),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_245),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

BUFx2_ASAP7_75t_SL g315 ( 
.A(n_237),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_239),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_237),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_275),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_291),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_287),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_284),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_292),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_268),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_277),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_277),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_297),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_276),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_283),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_308),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_300),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_283),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_271),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_269),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_317),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_317),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_288),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_272),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_279),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_287),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_280),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_267),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_310),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_312),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_314),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_316),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_270),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_289),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_307),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_276),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_224),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_319),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_224),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_304),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_325),
.B(n_352),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_327),
.B(n_333),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_285),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

CKINVDCx11_ASAP7_75t_R g377 ( 
.A(n_348),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_304),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_324),
.B(n_302),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_362),
.Y(n_380)
);

BUFx12f_ASAP7_75t_L g381 ( 
.A(n_332),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_282),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_337),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_342),
.B(n_350),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

BUFx12f_ASAP7_75t_L g388 ( 
.A(n_332),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_351),
.Y(n_389)
);

BUFx12f_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_325),
.B(n_302),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_355),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_338),
.B(n_303),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_356),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_295),
.Y(n_396)
);

BUFx12f_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_329),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

BUFx8_ASAP7_75t_SL g402 ( 
.A(n_326),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_363),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_347),
.B(n_181),
.Y(n_405)
);

BUFx12f_ASAP7_75t_L g406 ( 
.A(n_349),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_334),
.B(n_183),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_365),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_352),
.B(n_311),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_371),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_313),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_390),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_303),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

AND2x2_ASAP7_75t_SL g417 ( 
.A(n_389),
.B(n_181),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_395),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_370),
.B(n_197),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_399),
.A2(n_331),
.B1(n_346),
.B2(n_340),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_390),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_389),
.A2(n_227),
.B1(n_223),
.B2(n_208),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_389),
.A2(n_227),
.B1(n_223),
.B2(n_288),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_369),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_293),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_371),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_293),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_387),
.B(n_180),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_395),
.B(n_320),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_387),
.B(n_233),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_400),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_397),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_403),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_385),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_394),
.B(n_202),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_393),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_393),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_402),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_397),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_375),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_397),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_400),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_398),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_370),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_400),
.B(n_210),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_400),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_407),
.B(n_321),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_406),
.B(n_326),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_404),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_389),
.B(n_186),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_400),
.B(n_193),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_401),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_382),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_382),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_382),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_380),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_407),
.B(n_329),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_379),
.B(n_372),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_367),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_409),
.B(n_298),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_366),
.B(n_331),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_373),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_401),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_401),
.Y(n_478)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_366),
.B(n_335),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_380),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_410),
.B(n_202),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_366),
.B(n_368),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_383),
.B(n_335),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_409),
.B(n_298),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_401),
.B(n_203),
.Y(n_488)
);

AND2x6_ASAP7_75t_L g489 ( 
.A(n_378),
.B(n_197),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_396),
.B(n_340),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_366),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_406),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_430),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_438),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_R g495 ( 
.A(n_425),
.B(n_318),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_447),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_447),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_442),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_458),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_412),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_412),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_428),
.B(n_391),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_428),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_450),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_443),
.B(n_381),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_459),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_476),
.B(n_374),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_450),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_420),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_492),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_462),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_416),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_418),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_414),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_492),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_416),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_418),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_418),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_415),
.B(n_381),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_443),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_431),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_473),
.B(n_405),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_448),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_445),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_446),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_411),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_452),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_411),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_436),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_422),
.Y(n_534)
);

OA21x2_ASAP7_75t_L g535 ( 
.A1(n_466),
.A2(n_408),
.B(n_200),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_421),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_453),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_421),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_467),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_454),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_468),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_R g543 ( 
.A(n_461),
.B(n_346),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_422),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_433),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_444),
.B(n_348),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_441),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_434),
.Y(n_548)
);

NOR2xp67_ASAP7_75t_L g549 ( 
.A(n_473),
.B(n_406),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_479),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_441),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_434),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_500),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_514),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_508),
.B(n_415),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_552),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_552),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_525),
.A2(n_456),
.B(n_464),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_500),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_493),
.B(n_417),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_501),
.B(n_449),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_496),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_501),
.Y(n_563)
);

AOI21x1_ASAP7_75t_L g564 ( 
.A1(n_535),
.A2(n_456),
.B(n_464),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_514),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_496),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_514),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_546),
.B(n_444),
.Y(n_568)
);

AND2x2_ASAP7_75t_SL g569 ( 
.A(n_535),
.B(n_417),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_513),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_SL g571 ( 
.A(n_543),
.B(n_472),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_514),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_550),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_527),
.B(n_413),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_549),
.B(n_423),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_540),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_497),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_513),
.B(n_449),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_533),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_514),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_528),
.B(n_429),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_517),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_517),
.B(n_455),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_534),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_510),
.B(n_426),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_503),
.B(n_486),
.Y(n_586)
);

INVxp67_ASAP7_75t_SL g587 ( 
.A(n_534),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_504),
.Y(n_588)
);

CKINVDCx6p67_ASAP7_75t_R g589 ( 
.A(n_550),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_523),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_524),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_534),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_524),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_568),
.A2(n_482),
.B1(n_490),
.B2(n_510),
.Y(n_594)
);

INVx6_ASAP7_75t_L g595 ( 
.A(n_562),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_589),
.Y(n_596)
);

INVx6_ASAP7_75t_L g597 ( 
.A(n_562),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_568),
.A2(n_482),
.B1(n_405),
.B2(n_471),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_586),
.B(n_437),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_571),
.B(n_555),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_553),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_575),
.A2(n_405),
.B1(n_480),
.B2(n_475),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_554),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_573),
.B(n_479),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_559),
.Y(n_606)
);

AND2x6_ASAP7_75t_L g607 ( 
.A(n_565),
.B(n_534),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_554),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_588),
.B(n_437),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_589),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_559),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_574),
.B(n_506),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_574),
.B(n_460),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_573),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_589),
.Y(n_615)
);

INVx6_ASAP7_75t_L g616 ( 
.A(n_562),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_573),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_563),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_581),
.B(n_435),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_563),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_588),
.A2(n_388),
.B1(n_495),
.B2(n_479),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_579),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_554),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_585),
.A2(n_405),
.B1(n_480),
.B2(n_475),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_565),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_585),
.B(n_377),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_590),
.B(n_435),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_579),
.B(n_483),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_556),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_576),
.B(n_388),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_576),
.B(n_530),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_590),
.B(n_537),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_561),
.B(n_439),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_562),
.Y(n_634)
);

BUFx4f_ASAP7_75t_L g635 ( 
.A(n_565),
.Y(n_635)
);

AND2x6_ASAP7_75t_L g636 ( 
.A(n_565),
.B(n_534),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_554),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_566),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_577),
.B(n_388),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_577),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_577),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_577),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_561),
.B(n_439),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_565),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_567),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_557),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_567),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_560),
.B(n_526),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_560),
.B(n_526),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_561),
.B(n_483),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_565),
.B(n_542),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_558),
.A2(n_405),
.B1(n_419),
.B2(n_463),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_569),
.B(n_451),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_558),
.A2(n_405),
.B1(n_419),
.B2(n_463),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_557),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_578),
.B(n_519),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_565),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_580),
.B(n_521),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_570),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_578),
.B(n_522),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_569),
.B(n_451),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_584),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_578),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_570),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_570),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_582),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_583),
.B(n_432),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_582),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_584),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_572),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_572),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_599),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_594),
.A2(n_419),
.B(n_463),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_606),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_620),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_638),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_605),
.B(n_595),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_642),
.B(n_572),
.Y(n_678)
);

BUFx6f_ASAP7_75t_SL g679 ( 
.A(n_638),
.Y(n_679)
);

XOR2x2_ASAP7_75t_L g680 ( 
.A(n_626),
.B(n_515),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_602),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_611),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_618),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_646),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_613),
.B(n_667),
.Y(n_685)
);

BUFx2_ASAP7_75t_R g686 ( 
.A(n_630),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_646),
.Y(n_687)
);

INVxp33_ASAP7_75t_L g688 ( 
.A(n_627),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_655),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_612),
.B(n_464),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_655),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_666),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_619),
.B(n_591),
.Y(n_693)
);

AND2x6_ASAP7_75t_L g694 ( 
.A(n_604),
.B(n_584),
.Y(n_694)
);

AND2x6_ASAP7_75t_L g695 ( 
.A(n_604),
.B(n_584),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_668),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_668),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_634),
.B(n_572),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_601),
.A2(n_569),
.B(n_587),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_614),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_664),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_629),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_641),
.B(n_592),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_632),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_639),
.B(n_531),
.Y(n_705)
);

AND2x2_ASAP7_75t_SL g706 ( 
.A(n_596),
.B(n_485),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_SL g707 ( 
.A(n_596),
.B(n_497),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_622),
.B(n_591),
.Y(n_708)
);

INVxp33_ASAP7_75t_L g709 ( 
.A(n_628),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_610),
.B(n_505),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_659),
.Y(n_711)
);

XOR2x2_ASAP7_75t_SL g712 ( 
.A(n_631),
.B(n_191),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_665),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_647),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_609),
.Y(n_715)
);

XOR2xp5_ASAP7_75t_L g716 ( 
.A(n_600),
.B(n_515),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_656),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_628),
.B(n_505),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_650),
.B(n_488),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_660),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_663),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_645),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_645),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_614),
.B(n_488),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_R g725 ( 
.A(n_605),
.B(n_509),
.Y(n_725)
);

INVx4_ASAP7_75t_SL g726 ( 
.A(n_595),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_621),
.B(n_509),
.Y(n_727)
);

AND2x2_ASAP7_75t_SL g728 ( 
.A(n_610),
.B(n_584),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_614),
.B(n_488),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_670),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_648),
.B(n_511),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_670),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_649),
.Y(n_733)
);

XOR2xp5_ASAP7_75t_L g734 ( 
.A(n_624),
.B(n_511),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_633),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_643),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_640),
.B(n_516),
.Y(n_737)
);

INVx4_ASAP7_75t_SL g738 ( 
.A(n_597),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_617),
.B(n_516),
.Y(n_739)
);

NOR2xp67_ASAP7_75t_L g740 ( 
.A(n_615),
.B(n_531),
.Y(n_740)
);

INVxp33_ASAP7_75t_L g741 ( 
.A(n_617),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_597),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_671),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_616),
.Y(n_744)
);

XNOR2xp5_ASAP7_75t_L g745 ( 
.A(n_603),
.B(n_529),
.Y(n_745)
);

AOI21x1_ASAP7_75t_L g746 ( 
.A1(n_653),
.A2(n_564),
.B(n_661),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_615),
.B(n_542),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_704),
.B(n_558),
.Y(n_748)
);

AND2x2_ASAP7_75t_SL g749 ( 
.A(n_706),
.B(n_635),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_736),
.B(n_558),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_737),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_717),
.B(n_598),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_712),
.B(n_617),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_720),
.B(n_616),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_681),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_682),
.B(n_608),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_705),
.B(n_740),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_733),
.A2(n_405),
.B1(n_419),
.B2(n_191),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_683),
.B(n_608),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_715),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_672),
.B(n_623),
.Y(n_761)
);

AOI22x1_ASAP7_75t_L g762 ( 
.A1(n_734),
.A2(n_536),
.B1(n_547),
.B2(n_538),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_L g763 ( 
.A(n_742),
.B(n_536),
.Y(n_763)
);

INVx5_ASAP7_75t_L g764 ( 
.A(n_694),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_672),
.Y(n_765)
);

AND2x6_ASAP7_75t_L g766 ( 
.A(n_690),
.B(n_735),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_714),
.B(n_726),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_710),
.B(n_635),
.Y(n_768)
);

INVx8_ASAP7_75t_L g769 ( 
.A(n_677),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_744),
.B(n_538),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_685),
.B(n_658),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_721),
.B(n_658),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_707),
.B(n_625),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_688),
.B(n_662),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_727),
.B(n_625),
.Y(n_775)
);

BUFx8_ASAP7_75t_L g776 ( 
.A(n_679),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_716),
.B(n_529),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_731),
.B(n_726),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_674),
.B(n_637),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_738),
.B(n_625),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_709),
.B(n_547),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_711),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_718),
.B(n_551),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_700),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_739),
.B(n_551),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_738),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_693),
.B(n_637),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_673),
.A2(n_654),
.B(n_652),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_675),
.B(n_591),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_713),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_684),
.B(n_593),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_687),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_702),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_676),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_689),
.B(n_593),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_691),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_728),
.B(n_644),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_678),
.B(n_644),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_701),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_692),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_677),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_708),
.B(n_662),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_743),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_719),
.A2(n_419),
.B1(n_489),
.B2(n_200),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_678),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_SL g806 ( 
.A(n_686),
.B(n_657),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_696),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_697),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_722),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_725),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_699),
.B(n_593),
.Y(n_811)
);

NAND2x1_ASAP7_75t_L g812 ( 
.A(n_694),
.B(n_695),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_723),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_765),
.Y(n_814)
);

OAI221xp5_ASAP7_75t_L g815 ( 
.A1(n_753),
.A2(n_745),
.B1(n_219),
.B2(n_236),
.C(n_220),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_805),
.B(n_698),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_750),
.B(n_730),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_749),
.B(n_698),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_760),
.B(n_732),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_803),
.B(n_703),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_755),
.Y(n_821)
);

NAND2x1p5_ASAP7_75t_L g822 ( 
.A(n_764),
.B(n_644),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_792),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_796),
.Y(n_824)
);

NAND2x1p5_ASAP7_75t_L g825 ( 
.A(n_764),
.B(n_703),
.Y(n_825)
);

OAI221xp5_ASAP7_75t_L g826 ( 
.A1(n_810),
.A2(n_236),
.B1(n_680),
.B2(n_222),
.C(n_217),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_784),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_787),
.B(n_746),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_800),
.Y(n_829)
);

AO22x2_ASAP7_75t_L g830 ( 
.A1(n_750),
.A2(n_729),
.B1(n_724),
.B2(n_669),
.Y(n_830)
);

AO22x2_ASAP7_75t_L g831 ( 
.A1(n_748),
.A2(n_669),
.B1(n_580),
.B2(n_587),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_807),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_808),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_776),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_774),
.B(n_741),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_805),
.B(n_747),
.Y(n_836)
);

AO22x2_ASAP7_75t_L g837 ( 
.A1(n_748),
.A2(n_580),
.B1(n_592),
.B2(n_498),
.Y(n_837)
);

OAI221xp5_ASAP7_75t_L g838 ( 
.A1(n_751),
.A2(n_234),
.B1(n_229),
.B2(n_218),
.C(n_216),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_788),
.A2(n_679),
.B1(n_489),
.B2(n_211),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_767),
.B(n_694),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_771),
.B(n_694),
.Y(n_841)
);

NAND2x1p5_ASAP7_75t_L g842 ( 
.A(n_764),
.B(n_584),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_764),
.B(n_695),
.Y(n_843)
);

AO22x2_ASAP7_75t_L g844 ( 
.A1(n_799),
.A2(n_592),
.B1(n_499),
.B2(n_507),
.Y(n_844)
);

NAND2x1p5_ASAP7_75t_L g845 ( 
.A(n_773),
.B(n_584),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_782),
.B(n_695),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_790),
.B(n_695),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_809),
.Y(n_848)
);

AO22x2_ASAP7_75t_L g849 ( 
.A1(n_813),
.A2(n_592),
.B1(n_512),
.B2(n_494),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_801),
.B(n_778),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_780),
.B(n_542),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_788),
.A2(n_188),
.B(n_232),
.C(n_187),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_761),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_761),
.Y(n_854)
);

INVxp33_ASAP7_75t_SL g855 ( 
.A(n_777),
.Y(n_855)
);

AO22x2_ASAP7_75t_L g856 ( 
.A1(n_754),
.A2(n_541),
.B1(n_539),
.B2(n_532),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_756),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_759),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_762),
.A2(n_491),
.B1(n_548),
.B2(n_545),
.Y(n_859)
);

NAND2x1p5_ASAP7_75t_L g860 ( 
.A(n_786),
.B(n_542),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_754),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_775),
.A2(n_489),
.B1(n_429),
.B2(n_432),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_766),
.A2(n_489),
.B1(n_429),
.B2(n_368),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_776),
.Y(n_864)
);

AO22x2_ASAP7_75t_L g865 ( 
.A1(n_772),
.A2(n_502),
.B1(n_532),
.B2(n_544),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_767),
.B(n_607),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_779),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_793),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_811),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_785),
.B(n_794),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_789),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_789),
.Y(n_872)
);

BUFx8_ASAP7_75t_L g873 ( 
.A(n_784),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_811),
.Y(n_874)
);

NOR2xp67_ASAP7_75t_L g875 ( 
.A(n_786),
.B(n_0),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_784),
.Y(n_876)
);

NAND2x1p5_ASAP7_75t_L g877 ( 
.A(n_797),
.B(n_542),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_791),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_791),
.Y(n_879)
);

AO22x2_ASAP7_75t_L g880 ( 
.A1(n_812),
.A2(n_502),
.B1(n_532),
.B2(n_544),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_795),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_814),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_839),
.A2(n_768),
.B(n_757),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_841),
.B(n_766),
.Y(n_884)
);

CKINVDCx8_ASAP7_75t_R g885 ( 
.A(n_864),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_852),
.A2(n_798),
.B(n_806),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_831),
.A2(n_752),
.B(n_769),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_861),
.B(n_769),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_855),
.B(n_769),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_840),
.B(n_781),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_869),
.A2(n_752),
.B(n_763),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_857),
.B(n_802),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_838),
.A2(n_783),
.B(n_770),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_818),
.A2(n_758),
.B(n_804),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_850),
.B(n_766),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_843),
.B(n_766),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_SL g897 ( 
.A(n_834),
.B(n_607),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_828),
.A2(n_535),
.B(n_477),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_823),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_874),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_815),
.A2(n_187),
.B(n_188),
.C(n_232),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_842),
.A2(n_544),
.B(n_502),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_876),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_856),
.A2(n_487),
.B(n_474),
.Y(n_904)
);

AOI33xp33_ASAP7_75t_L g905 ( 
.A1(n_858),
.A2(n_368),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.B3(n_6),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_873),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_870),
.B(n_1),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_826),
.A2(n_368),
.B(n_607),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_853),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_843),
.B(n_211),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_865),
.A2(n_440),
.B(n_469),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_SL g912 ( 
.A1(n_819),
.A2(n_1),
.B(n_5),
.C(n_6),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_867),
.B(n_636),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_L g914 ( 
.A(n_825),
.B(n_211),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_831),
.A2(n_440),
.B(n_451),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_865),
.A2(n_470),
.B(n_469),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_875),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_837),
.A2(n_481),
.B(n_470),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_854),
.B(n_636),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_830),
.B(n_636),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_837),
.A2(n_484),
.B(n_481),
.Y(n_921)
);

AO21x1_ASAP7_75t_L g922 ( 
.A1(n_824),
.A2(n_7),
.B(n_8),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_844),
.A2(n_457),
.B(n_451),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_844),
.A2(n_465),
.B(n_457),
.Y(n_924)
);

NOR2x1p5_ASAP7_75t_L g925 ( 
.A(n_820),
.B(n_211),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_829),
.Y(n_926)
);

AO21x1_ASAP7_75t_L g927 ( 
.A1(n_832),
.A2(n_9),
.B(n_10),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_827),
.Y(n_928)
);

NOR3xp33_ASAP7_75t_SL g929 ( 
.A(n_893),
.B(n_847),
.C(n_846),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_900),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_884),
.B(n_830),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_909),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_SL g933 ( 
.A(n_901),
.B(n_213),
.C(n_212),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_891),
.B(n_892),
.Y(n_934)
);

HAxp5_ASAP7_75t_L g935 ( 
.A(n_925),
.B(n_11),
.CON(n_935),
.SN(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_906),
.Y(n_936)
);

BUFx4f_ASAP7_75t_L g937 ( 
.A(n_885),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_903),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_887),
.B(n_821),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_887),
.B(n_816),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_882),
.Y(n_941)
);

INVx6_ASAP7_75t_L g942 ( 
.A(n_903),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_899),
.Y(n_943)
);

INVx5_ASAP7_75t_L g944 ( 
.A(n_920),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_922),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_926),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_896),
.B(n_836),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_919),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_928),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_889),
.B(n_866),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_913),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_R g952 ( 
.A(n_914),
.B(n_12),
.Y(n_952)
);

AO21x1_ASAP7_75t_L g953 ( 
.A1(n_907),
.A2(n_833),
.B(n_851),
.Y(n_953)
);

AOI211xp5_ASAP7_75t_L g954 ( 
.A1(n_927),
.A2(n_817),
.B(n_835),
.C(n_848),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_888),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_890),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_895),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_902),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_910),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_915),
.B(n_871),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_923),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_897),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_915),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_912),
.B(n_872),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_883),
.B(n_863),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_883),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_SL g967 ( 
.A(n_905),
.B(n_878),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_923),
.Y(n_968)
);

CKINVDCx11_ASAP7_75t_R g969 ( 
.A(n_917),
.Y(n_969)
);

NOR2xp67_ASAP7_75t_L g970 ( 
.A(n_924),
.B(n_879),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_924),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_908),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_886),
.B(n_881),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_916),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_918),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_921),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_886),
.Y(n_977)
);

NOR3xp33_ASAP7_75t_SL g978 ( 
.A(n_894),
.B(n_225),
.C(n_214),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_911),
.Y(n_979)
);

BUFx4f_ASAP7_75t_L g980 ( 
.A(n_904),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_898),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_907),
.B(n_868),
.Y(n_982)
);

AND3x1_ASAP7_75t_SL g983 ( 
.A(n_925),
.B(n_13),
.C(n_14),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_906),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_977),
.A2(n_862),
.B1(n_880),
.B2(n_849),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_945),
.A2(n_880),
.B(n_849),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_943),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_943),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_973),
.B(n_877),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_937),
.B(n_845),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_941),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_973),
.B(n_860),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_984),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_934),
.B(n_822),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_942),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_954),
.B(n_859),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_929),
.B(n_14),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_966),
.B(n_211),
.Y(n_998)
);

BUFx12f_ASAP7_75t_L g999 ( 
.A(n_936),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_937),
.B(n_15),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_969),
.B(n_15),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_945),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_980),
.A2(n_230),
.B1(n_231),
.B2(n_520),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_938),
.A2(n_940),
.B(n_963),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_1004),
.A2(n_940),
.B(n_939),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_993),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_999),
.B(n_956),
.Y(n_1007)
);

INVx8_ASAP7_75t_L g1008 ( 
.A(n_993),
.Y(n_1008)
);

BUFx4f_ASAP7_75t_L g1009 ( 
.A(n_993),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_995),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_995),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_996),
.A2(n_972),
.B1(n_980),
.B2(n_965),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_994),
.B(n_931),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_987),
.Y(n_1014)
);

CKINVDCx6p67_ASAP7_75t_R g1015 ( 
.A(n_997),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_991),
.B(n_964),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_985),
.A2(n_942),
.B1(n_957),
.B2(n_944),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_988),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_1001),
.A2(n_942),
.B1(n_944),
.B2(n_949),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_1000),
.B(n_950),
.Y(n_1020)
);

AOI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_1002),
.A2(n_981),
.B(n_976),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_990),
.B(n_949),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_989),
.A2(n_944),
.B1(n_929),
.B2(n_964),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_998),
.B(n_962),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_986),
.A2(n_935),
.B(n_953),
.C(n_963),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_992),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1003),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_1001),
.A2(n_967),
.B(n_978),
.C(n_933),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_991),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_1025),
.B(n_944),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_SL g1031 ( 
.A(n_1006),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1015),
.B(n_982),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_1005),
.A2(n_978),
.B(n_933),
.C(n_979),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1011),
.B(n_982),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1018),
.Y(n_1035)
);

AO31x2_ASAP7_75t_L g1036 ( 
.A1(n_1019),
.A2(n_932),
.A3(n_961),
.B(n_971),
.Y(n_1036)
);

AO21x2_ASAP7_75t_L g1037 ( 
.A1(n_1030),
.A2(n_1023),
.B(n_1017),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1035),
.B(n_1006),
.Y(n_1038)
);

AO21x1_ASAP7_75t_L g1039 ( 
.A1(n_1038),
.A2(n_1010),
.B(n_1014),
.Y(n_1039)
);

BUFx8_ASAP7_75t_L g1040 ( 
.A(n_1037),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1040),
.A2(n_1033),
.B(n_1028),
.Y(n_1041)
);

CKINVDCx6p67_ASAP7_75t_R g1042 ( 
.A(n_1039),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1042),
.A2(n_1031),
.B1(n_1012),
.B2(n_1009),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_SL g1044 ( 
.A1(n_1041),
.A2(n_1006),
.B1(n_1032),
.B2(n_1027),
.Y(n_1044)
);

AO31x2_ASAP7_75t_L g1045 ( 
.A1(n_1042),
.A2(n_1010),
.A3(n_1007),
.B(n_1014),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_1045),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1044),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1043),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1046),
.Y(n_1049)
);

NOR2x1p5_ASAP7_75t_L g1050 ( 
.A(n_1047),
.B(n_1034),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1050),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_1049),
.B(n_1047),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1051),
.B(n_1048),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1052),
.B(n_1008),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1053),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1054),
.B(n_1008),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_SL g1057 ( 
.A1(n_1055),
.A2(n_1022),
.B(n_1020),
.Y(n_1057)
);

OAI21xp33_ASAP7_75t_L g1058 ( 
.A1(n_1056),
.A2(n_1016),
.B(n_1026),
.Y(n_1058)
);

AOI33xp33_ASAP7_75t_L g1059 ( 
.A1(n_1057),
.A2(n_1029),
.A3(n_1013),
.B1(n_1036),
.B2(n_955),
.B3(n_959),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_1058),
.B(n_1036),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1060),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_1059),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1059),
.B(n_1021),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_1063),
.B(n_1061),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1062),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1063),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1065),
.B(n_930),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_1064),
.B(n_930),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_1067),
.B(n_1066),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1068),
.B(n_1024),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1070),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1069),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1072),
.B(n_16),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1071),
.B(n_17),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_1074),
.B(n_294),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1073),
.B(n_951),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_1075),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_1076),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1078),
.A2(n_408),
.B(n_18),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1077),
.A2(n_968),
.B1(n_951),
.B2(n_979),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1078),
.B(n_19),
.Y(n_1081)
);

O2A1O1Ixp5_ASAP7_75t_L g1082 ( 
.A1(n_1079),
.A2(n_1081),
.B(n_1080),
.C(n_408),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_1081),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1081),
.Y(n_1084)
);

OAI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_1083),
.A2(n_1082),
.B1(n_1084),
.B2(n_22),
.C(n_23),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1083),
.A2(n_968),
.B1(n_21),
.B2(n_22),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1085),
.B(n_19),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_1086),
.B(n_294),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1087),
.B(n_948),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1088),
.A2(n_294),
.B1(n_23),
.B2(n_24),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1089),
.B(n_21),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_1090),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1092),
.A2(n_294),
.B1(n_25),
.B2(n_26),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_L g1094 ( 
.A1(n_1091),
.A2(n_408),
.B1(n_276),
.B2(n_27),
.C(n_28),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_1094),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1093),
.A2(n_270),
.B(n_26),
.C(n_27),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_1095),
.Y(n_1097)
);

AOI221xp5_ASAP7_75t_L g1098 ( 
.A1(n_1096),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_1098)
);

XOR2x2_ASAP7_75t_L g1099 ( 
.A(n_1095),
.B(n_29),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_SL g1100 ( 
.A(n_1097),
.B(n_952),
.C(n_30),
.Y(n_1100)
);

NAND4xp25_ASAP7_75t_L g1101 ( 
.A(n_1098),
.B(n_1099),
.C(n_31),
.D(n_33),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1099),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_1102),
.Y(n_1103)
);

OAI222xp33_ASAP7_75t_L g1104 ( 
.A1(n_1101),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.C1(n_35),
.C2(n_36),
.Y(n_1104)
);

NOR2x1p5_ASAP7_75t_L g1105 ( 
.A(n_1103),
.B(n_1100),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_L g1106 ( 
.A(n_1104),
.B(n_298),
.C(n_37),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1105),
.B(n_1106),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_1105),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1108),
.B(n_38),
.Y(n_1109)
);

AOI221xp5_ASAP7_75t_L g1110 ( 
.A1(n_1107),
.A2(n_952),
.B1(n_40),
.B2(n_41),
.C(n_46),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_1109),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1110),
.B(n_39),
.Y(n_1112)
);

AND4x1_ASAP7_75t_L g1113 ( 
.A(n_1112),
.B(n_47),
.C(n_50),
.D(n_51),
.Y(n_1113)
);

XNOR2x1_ASAP7_75t_L g1114 ( 
.A(n_1111),
.B(n_53),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_R g1115 ( 
.A(n_1113),
.B(n_56),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_1114),
.B(n_57),
.Y(n_1116)
);

NAND2xp33_ASAP7_75t_SL g1117 ( 
.A(n_1114),
.B(n_58),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1115),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1117),
.B(n_59),
.Y(n_1119)
);

AND3x4_ASAP7_75t_L g1120 ( 
.A(n_1116),
.B(n_60),
.C(n_61),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1118),
.Y(n_1121)
);

OAI22x1_ASAP7_75t_L g1122 ( 
.A1(n_1119),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1121),
.B(n_1120),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1122),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1123),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_SL g1126 ( 
.A1(n_1124),
.A2(n_67),
.B1(n_71),
.B2(n_72),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1125),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1126),
.A2(n_983),
.B1(n_74),
.B2(n_75),
.Y(n_1128)
);

XNOR2xp5_ASAP7_75t_L g1129 ( 
.A(n_1127),
.B(n_73),
.Y(n_1129)
);

AOI31xp33_ASAP7_75t_L g1130 ( 
.A1(n_1128),
.A2(n_78),
.A3(n_79),
.B(n_80),
.Y(n_1130)
);

AO21x2_ASAP7_75t_L g1131 ( 
.A1(n_1130),
.A2(n_81),
.B(n_83),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1129),
.A2(n_84),
.B(n_86),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1131),
.Y(n_1133)
);

XNOR2xp5_ASAP7_75t_L g1134 ( 
.A(n_1132),
.B(n_87),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1131),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1133),
.Y(n_1136)
);

NOR2x1p5_ASAP7_75t_L g1137 ( 
.A(n_1135),
.B(n_1134),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1133),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1136),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_1138),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1139),
.B(n_1137),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1140),
.B(n_89),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1141),
.A2(n_983),
.B1(n_520),
.B2(n_518),
.Y(n_1143)
);

OAI322xp33_ASAP7_75t_L g1144 ( 
.A1(n_1142),
.A2(n_90),
.A3(n_92),
.B1(n_93),
.B2(n_94),
.C1(n_96),
.C2(n_97),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1144),
.Y(n_1145)
);

XOR2xp5_ASAP7_75t_L g1146 ( 
.A(n_1143),
.B(n_98),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1144),
.A2(n_99),
.B(n_100),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1145),
.A2(n_520),
.B1(n_518),
.B2(n_651),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1146),
.A2(n_520),
.B1(n_518),
.B2(n_651),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1147),
.A2(n_518),
.B1(n_651),
.B2(n_104),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1150),
.A2(n_101),
.B(n_102),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1149),
.A2(n_105),
.B(n_106),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1148),
.A2(n_107),
.B(n_109),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1151),
.A2(n_110),
.B(n_113),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1152),
.B(n_114),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1153),
.Y(n_1156)
);

NAND2x1p5_ASAP7_75t_L g1157 ( 
.A(n_1151),
.B(n_116),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1151),
.A2(n_117),
.B(n_120),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_L g1159 ( 
.A(n_1151),
.B(n_121),
.C(n_122),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1151),
.B(n_123),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_1151),
.B(n_124),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1151),
.A2(n_125),
.B(n_127),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1151),
.A2(n_128),
.B(n_130),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1151),
.B(n_131),
.Y(n_1164)
);

AOI21xp33_ASAP7_75t_SL g1165 ( 
.A1(n_1151),
.A2(n_132),
.B(n_133),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1151),
.B(n_134),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1156),
.A2(n_1161),
.B1(n_1157),
.B2(n_1164),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1160),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1166),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1155),
.A2(n_135),
.B1(n_139),
.B2(n_140),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1154),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1158),
.A2(n_1162),
.B1(n_1163),
.B2(n_1165),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1159),
.A2(n_651),
.B1(n_143),
.B2(n_144),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1156),
.Y(n_1174)
);

AOI322xp5_ASAP7_75t_L g1175 ( 
.A1(n_1156),
.A2(n_142),
.A3(n_145),
.B1(n_146),
.B2(n_147),
.C1(n_148),
.C2(n_149),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1174),
.A2(n_150),
.B(n_153),
.Y(n_1176)
);

AO221x2_ASAP7_75t_L g1177 ( 
.A1(n_1171),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.C(n_158),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1167),
.A2(n_159),
.B(n_161),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1168),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1169),
.A2(n_168),
.B(n_169),
.Y(n_1180)
);

AO221x2_ASAP7_75t_L g1181 ( 
.A1(n_1172),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.C(n_176),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_L g1182 ( 
.A1(n_1180),
.A2(n_1173),
.B1(n_1170),
.B2(n_1175),
.C(n_478),
.Y(n_1182)
);

AOI221xp5_ASAP7_75t_L g1183 ( 
.A1(n_1178),
.A2(n_478),
.B1(n_465),
.B2(n_457),
.C(n_958),
.Y(n_1183)
);

AOI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1176),
.A2(n_478),
.B1(n_465),
.B2(n_457),
.C(n_380),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1182),
.A2(n_1177),
.B1(n_1181),
.B2(n_1179),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1185),
.A2(n_1184),
.B1(n_1183),
.B2(n_947),
.Y(n_1186)
);

AOI211xp5_ASAP7_75t_L g1187 ( 
.A1(n_1186),
.A2(n_947),
.B(n_970),
.C(n_946),
.Y(n_1187)
);

AOI211xp5_ASAP7_75t_L g1188 ( 
.A1(n_1187),
.A2(n_975),
.B(n_960),
.C(n_974),
.Y(n_1188)
);


endmodule