module fake_aes_4303_n_149 (n_45, n_20, n_2, n_38, n_44, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_49, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_12, n_9, n_17, n_14, n_10, n_15, n_42, n_24, n_19, n_21, n_6, n_4, n_29, n_43, n_7, n_40, n_27, n_39, n_149);
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_49;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_149;
wire n_117;
wire n_133;
wire n_81;
wire n_69;
wire n_57;
wire n_88;
wire n_52;
wire n_102;
wire n_73;
wire n_119;
wire n_141;
wire n_115;
wire n_97;
wire n_80;
wire n_107;
wire n_60;
wire n_114;
wire n_121;
wire n_94;
wire n_65;
wire n_125;
wire n_130;
wire n_103;
wire n_87;
wire n_137;
wire n_104;
wire n_98;
wire n_74;
wire n_146;
wire n_85;
wire n_101;
wire n_62;
wire n_91;
wire n_108;
wire n_116;
wire n_139;
wire n_113;
wire n_95;
wire n_124;
wire n_128;
wire n_120;
wire n_129;
wire n_70;
wire n_90;
wire n_71;
wire n_63;
wire n_56;
wire n_135;
wire n_78;
wire n_127;
wire n_111;
wire n_79;
wire n_64;
wire n_142;
wire n_58;
wire n_122;
wire n_138;
wire n_126;
wire n_118;
wire n_84;
wire n_131;
wire n_112;
wire n_55;
wire n_86;
wire n_143;
wire n_75;
wire n_105;
wire n_72;
wire n_136;
wire n_76;
wire n_89;
wire n_68;
wire n_144;
wire n_53;
wire n_77;
wire n_67;
wire n_147;
wire n_54;
wire n_148;
wire n_123;
wire n_83;
wire n_100;
wire n_92;
wire n_59;
wire n_110;
wire n_66;
wire n_134;
wire n_82;
wire n_106;
wire n_145;
wire n_61;
wire n_99;
wire n_109;
wire n_93;
wire n_132;
wire n_51;
wire n_140;
wire n_96;
CKINVDCx5p33_ASAP7_75t_R g51 ( .A(n_45), .Y(n_51) );
INVx1_ASAP7_75t_L g52 ( .A(n_48), .Y(n_52) );
INVx1_ASAP7_75t_L g53 ( .A(n_8), .Y(n_53) );
INVx1_ASAP7_75t_L g54 ( .A(n_31), .Y(n_54) );
INVx1_ASAP7_75t_L g55 ( .A(n_24), .Y(n_55) );
CKINVDCx5p33_ASAP7_75t_R g56 ( .A(n_25), .Y(n_56) );
INVx2_ASAP7_75t_SL g57 ( .A(n_49), .Y(n_57) );
INVx1_ASAP7_75t_L g58 ( .A(n_18), .Y(n_58) );
CKINVDCx5p33_ASAP7_75t_R g59 ( .A(n_6), .Y(n_59) );
CKINVDCx5p33_ASAP7_75t_R g60 ( .A(n_44), .Y(n_60) );
INVx3_ASAP7_75t_L g61 ( .A(n_23), .Y(n_61) );
CKINVDCx5p33_ASAP7_75t_R g62 ( .A(n_20), .Y(n_62) );
INVx1_ASAP7_75t_L g63 ( .A(n_13), .Y(n_63) );
INVx3_ASAP7_75t_L g64 ( .A(n_47), .Y(n_64) );
INVx2_ASAP7_75t_L g65 ( .A(n_11), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_7), .Y(n_66) );
INVx2_ASAP7_75t_L g67 ( .A(n_42), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_21), .Y(n_68) );
OR2x2_ASAP7_75t_L g69 ( .A(n_46), .B(n_9), .Y(n_69) );
CKINVDCx5p33_ASAP7_75t_R g70 ( .A(n_36), .Y(n_70) );
INVx2_ASAP7_75t_SL g71 ( .A(n_22), .Y(n_71) );
HB1xp67_ASAP7_75t_L g72 ( .A(n_5), .Y(n_72) );
CKINVDCx5p33_ASAP7_75t_R g73 ( .A(n_43), .Y(n_73) );
INVx2_ASAP7_75t_SL g74 ( .A(n_26), .Y(n_74) );
HB1xp67_ASAP7_75t_L g75 ( .A(n_3), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_1), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_4), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_34), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_41), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_0), .Y(n_80) );
BUFx6f_ASAP7_75t_L g81 ( .A(n_61), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_75), .B(n_0), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_72), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_64), .Y(n_84) );
OA21x2_ASAP7_75t_L g85 ( .A1(n_52), .A2(n_27), .B(n_50), .Y(n_85) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_57), .B(n_2), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_76), .Y(n_87) );
AND2x4_ASAP7_75t_L g88 ( .A(n_77), .B(n_2), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_53), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_80), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g91 ( .A(n_89), .B(n_71), .Y(n_91) );
NOR2xp33_ASAP7_75t_L g92 ( .A(n_83), .B(n_74), .Y(n_92) );
HB1xp67_ASAP7_75t_L g93 ( .A(n_82), .Y(n_93) );
AOI21x1_ASAP7_75t_L g94 ( .A1(n_85), .A2(n_55), .B(n_54), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_81), .Y(n_95) );
AND2x4_ASAP7_75t_L g96 ( .A(n_84), .B(n_58), .Y(n_96) );
INVx3_ASAP7_75t_L g97 ( .A(n_88), .Y(n_97) );
AOI22xp33_ASAP7_75t_L g98 ( .A1(n_93), .A2(n_89), .B1(n_90), .B2(n_87), .Y(n_98) );
BUFx8_ASAP7_75t_L g99 ( .A(n_96), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g100 ( .A(n_97), .B(n_86), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_95), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_94), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_100), .A2(n_91), .B(n_92), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g104 ( .A(n_98), .B(n_51), .Y(n_104) );
INVx5_ASAP7_75t_L g105 ( .A(n_102), .Y(n_105) );
BUFx12f_ASAP7_75t_L g106 ( .A(n_99), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_101), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g108 ( .A1(n_103), .A2(n_102), .B(n_69), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_107), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_106), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g111 ( .A1(n_105), .A2(n_102), .B(n_63), .Y(n_111) );
AOI21x1_ASAP7_75t_L g112 ( .A1(n_104), .A2(n_68), .B(n_66), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_109), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_110), .Y(n_114) );
AOI21x1_ASAP7_75t_L g115 ( .A1(n_112), .A2(n_79), .B(n_78), .Y(n_115) );
OAI21x1_ASAP7_75t_L g116 ( .A1(n_111), .A2(n_67), .B(n_65), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_108), .A2(n_59), .B(n_56), .Y(n_117) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_108), .A2(n_62), .B(n_60), .Y(n_118) );
BUFx10_ASAP7_75t_L g119 ( .A(n_114), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_113), .Y(n_120) );
AOI21x1_ASAP7_75t_L g121 ( .A1(n_115), .A2(n_73), .B(n_70), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_118), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_116), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_117), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_113), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_113), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_120), .B(n_10), .Y(n_127) );
AO31x2_ASAP7_75t_L g128 ( .A1(n_123), .A2(n_12), .A3(n_14), .B(n_15), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_125), .B(n_16), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_126), .B(n_17), .Y(n_130) );
INVx11_ASAP7_75t_L g131 ( .A(n_119), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_124), .B(n_19), .Y(n_132) );
INVx5_ASAP7_75t_L g133 ( .A(n_122), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_133), .Y(n_134) );
AND2x6_ASAP7_75t_SL g135 ( .A(n_131), .B(n_121), .Y(n_135) );
INVx1_ASAP7_75t_SL g136 ( .A(n_134), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_136), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_137), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_138), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_139), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_140), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_141), .Y(n_142) );
AO22x2_ASAP7_75t_L g143 ( .A1(n_142), .A2(n_135), .B1(n_132), .B2(n_130), .Y(n_143) );
AOI211x1_ASAP7_75t_L g144 ( .A1(n_143), .A2(n_135), .B(n_129), .C(n_127), .Y(n_144) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_144), .A2(n_128), .B1(n_28), .B2(n_29), .Y(n_145) );
AND3x1_ASAP7_75t_L g146 ( .A(n_145), .B(n_128), .C(n_30), .Y(n_146) );
AO21x2_ASAP7_75t_L g147 ( .A1(n_146), .A2(n_32), .B(n_33), .Y(n_147) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_147), .A2(n_35), .B(n_37), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_148), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_149) );
endmodule