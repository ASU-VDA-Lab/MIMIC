module fake_jpeg_24279_n_251 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_46),
.Y(n_50)
);

HAxp5_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_0),
.CON(n_39),
.SN(n_39)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_22),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_0),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_67),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_17),
.B1(n_35),
.B2(n_21),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_35),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_64),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_29),
.B1(n_30),
.B2(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_33),
.B1(n_26),
.B2(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_17),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_79),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_25),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_44),
.B1(n_30),
.B2(n_45),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_99),
.B1(n_18),
.B2(n_2),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_45),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_78),
.A2(n_86),
.B(n_89),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_85),
.Y(n_108)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_21),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_97),
.B1(n_61),
.B2(n_31),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_19),
.A3(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_33),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_98),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_33),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_57),
.B(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_102),
.B(n_124),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_98),
.B1(n_77),
.B2(n_75),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_115),
.Y(n_131)
);

OAI22x1_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_65),
.B1(n_57),
.B2(n_60),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_71),
.B1(n_101),
.B2(n_93),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_73),
.A2(n_24),
.B1(n_20),
.B2(n_18),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_18),
.B1(n_16),
.B2(n_15),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_120),
.B1(n_90),
.B2(n_96),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_16),
.B1(n_15),
.B2(n_3),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_123),
.B(n_83),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_125),
.B(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_3),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_85),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_86),
.B(n_90),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_124),
.B(n_123),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_78),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_137),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_84),
.C(n_76),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_113),
.C(n_118),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_78),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_133),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_74),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_144),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_135),
.B(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_74),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_125),
.B(n_114),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_101),
.B1(n_99),
.B2(n_80),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_139),
.A2(n_119),
.B1(n_121),
.B2(n_114),
.Y(n_163)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_140),
.B(n_153),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_4),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_141),
.A2(n_121),
.B(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_104),
.B(n_105),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_4),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_4),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_6),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_7),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_7),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_117),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_116),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_164),
.B(n_9),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_169),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_173),
.B1(n_141),
.B2(n_139),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_120),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_170),
.C(n_176),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_113),
.Y(n_169)
);

AO21x2_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_116),
.B(n_118),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_116),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_148),
.B(n_8),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_12),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_168),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_179),
.B(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_146),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_133),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_157),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_137),
.A3(n_128),
.B1(n_141),
.B2(n_132),
.C1(n_142),
.C2(n_131),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_191),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_145),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_194),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_131),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_195),
.C(n_176),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_134),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_152),
.C(n_10),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_9),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_198),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_162),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_206),
.C(n_208),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_203),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_173),
.B1(n_158),
.B2(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_170),
.C(n_164),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_173),
.C(n_158),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_189),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_173),
.B(n_159),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_197),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_205),
.B(n_179),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_219),
.C(n_222),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_221),
.B(n_223),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_201),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_R g218 ( 
.A1(n_212),
.A2(n_191),
.B(n_187),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_193),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_184),
.B1(n_175),
.B2(n_195),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_224),
.B1(n_213),
.B2(n_207),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_205),
.B(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_206),
.C(n_200),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_217),
.C(n_185),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_180),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_232),
.A2(n_216),
.B1(n_221),
.B2(n_202),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_161),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_234),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_162),
.Y(n_234)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_239),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_209),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_241),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_180),
.C(n_198),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_231),
.B1(n_229),
.B2(n_227),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_246),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_231),
.B1(n_11),
.B2(n_12),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_241),
.C(n_238),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_10),
.A3(n_243),
.B1(n_244),
.B2(n_233),
.C1(n_227),
.C2(n_237),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_247),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_244),
.Y(n_251)
);


endmodule