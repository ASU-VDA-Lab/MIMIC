module fake_jpeg_10957_n_133 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_29),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_3),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_3),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_48),
.B1(n_15),
.B2(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_11),
.B(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_8),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_17),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_21),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_25),
.A2(n_15),
.B1(n_21),
.B2(n_12),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_20),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_67),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_20),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_34),
.B(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_72),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_59),
.B(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_37),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_54),
.C(n_52),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_80),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_79),
.B(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_90),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_62),
.B(n_57),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_60),
.B(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_55),
.B1(n_66),
.B2(n_73),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_89),
.B1(n_76),
.B2(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_77),
.Y(n_100)
);

NOR2xp67_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_87),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_63),
.B1(n_54),
.B2(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_78),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_97),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_83),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_104),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_89),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

XOR2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_79),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_95),
.B1(n_99),
.B2(n_98),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_82),
.C(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_102),
.B(n_101),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_106),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_117),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_119),
.B(n_105),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_123),
.C(n_125),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_100),
.Y(n_125)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_128),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_117),
.C(n_118),
.Y(n_128)
);

AOI21x1_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_124),
.B(n_118),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_108),
.B(n_121),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_108),
.A3(n_130),
.B1(n_119),
.B2(n_94),
.C1(n_117),
.C2(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_126),
.Y(n_133)
);


endmodule