module fake_jpeg_28597_n_410 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_410);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_10),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_46),
.Y(n_90)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_10),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_10),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_23),
.A2(n_9),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_57),
.B(n_23),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_69),
.Y(n_116)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_67),
.Y(n_103)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_36),
.B(n_11),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_11),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_71),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_28),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_74),
.B(n_87),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx2_ASAP7_75t_R g122 ( 
.A(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_21),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_111),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_38),
.B1(n_50),
.B2(n_25),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_104),
.B1(n_77),
.B2(n_75),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_46),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_119),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_38),
.B1(n_25),
.B2(n_26),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_30),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_105),
.B(n_32),
.Y(n_161)
);

NAND2x1_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_43),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_71),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_37),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_129),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_61),
.A2(n_44),
.B1(n_26),
.B2(n_29),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_44),
.B1(n_25),
.B2(n_29),
.Y(n_144)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_152),
.Y(n_173)
);

BUFx2_ASAP7_75t_SL g134 ( 
.A(n_122),
.Y(n_134)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_51),
.B1(n_81),
.B2(n_84),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_135),
.A2(n_62),
.B1(n_83),
.B2(n_107),
.Y(n_184)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_136),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_143),
.A2(n_148),
.B1(n_103),
.B2(n_93),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_94),
.B1(n_110),
.B2(n_89),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_31),
.B(n_44),
.C(n_29),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_32),
.B(n_42),
.C(n_41),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_104),
.A2(n_73),
.B1(n_26),
.B2(n_38),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_98),
.B(n_35),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_157),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_59),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_77),
.Y(n_182)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_118),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_161),
.Y(n_178)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_163),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_187),
.B1(n_144),
.B2(n_156),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_117),
.C(n_31),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_145),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_154),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_186),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_184),
.A2(n_82),
.B1(n_142),
.B2(n_141),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_185),
.B(n_147),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_121),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_146),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_204),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_202),
.B1(n_208),
.B2(n_176),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_137),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_200),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_132),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_137),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_207),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_166),
.A2(n_131),
.B1(n_159),
.B2(n_140),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_211),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_185),
.A2(n_156),
.B(n_103),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_181),
.B(n_176),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_174),
.A3(n_187),
.B1(n_181),
.B2(n_175),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

AO22x1_ASAP7_75t_SL g207 ( 
.A1(n_175),
.A2(n_150),
.B1(n_107),
.B2(n_149),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_128),
.B1(n_93),
.B2(n_106),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_128),
.B1(n_106),
.B2(n_109),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_210),
.A2(n_182),
.B(n_176),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_174),
.B(n_120),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_212),
.A2(n_218),
.B(n_111),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_206),
.A2(n_177),
.B1(n_182),
.B2(n_164),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_219),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_211),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_221),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_216),
.A2(n_202),
.B1(n_209),
.B2(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_195),
.B(n_189),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_191),
.C(n_189),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_192),
.C(n_196),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_205),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_228),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_170),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_207),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_207),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_191),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_208),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_232),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_197),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_234),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_239),
.C(n_242),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_236),
.A2(n_243),
.B1(n_250),
.B2(n_254),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_221),
.B(n_203),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_238),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_206),
.C(n_194),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_222),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_183),
.C(n_157),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_180),
.B1(n_190),
.B2(n_168),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_220),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_223),
.Y(n_257)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_170),
.B(n_183),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_252),
.B(n_231),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_230),
.B1(n_232),
.B2(n_216),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_199),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_226),
.A2(n_167),
.B1(n_168),
.B2(n_180),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_190),
.B1(n_199),
.B2(n_167),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_214),
.B1(n_220),
.B2(n_245),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_162),
.C(n_153),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_212),
.C(n_213),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_263),
.Y(n_292)
);

AO22x1_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_213),
.B1(n_224),
.B2(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_253),
.Y(n_259)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_227),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_271),
.C(n_272),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_227),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_265),
.Y(n_305)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_215),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_215),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_217),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_256),
.C(n_246),
.Y(n_296)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_217),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_278),
.B(n_35),
.Y(n_302)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_248),
.A2(n_212),
.B1(n_190),
.B2(n_165),
.Y(n_280)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_251),
.Y(n_281)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

OA22x2_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_247),
.B1(n_234),
.B2(n_250),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_294),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_247),
.B1(n_238),
.B2(n_237),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_285),
.A2(n_287),
.B1(n_298),
.B2(n_303),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_267),
.A2(n_252),
.B(n_249),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_301),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_236),
.B1(n_255),
.B2(n_245),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_271),
.B(n_42),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_273),
.B(n_254),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_270),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_41),
.B1(n_37),
.B2(n_39),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_263),
.Y(n_299)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_261),
.B(n_39),
.Y(n_301)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_259),
.A2(n_139),
.B1(n_138),
.B2(n_112),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_304),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_257),
.C(n_272),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_279),
.C(n_280),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_311),
.C(n_317),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_326),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_270),
.C(n_258),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_321),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_136),
.C(n_125),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_170),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_319),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_172),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_172),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_295),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_322),
.Y(n_333)
);

XOR2x2_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_291),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_288),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_325),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_291),
.A2(n_171),
.B(n_152),
.Y(n_326)
);

NOR3xp33_ASAP7_75t_SL g327 ( 
.A(n_305),
.B(n_21),
.C(n_18),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_16),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_297),
.A2(n_131),
.B1(n_86),
.B2(n_85),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_328),
.A2(n_329),
.B1(n_151),
.B2(n_109),
.Y(n_339)
);

AOI211xp5_ASAP7_75t_SL g329 ( 
.A1(n_290),
.A2(n_172),
.B(n_171),
.C(n_2),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_308),
.A2(n_297),
.B1(n_289),
.B2(n_288),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_335),
.A2(n_304),
.B1(n_283),
.B2(n_322),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_296),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_312),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_289),
.C(n_300),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_338),
.C(n_340),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_300),
.C(n_290),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_339),
.A2(n_346),
.B1(n_333),
.B2(n_332),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_282),
.C(n_286),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_341),
.Y(n_352)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_342),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_282),
.C(n_284),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_345),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_282),
.C(n_284),
.Y(n_345)
);

OAI321xp33_ASAP7_75t_L g354 ( 
.A1(n_347),
.A2(n_327),
.A3(n_310),
.B1(n_315),
.B2(n_320),
.C(n_314),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_330),
.B(n_313),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_348),
.B(n_350),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_318),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_354),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_338),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_356),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_309),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_359),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_340),
.Y(n_359)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_283),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_360),
.B(n_344),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_171),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_357),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_352),
.A2(n_332),
.B1(n_331),
.B2(n_337),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_366),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_350),
.B(n_343),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_60),
.C(n_79),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_368),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_91),
.C(n_72),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_0),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_353),
.A2(n_171),
.B1(n_96),
.B2(n_91),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_371),
.A2(n_372),
.B(n_43),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_360),
.A2(n_96),
.B1(n_66),
.B2(n_43),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_374),
.B(n_376),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_348),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_351),
.C(n_43),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_377),
.B(n_378),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_43),
.C(n_8),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_4),
.Y(n_394)
);

AO22x1_ASAP7_75t_L g380 ( 
.A1(n_364),
.A2(n_6),
.B1(n_16),
.B2(n_2),
.Y(n_380)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_380),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_17),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_5),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_6),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_385),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_8),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_6),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_387),
.B(n_388),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_376),
.C(n_383),
.Y(n_388)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_390),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_385),
.B(n_8),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_391),
.A2(n_392),
.B(n_382),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_394),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_386),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_396),
.B(n_397),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_393),
.A2(n_4),
.B(n_14),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_400),
.A2(n_393),
.B(n_12),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_403),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_395),
.B(n_2),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_402),
.A2(n_399),
.B(n_398),
.Y(n_404)
);

AOI322xp5_ASAP7_75t_L g406 ( 
.A1(n_404),
.A2(n_3),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.C1(n_0),
.C2(n_1),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_407),
.A2(n_405),
.B(n_14),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_0),
.C(n_1),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_409),
.B(n_1),
.Y(n_410)
);


endmodule