module real_jpeg_4435_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_1),
.B(n_90),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_1),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_1),
.B(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_1),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_1),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_1),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_2),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_2),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_2),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_2),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_2),
.B(n_181),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_2),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_2),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_3),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_3),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_3),
.B(n_408),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_4),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_4),
.Y(n_191)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_4),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_5),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_5),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_5),
.B(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_5),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g299 ( 
.A(n_5),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_5),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_5),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_5),
.B(n_399),
.Y(n_398)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_7),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_7),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_7),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_7),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_7),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_7),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_7),
.B(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_8),
.Y(n_156)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_8),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_9),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_9),
.B(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_9),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_9),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_9),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_9),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_9),
.B(n_63),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_12),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_12),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_12),
.B(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_12),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_12),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_12),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_12),
.B(n_337),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_13),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_13),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_13),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_13),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_14),
.Y(n_163)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_14),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_14),
.Y(n_431)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_15),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_15),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_15),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_104),
.B(n_328),
.C(n_502),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_26),
.C(n_31),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_20),
.A2(n_31),
.B1(n_73),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_20),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_20),
.A2(n_83),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_20),
.B(n_226),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g502 ( 
.A(n_20),
.B(n_48),
.C(n_98),
.Y(n_502)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_25),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_25),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_26),
.A2(n_27),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_26),
.A2(n_27),
.B1(n_335),
.B2(n_341),
.Y(n_334)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_27),
.B(n_336),
.C(n_340),
.Y(n_483)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_31),
.A2(n_42),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_31),
.A2(n_73),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_31),
.B(n_144),
.C(n_148),
.Y(n_252)
);

OR2x2_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_32),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_34),
.Y(n_275)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_35),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_35),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_43),
.Y(n_42)
);

OR2x2_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_36),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_92),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_78),
.C(n_79),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_39),
.B(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_61),
.C(n_70),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_40),
.B(n_490),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_54),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_57),
.C(n_59),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.C(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_42),
.B(n_73),
.C(n_77),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_42),
.A2(n_74),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_42),
.B(n_115),
.C(n_118),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_42),
.A2(n_74),
.B1(n_478),
.B2(n_479),
.Y(n_477)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_46),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_46),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_46),
.Y(n_376)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_47),
.Y(n_251)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_47),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_48),
.A2(n_95),
.B1(n_96),
.B2(n_102),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_48),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_102),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_50),
.A2(n_51),
.B1(n_128),
.B2(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_50),
.A2(n_51),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_51),
.B(n_125),
.C(n_128),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_51),
.B(n_189),
.C(n_328),
.Y(n_482)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_53),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_61),
.B(n_70),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.C(n_69),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_62),
.Y(n_473)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_65),
.A2(n_66),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_66),
.B(n_133),
.C(n_236),
.Y(n_316)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_68),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_69),
.B(n_472),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_75),
.B2(n_77),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_75),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_75),
.A2(n_77),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_77),
.B(n_189),
.C(n_294),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_78),
.B(n_79),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_84),
.B1(n_85),
.B2(n_91),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_83),
.B(n_227),
.C(n_230),
.Y(n_289)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_88),
.C(n_91),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_97),
.A2(n_98),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_97),
.A2(n_98),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_97),
.B(n_349),
.C(n_354),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_98),
.B(n_311),
.C(n_316),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_99),
.Y(n_166)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_100),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_497),
.B(n_501),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_465),
.B(n_494),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_355),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_283),
.B(n_318),
.C(n_319),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_253),
.B(n_282),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_109),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_219),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_110),
.B(n_219),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_167),
.C(n_203),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_111),
.B(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_140),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_112),
.B(n_141),
.C(n_149),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_124),
.C(n_131),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_113),
.B(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_122),
.B(n_170),
.Y(n_423)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_124),
.A2(n_131),
.B1(n_132),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_124),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_125),
.B(n_261),
.Y(n_260)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_128),
.Y(n_262)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_133),
.A2(n_235),
.B1(n_236),
.B2(n_238),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_133),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_238),
.Y(n_276)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_149),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_145),
.B(n_189),
.Y(n_371)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_146),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_157),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_151),
.B(n_153),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_150),
.B(n_158),
.C(n_164),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_165),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_167),
.B(n_203),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_184),
.C(n_186),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_168),
.A2(n_184),
.B1(n_185),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_168),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_173),
.C(n_178),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_170),
.B(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_177),
.B1(n_178),
.B2(n_183),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_177),
.A2(n_178),
.B1(n_298),
.B2(n_302),
.Y(n_297)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_178),
.B(n_236),
.C(n_299),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_186),
.B(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.C(n_198),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_187),
.A2(n_188),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_189),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_189),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_189),
.A2(n_291),
.B1(n_328),
.B2(n_331),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx8_ASAP7_75t_L g366 ( 
.A(n_191),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_192),
.A2(n_193),
.B1(n_198),
.B2(n_199),
.Y(n_453)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_197),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_197),
.Y(n_427)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_218),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_206),
.C(n_218),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_214),
.C(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_212),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_212),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_214),
.A2(n_336),
.B1(n_339),
.B2(n_340),
.Y(n_335)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_214),
.Y(n_340)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_220),
.B(n_222),
.C(n_239),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_239),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_232),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_224),
.B(n_225),
.C(n_232),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_235),
.A2(n_236),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_235),
.A2(n_236),
.B1(n_363),
.B2(n_364),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_236),
.B(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_245),
.B(n_247),
.C(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_252),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_280),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_254),
.B(n_280),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_259),
.C(n_277),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_255),
.A2(n_256),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_259),
.B(n_277),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.C(n_276),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_260),
.B(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_263),
.B(n_276),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_269),
.C(n_272),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_264),
.A2(n_265),
.B1(n_272),
.B2(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_269),
.B(n_383),
.Y(n_382)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_271),
.Y(n_408)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_272),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_273),
.B(n_375),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_273),
.B(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_284),
.B(n_320),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_286),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_321),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_286),
.B(n_321),
.Y(n_464)
);

FAx1_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_303),
.CI(n_317),
.CON(n_286),
.SN(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_297),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_289),
.B(n_290),
.C(n_297),
.Y(n_344)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_299),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_306),
.C(n_308),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_322),
.B(n_324),
.C(n_342),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_342),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_325),
.B(n_333),
.C(n_334),
.Y(n_474)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_335),
.Y(n_341)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_336),
.Y(n_339)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_345),
.B2(n_346),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_343),
.B(n_347),
.C(n_348),
.Y(n_484)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

AO22x1_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_353),
.Y(n_354)
);

OAI31xp33_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_461),
.A3(n_462),
.B(n_464),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_455),
.B(n_460),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_442),
.B(n_454),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_402),
.B(n_441),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_385),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_360),
.B(n_385),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_372),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_361),
.B(n_373),
.C(n_382),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_367),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_362),
.B(n_368),
.C(n_371),
.Y(n_450)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_382),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_377),
.C(n_380),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_374),
.B(n_387),
.Y(n_386)
);

INVx11_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_377),
.A2(n_378),
.B1(n_380),
.B2(n_381),
.Y(n_387)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.C(n_401),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_386),
.B(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_388),
.A2(n_389),
.B1(n_401),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_397),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_390),
.A2(n_391),
.B1(n_397),
.B2(n_398),
.Y(n_411)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_401),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_435),
.B(n_440),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_421),
.B(n_434),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_412),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_412),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_411),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_409),
.C(n_411),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_418),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_413),
.A2(n_414),
.B1(n_418),
.B2(n_419),
.Y(n_432)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_419),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_428),
.B(n_433),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx8_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_432),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_429),
.B(n_432),
.Y(n_433)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_437),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_444),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_450),
.C(n_451),
.Y(n_459)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_459),
.Y(n_460)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_457),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_491),
.Y(n_465)
);

OAI21xp33_ASAP7_75t_L g494 ( 
.A1(n_466),
.A2(n_495),
.B(n_496),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_485),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_467),
.B(n_485),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_475),
.C(n_484),
.Y(n_467)
);

FAx1_ASAP7_75t_SL g493 ( 
.A(n_468),
.B(n_475),
.CI(n_484),
.CON(n_493),
.SN(n_493)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_474),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_471),
.C(n_474),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_477),
.B1(n_480),
.B2(n_481),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_482),
.C(n_483),
.Y(n_488)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_488),
.C(n_489),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_493),
.Y(n_495)
);

BUFx24_ASAP7_75t_SL g503 ( 
.A(n_493),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_500),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_500),
.Y(n_501)
);


endmodule