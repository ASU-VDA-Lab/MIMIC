module fake_jpeg_10342_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_4),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_1),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_5),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_18),
.B(n_19),
.Y(n_20)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

AO22x1_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_13),
.A2(n_6),
.B(n_7),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_19),
.B(n_18),
.C(n_16),
.Y(n_25)
);

AOI221xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_28),
.B1(n_19),
.B2(n_17),
.C(n_16),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_14),
.C(n_16),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_27),
.B(n_29),
.Y(n_31)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_32),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_10),
.B1(n_7),
.B2(n_12),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_22),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_35),
.B1(n_10),
.B2(n_25),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_38),
.B1(n_3),
.B2(n_4),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_31),
.C(n_17),
.Y(n_38)
);

AOI211xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_0),
.B(n_4),
.C(n_20),
.Y(n_40)
);


endmodule