module fake_jpeg_27083_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_20),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_11),
.B(n_20),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_13),
.B1(n_19),
.B2(n_12),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_16),
.B1(n_17),
.B2(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_31),
.B1(n_19),
.B2(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_37),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_25),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_41),
.C(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_42),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_12),
.B1(n_27),
.B2(n_11),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_13),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_48),
.B1(n_36),
.B2(n_44),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_46),
.B(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_18),
.B1(n_14),
.B2(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_36),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_57),
.B1(n_50),
.B2(n_49),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_36),
.B(n_34),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_58),
.B(n_44),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_14),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_8),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_61),
.B(n_63),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_8),
.C(n_3),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_2),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_69),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_66),
.C(n_5),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_7),
.C(n_70),
.Y(n_72)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_72),
.Y(n_73)
);


endmodule