module fake_jpeg_11229_n_630 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_630);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_630;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_539;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_5),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_2),
.B(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_78),
.Y(n_176)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_81),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_82),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_83),
.Y(n_184)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_85),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_35),
.B(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_96),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_35),
.B(n_10),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_87),
.A2(n_99),
.B(n_111),
.C(n_112),
.Y(n_173)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_90),
.Y(n_182)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_92),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_93),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_94),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_10),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_97),
.Y(n_187)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_10),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_103),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_9),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_60),
.B(n_9),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_19),
.B(n_11),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_117),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

CKINVDCx6p67_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_19),
.B(n_11),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_25),
.Y(n_121)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_20),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_49),
.Y(n_136)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_25),
.Y(n_127)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_30),
.Y(n_128)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_30),
.Y(n_129)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_136),
.B(n_151),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_60),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_141),
.B(n_160),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_22),
.B1(n_58),
.B2(n_42),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_146),
.A2(n_149),
.B1(n_155),
.B2(n_157),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_74),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_96),
.B(n_22),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_85),
.A2(n_31),
.B1(n_33),
.B2(n_45),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_156),
.B(n_170),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_112),
.A2(n_46),
.B1(n_58),
.B2(n_42),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_93),
.B(n_46),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_82),
.B(n_52),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_165),
.B(n_90),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_83),
.B(n_52),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_92),
.B(n_55),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_171),
.B(n_211),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_62),
.A2(n_31),
.B1(n_33),
.B2(n_49),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_174),
.A2(n_204),
.B1(n_59),
.B2(n_53),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_103),
.A2(n_55),
.B1(n_27),
.B2(n_34),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_209),
.B(n_0),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_64),
.A2(n_34),
.B1(n_27),
.B2(n_32),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_201),
.A2(n_213),
.B1(n_59),
.B2(n_53),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_65),
.A2(n_34),
.B1(n_32),
.B2(n_27),
.Y(n_204)
);

INVx6_ASAP7_75t_SL g206 ( 
.A(n_126),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_121),
.B(n_32),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_208),
.B(n_0),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_68),
.A2(n_56),
.B1(n_14),
.B2(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_102),
.B(n_13),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_67),
.A2(n_53),
.B1(n_47),
.B2(n_20),
.Y(n_213)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_105),
.Y(n_214)
);

BUFx2_ASAP7_75t_SL g220 ( 
.A(n_214),
.Y(n_220)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_134),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_216),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_164),
.A2(n_63),
.B1(n_128),
.B2(n_127),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_217),
.A2(n_253),
.B1(n_256),
.B2(n_273),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_218),
.Y(n_343)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_223),
.Y(n_311)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_224),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_204),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_226),
.B(n_240),
.Y(n_302)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_227),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_228),
.Y(n_325)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_143),
.Y(n_229)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_229),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_230),
.A2(n_231),
.B(n_262),
.Y(n_348)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_140),
.B(n_129),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_232),
.Y(n_339)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_144),
.Y(n_234)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_234),
.Y(n_298)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_152),
.B(n_104),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_236),
.B(n_261),
.Y(n_307)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_238),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_175),
.Y(n_239)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_239),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_149),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_137),
.Y(n_241)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_168),
.Y(n_242)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_242),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_243),
.Y(n_300)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_251),
.Y(n_296)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_131),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_245),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_175),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_247),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_188),
.B(n_116),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_248),
.B(n_254),
.C(n_287),
.Y(n_297)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_131),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_249),
.B(n_252),
.Y(n_310)
);

BUFx2_ASAP7_75t_SL g251 ( 
.A(n_195),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_198),
.A2(n_101),
.B1(n_95),
.B2(n_107),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_180),
.B(n_78),
.C(n_81),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_199),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_255),
.B(n_258),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_158),
.Y(n_256)
);

O2A1O1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_173),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g323 ( 
.A1(n_257),
.A2(n_269),
.B1(n_183),
.B2(n_167),
.Y(n_323)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

INVx11_ASAP7_75t_L g259 ( 
.A(n_134),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_259),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_155),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_260),
.B(n_264),
.Y(n_349)
);

OR2x2_ASAP7_75t_SL g262 ( 
.A(n_148),
.B(n_59),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_172),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_263),
.B(n_266),
.Y(n_334)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_202),
.Y(n_264)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_166),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_267),
.A2(n_278),
.B1(n_279),
.B2(n_288),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_130),
.B(n_14),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_268),
.B(n_271),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_192),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_212),
.B1(n_138),
.B2(n_167),
.Y(n_299)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_158),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_145),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_275),
.Y(n_295)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_172),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_147),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_277),
.Y(n_292)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_154),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_196),
.A2(n_59),
.B1(n_53),
.B2(n_47),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_159),
.A2(n_59),
.B1(n_53),
.B2(n_47),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_163),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_280),
.A2(n_289),
.B1(n_290),
.B2(n_183),
.Y(n_314)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_161),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_282),
.Y(n_301)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_166),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_185),
.B(n_5),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_283),
.B(n_285),
.Y(n_313)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_162),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_286),
.Y(n_316)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_135),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_140),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_139),
.B(n_47),
.C(n_20),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_159),
.A2(n_47),
.B1(n_20),
.B2(n_7),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_191),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_184),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_236),
.A2(n_174),
.B1(n_163),
.B2(n_169),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_293),
.A2(n_324),
.B1(n_330),
.B2(n_331),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_299),
.A2(n_315),
.B1(n_329),
.B2(n_238),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

AO21x2_ASAP7_75t_L g315 ( 
.A1(n_231),
.A2(n_214),
.B(n_142),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_262),
.B(n_177),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_327),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_323),
.B(n_315),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_267),
.A2(n_169),
.B1(n_176),
.B2(n_186),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_272),
.B(n_215),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_233),
.B(n_193),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_333),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_228),
.A2(n_269),
.B1(n_257),
.B2(n_254),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_230),
.A2(n_186),
.B1(n_176),
.B2(n_182),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_265),
.A2(n_287),
.B1(n_250),
.B2(n_235),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_219),
.A2(n_182),
.B1(n_194),
.B2(n_187),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_332),
.A2(n_338),
.B1(n_345),
.B2(n_220),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_222),
.B(n_189),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_241),
.B(n_205),
.C(n_142),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_347),
.C(n_218),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_237),
.A2(n_194),
.B1(n_153),
.B2(n_178),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_229),
.B(n_5),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_340),
.B(n_341),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_234),
.B(n_6),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_7),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_342),
.B(n_346),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_263),
.A2(n_142),
.B1(n_184),
.B2(n_20),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_225),
.B(n_7),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_248),
.B(n_12),
.C(n_13),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_348),
.A2(n_221),
.B(n_290),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_351),
.A2(n_357),
.B(n_315),
.Y(n_424)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_343),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_352),
.Y(n_402)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_353),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_348),
.A2(n_242),
.B(n_248),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_354),
.A2(n_384),
.B(n_387),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_328),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_355),
.B(n_359),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_325),
.A2(n_329),
.B(n_302),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_282),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_358),
.B(n_361),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_313),
.B(n_247),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_327),
.A2(n_307),
.B1(n_318),
.B2(n_297),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_360),
.A2(n_385),
.B1(n_388),
.B2(n_317),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_331),
.B(n_244),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_362),
.B(n_368),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_363),
.A2(n_395),
.B1(n_334),
.B2(n_309),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_293),
.A2(n_275),
.B1(n_232),
.B2(n_224),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_364),
.A2(n_377),
.B1(n_380),
.B2(n_389),
.Y(n_423)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_295),
.Y(n_366)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_366),
.Y(n_409)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_297),
.B(n_259),
.C(n_216),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_301),
.Y(n_369)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_370),
.B(n_372),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_296),
.Y(n_371)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_296),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_344),
.B(n_310),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_394),
.Y(n_397)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_316),
.Y(n_375)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_375),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_223),
.C(n_280),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_376),
.B(n_391),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_324),
.A2(n_273),
.B1(n_256),
.B2(n_266),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_316),
.Y(n_378)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_330),
.A2(n_249),
.B1(n_245),
.B2(n_289),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_326),
.Y(n_381)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_304),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_382),
.Y(n_405)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_383),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_294),
.A2(n_323),
.B1(n_345),
.B2(n_347),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_299),
.A2(n_239),
.B1(n_246),
.B2(n_16),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_323),
.A2(n_12),
.B(n_15),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_315),
.A2(n_17),
.B1(n_336),
.B2(n_323),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_340),
.A2(n_17),
.B1(n_342),
.B2(n_341),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_291),
.B(n_17),
.C(n_333),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_322),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_392),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_291),
.B(n_296),
.C(n_300),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_393),
.B(n_298),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_319),
.B(n_292),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_379),
.A2(n_312),
.B1(n_309),
.B2(n_339),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_396),
.A2(n_421),
.B1(n_425),
.B2(n_379),
.Y(n_438)
);

INVx5_ASAP7_75t_SL g399 ( 
.A(n_358),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_399),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_346),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_433),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_358),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_407),
.B(n_408),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_393),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_356),
.A2(n_315),
.B1(n_314),
.B2(n_292),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_410),
.A2(n_395),
.B1(n_387),
.B2(n_385),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_362),
.B(n_303),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_413),
.C(n_419),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_360),
.B(n_322),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_352),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_415),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_370),
.B(n_298),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_386),
.B(n_367),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_422),
.B(n_390),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_424),
.A2(n_430),
.B(n_351),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_388),
.A2(n_395),
.B1(n_350),
.B2(n_378),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_357),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_428),
.B(n_382),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_369),
.B(n_300),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_354),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_433),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_436),
.B(n_445),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_438),
.A2(n_463),
.B1(n_410),
.B2(n_423),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_439),
.B(n_442),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_440),
.A2(n_458),
.B(n_461),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_368),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_444),
.C(n_447),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_376),
.C(n_373),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_399),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_397),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_457),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_367),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_401),
.B(n_386),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_448),
.B(n_450),
.C(n_454),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_449),
.B(n_427),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_384),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_400),
.B(n_366),
.Y(n_451)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_417),
.B(n_353),
.Y(n_452)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_429),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_453),
.B(n_466),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_411),
.B(n_371),
.C(n_350),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_455),
.A2(n_398),
.B1(n_421),
.B2(n_431),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_356),
.C(n_391),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_469),
.C(n_427),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_429),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_424),
.A2(n_380),
.B(n_361),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_432),
.Y(n_459)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_459),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_429),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_467),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_364),
.B(n_377),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_425),
.A2(n_389),
.B1(n_392),
.B2(n_383),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_405),
.Y(n_464)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_464),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_381),
.Y(n_465)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_465),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_321),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_431),
.B(n_365),
.Y(n_468)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_468),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_422),
.B(n_305),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_472),
.A2(n_479),
.B1(n_484),
.B2(n_493),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_465),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_475),
.B(n_480),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_476),
.A2(n_496),
.B1(n_499),
.B2(n_437),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_436),
.A2(n_414),
.B1(n_406),
.B2(n_409),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_446),
.B(n_462),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_457),
.A2(n_414),
.B1(n_416),
.B2(n_398),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_468),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_485),
.B(n_487),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_486),
.B(n_490),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_452),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_448),
.Y(n_502)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_459),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_489),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_440),
.B(n_437),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_492),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_460),
.A2(n_404),
.B1(n_426),
.B2(n_418),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_441),
.B(n_404),
.C(n_426),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_498),
.C(n_454),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_455),
.A2(n_418),
.B1(n_432),
.B2(n_403),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_441),
.B(n_444),
.C(n_450),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_461),
.A2(n_403),
.B1(n_402),
.B2(n_405),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_456),
.B(n_415),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_501),
.B(n_402),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_502),
.B(n_503),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_439),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_504),
.B(n_520),
.Y(n_532)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_470),
.Y(n_506)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_506),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_507),
.A2(n_521),
.B1(n_495),
.B2(n_471),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_477),
.B(n_447),
.C(n_469),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_508),
.B(n_515),
.C(n_516),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_449),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_509),
.B(n_519),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_492),
.A2(n_445),
.B(n_458),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_511),
.B(n_518),
.Y(n_542)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_483),
.Y(n_512)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_512),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_471),
.A2(n_435),
.B(n_451),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_513),
.B(n_517),
.Y(n_545)
);

XNOR2x1_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_435),
.Y(n_514)
);

XNOR2x1_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_476),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_477),
.B(n_463),
.C(n_321),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_486),
.B(n_464),
.C(n_402),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_483),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_482),
.B(n_443),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_498),
.B(n_443),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_496),
.A2(n_311),
.B1(n_312),
.B2(n_343),
.Y(n_521)
);

XNOR2x2_ASAP7_75t_L g522 ( 
.A(n_484),
.B(n_308),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_522),
.B(n_481),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_495),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_528),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_472),
.A2(n_311),
.B1(n_308),
.B2(n_305),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_527),
.A2(n_499),
.B1(n_497),
.B2(n_491),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_494),
.B(n_490),
.C(n_493),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_479),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_529),
.A2(n_320),
.B1(n_306),
.B2(n_335),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_535),
.B(n_507),
.Y(n_569)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_536),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_524),
.A2(n_478),
.B1(n_497),
.B2(n_473),
.Y(n_537)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_537),
.Y(n_570)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_505),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_539),
.Y(n_565)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_530),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_SL g556 ( 
.A1(n_543),
.A2(n_551),
.B1(n_552),
.B2(n_553),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_510),
.B(n_500),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_544),
.Y(n_558)
);

INVxp33_ASAP7_75t_SL g546 ( 
.A(n_524),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_546),
.B(n_550),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_547),
.A2(n_502),
.B1(n_503),
.B2(n_521),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_527),
.A2(n_478),
.B1(n_473),
.B2(n_500),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_548),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_554),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_522),
.A2(n_491),
.B1(n_489),
.B2(n_474),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_526),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_525),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_525),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_533),
.Y(n_555)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_555),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_544),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_557),
.B(n_560),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_541),
.B(n_516),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_559),
.B(n_568),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_544),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_545),
.A2(n_513),
.B(n_514),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_561),
.A2(n_542),
.B(n_538),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_534),
.B(n_520),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_564),
.B(n_567),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_534),
.B(n_519),
.C(n_528),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_549),
.B(n_515),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_569),
.B(n_535),
.Y(n_584)
);

INVxp33_ASAP7_75t_L g581 ( 
.A(n_571),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_532),
.B(n_504),
.C(n_523),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_573),
.B(n_532),
.C(n_523),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_550),
.B(n_508),
.Y(n_574)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_574),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_576),
.A2(n_580),
.B(n_561),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_577),
.B(n_579),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_573),
.B(n_540),
.C(n_531),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_572),
.B(n_537),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_567),
.B(n_540),
.C(n_531),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_582),
.B(n_588),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_584),
.B(n_587),
.Y(n_603)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_565),
.Y(n_586)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_586),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_562),
.B(n_547),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_571),
.B(n_509),
.C(n_548),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_556),
.Y(n_589)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_589),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_580),
.A2(n_566),
.B1(n_570),
.B2(n_572),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_592),
.B(n_594),
.Y(n_607)
);

OAI21xp33_ASAP7_75t_L g593 ( 
.A1(n_578),
.A2(n_560),
.B(n_558),
.Y(n_593)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_593),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_576),
.A2(n_566),
.B1(n_570),
.B2(n_563),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_595),
.B(n_600),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_583),
.B(n_558),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_597),
.B(n_581),
.Y(n_610)
);

NAND2x1_ASAP7_75t_SL g600 ( 
.A(n_588),
.B(n_569),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_575),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_601),
.B(n_602),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_590),
.B(n_562),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_598),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_606),
.B(n_608),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_599),
.B(n_585),
.Y(n_608)
);

AO21x1_ASAP7_75t_L g609 ( 
.A1(n_596),
.A2(n_581),
.B(n_563),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_609),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_610),
.B(n_612),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_603),
.B(n_577),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_603),
.B(n_582),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_613),
.B(n_584),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_605),
.B(n_579),
.C(n_595),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_614),
.B(n_618),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_604),
.A2(n_593),
.B(n_591),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_615),
.A2(n_617),
.B(n_619),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_604),
.A2(n_600),
.B(n_594),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_621),
.A2(n_622),
.B(n_624),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_616),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_620),
.B(n_611),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_623),
.A2(n_607),
.B(n_592),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_625),
.B(n_587),
.Y(n_627)
);

OAI321xp33_ASAP7_75t_L g628 ( 
.A1(n_627),
.A2(n_626),
.A3(n_536),
.B1(n_320),
.B2(n_334),
.C(n_335),
.Y(n_628)
);

BUFx24_ASAP7_75t_SL g629 ( 
.A(n_628),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_629),
.B(n_334),
.C(n_306),
.Y(n_630)
);


endmodule