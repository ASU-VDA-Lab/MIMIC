module fake_netlist_6_911_n_937 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_937);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_937;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_671;
wire n_607;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_703;
wire n_578;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_742;
wire n_532;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_624;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_527;
wire n_608;
wire n_261;
wire n_683;
wire n_474;
wire n_420;
wire n_620;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_652;
wire n_553;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_71),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_128),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_88),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_30),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_173),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_150),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_77),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_49),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_47),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_65),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_28),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_139),
.Y(n_190)
);

INVxp33_ASAP7_75t_SL g191 ( 
.A(n_161),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_169),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_119),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_50),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_16),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_75),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_42),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_89),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_28),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_68),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_13),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_81),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_57),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_62),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_122),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_72),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_83),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_51),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_46),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_55),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_172),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_66),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_113),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_19),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_20),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_100),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_58),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_165),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_93),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_69),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_53),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_115),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_60),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_8),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_9),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_129),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_123),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_24),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_26),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_3),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_102),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_8),
.Y(n_241)
);

BUFx2_ASAP7_75t_SL g242 ( 
.A(n_106),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_20),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_52),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_54),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_31),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_91),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_192),
.B(n_214),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_0),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_197),
.B(n_0),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_174),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_192),
.B(n_1),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_205),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_214),
.B(n_1),
.Y(n_261)
);

AND2x4_ASAP7_75t_L g262 ( 
.A(n_204),
.B(n_170),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_241),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_191),
.B(n_2),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g265 ( 
.A(n_204),
.B(n_32),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_191),
.B(n_246),
.Y(n_266)
);

BUFx8_ASAP7_75t_SL g267 ( 
.A(n_237),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_180),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_2),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_3),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_222),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g274 ( 
.A(n_202),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_166),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_4),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_233),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_224),
.B(n_4),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_233),
.B(n_5),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_175),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_186),
.B(n_5),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_189),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_194),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_178),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_202),
.B(n_6),
.Y(n_286)
);

BUFx8_ASAP7_75t_L g287 ( 
.A(n_196),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_199),
.B(n_6),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_201),
.B(n_164),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_208),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_215),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_234),
.B(n_7),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_219),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_221),
.B(n_33),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_241),
.B(n_7),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_226),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_235),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_236),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_176),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_255),
.A2(n_237),
.B1(n_240),
.B2(n_210),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_247),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_286),
.A2(n_188),
.B1(n_203),
.B2(n_243),
.Y(n_305)
);

AO22x2_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_242),
.B1(n_10),
.B2(n_11),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_177),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_267),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_179),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_220),
.B1(n_207),
.B2(n_240),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_266),
.A2(n_207),
.B1(n_210),
.B2(n_225),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_264),
.A2(n_225),
.B1(n_244),
.B2(n_231),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_270),
.A2(n_245),
.B1(n_230),
.B2(n_229),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_263),
.B(n_9),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_181),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_R g317 ( 
.A1(n_263),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_182),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_L g321 ( 
.A1(n_258),
.A2(n_228),
.B1(n_218),
.B2(n_216),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_278),
.B(n_183),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_R g323 ( 
.A1(n_282),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_L g324 ( 
.A1(n_258),
.A2(n_213),
.B1(n_212),
.B2(n_211),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_255),
.A2(n_209),
.B1(n_206),
.B2(n_200),
.Y(n_327)
);

NAND2xp33_ASAP7_75t_SL g328 ( 
.A(n_295),
.B(n_184),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_251),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_248),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_284),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_268),
.A2(n_198),
.B1(n_193),
.B2(n_190),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_271),
.A2(n_187),
.B1(n_185),
.B2(n_16),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_278),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_251),
.B(n_15),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_278),
.B(n_34),
.Y(n_337)
);

AO22x2_ASAP7_75t_L g338 ( 
.A1(n_256),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_278),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_L g340 ( 
.A1(n_271),
.A2(n_272),
.B1(n_292),
.B2(n_274),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_290),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_252),
.B(n_35),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_290),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_L g344 ( 
.A1(n_272),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_256),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_276),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_252),
.B(n_27),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_252),
.B(n_36),
.Y(n_348)
);

AO22x2_ASAP7_75t_L g349 ( 
.A1(n_276),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_278),
.B(n_38),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_250),
.Y(n_351)
);

AO22x2_ASAP7_75t_L g352 ( 
.A1(n_280),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_278),
.B(n_41),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_L g354 ( 
.A1(n_292),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_280),
.A2(n_48),
.B1(n_56),
.B2(n_59),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_261),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_278),
.A2(n_67),
.B1(n_70),
.B2(n_73),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_262),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_299),
.B(n_79),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_262),
.A2(n_265),
.B1(n_275),
.B2(n_279),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_304),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_R g365 ( 
.A(n_307),
.B(n_262),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_329),
.A2(n_294),
.B(n_289),
.Y(n_366)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_353),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_302),
.B(n_262),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_340),
.B(n_248),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_320),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_309),
.B(n_248),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_326),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_303),
.B(n_249),
.Y(n_374)
);

NAND2x1p5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_265),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_327),
.B(n_249),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_315),
.B(n_249),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_302),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_311),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_319),
.B(n_274),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_314),
.B(n_299),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_312),
.B(n_274),
.Y(n_384)
);

BUFx6f_ASAP7_75t_SL g385 ( 
.A(n_308),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_277),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_330),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_328),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_332),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_321),
.B(n_265),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_342),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_310),
.B(n_265),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_359),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_R g400 ( 
.A(n_336),
.B(n_275),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_333),
.B(n_299),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_324),
.B(n_275),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_313),
.B(n_275),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_305),
.B(n_289),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_334),
.B(n_289),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_322),
.A2(n_294),
.B(n_289),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_337),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_345),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_R g411 ( 
.A(n_352),
.B(n_294),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_356),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_345),
.B(n_288),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_356),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_349),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_335),
.B(n_294),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_344),
.B(n_290),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_306),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_306),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_358),
.A2(n_293),
.B(n_291),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_339),
.B(n_291),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_357),
.Y(n_424)
);

NAND2x1p5_ASAP7_75t_L g425 ( 
.A(n_346),
.B(n_281),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_338),
.B(n_300),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_338),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_354),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_317),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_323),
.B(n_80),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_302),
.B(n_82),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_302),
.B(n_84),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_302),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_375),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_254),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_300),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_375),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_425),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_405),
.B(n_300),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_385),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_372),
.B(n_85),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_370),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_423),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_373),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_366),
.B(n_281),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_401),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_406),
.B(n_254),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_386),
.B(n_260),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_424),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_361),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_395),
.B(n_281),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_382),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_386),
.B(n_260),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_363),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_399),
.B(n_281),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_407),
.B(n_273),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_423),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_422),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_407),
.B(n_273),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_367),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_409),
.B(n_296),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_364),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_298),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_414),
.B(n_404),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_396),
.B(n_296),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_367),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_402),
.A2(n_293),
.B1(n_291),
.B2(n_296),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_365),
.Y(n_479)
);

AND2x2_ASAP7_75t_SL g480 ( 
.A(n_403),
.B(n_402),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_383),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_403),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_404),
.B(n_298),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_389),
.B(n_293),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_367),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_394),
.A2(n_296),
.B(n_250),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_427),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_418),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_367),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_418),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_367),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_408),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_420),
.B(n_284),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_421),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_374),
.B(n_284),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_428),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_377),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_419),
.B(n_250),
.Y(n_500)
);

AND2x2_ASAP7_75t_SL g501 ( 
.A(n_416),
.B(n_297),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_417),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_381),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_371),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_387),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_398),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_374),
.B(n_376),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_430),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_410),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_376),
.B(n_297),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_397),
.B(n_369),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_384),
.B(n_297),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_368),
.Y(n_514)
);

AND2x2_ASAP7_75t_SL g515 ( 
.A(n_411),
.B(n_297),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_400),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_284),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_450),
.B(n_434),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_439),
.B(n_380),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_287),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_455),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_453),
.Y(n_522)
);

INVx6_ASAP7_75t_L g523 ( 
.A(n_471),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_287),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_457),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_506),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_457),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_439),
.B(n_379),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_493),
.B(n_287),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_435),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_435),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_435),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_453),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_450),
.B(n_432),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_493),
.B(n_287),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_446),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_452),
.B(n_433),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_439),
.B(n_86),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_453),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_497),
.B(n_87),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_497),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_497),
.B(n_90),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_482),
.B(n_385),
.Y(n_544)
);

BUFx12f_ASAP7_75t_L g545 ( 
.A(n_443),
.Y(n_545)
);

CKINVDCx8_ASAP7_75t_R g546 ( 
.A(n_500),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_462),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_437),
.B(n_297),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_499),
.B(n_92),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_437),
.B(n_297),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_462),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_446),
.Y(n_552)
);

BUFx5_ASAP7_75t_L g553 ( 
.A(n_476),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_489),
.B(n_284),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_446),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_482),
.B(n_431),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_489),
.B(n_284),
.Y(n_557)
);

BUFx12f_ASAP7_75t_L g558 ( 
.A(n_438),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_498),
.B(n_94),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_462),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_448),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_491),
.B(n_269),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_499),
.B(n_95),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_463),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_452),
.B(n_96),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_448),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_448),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_452),
.B(n_458),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_498),
.B(n_97),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_458),
.B(n_461),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_498),
.B(n_98),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_491),
.B(n_269),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_499),
.B(n_99),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_480),
.B(n_269),
.Y(n_574)
);

CKINVDCx8_ASAP7_75t_R g575 ( 
.A(n_500),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_510),
.B(n_101),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_463),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_480),
.B(n_269),
.Y(n_578)
);

NOR2x1_ASAP7_75t_L g579 ( 
.A(n_463),
.B(n_103),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_500),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_522),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_523),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_558),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_580),
.Y(n_584)
);

BUFx2_ASAP7_75t_SL g585 ( 
.A(n_527),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_580),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_523),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_546),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_545),
.Y(n_589)
);

BUFx12f_ASAP7_75t_L g590 ( 
.A(n_529),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_522),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_522),
.Y(n_592)
);

CKINVDCx16_ASAP7_75t_R g593 ( 
.A(n_519),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_568),
.B(n_480),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_519),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_540),
.Y(n_596)
);

BUFx4f_ASAP7_75t_L g597 ( 
.A(n_540),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_537),
.Y(n_598)
);

BUFx2_ASAP7_75t_SL g599 ( 
.A(n_540),
.Y(n_599)
);

INVx5_ASAP7_75t_SL g600 ( 
.A(n_571),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_561),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_547),
.Y(n_602)
);

INVx3_ASAP7_75t_SL g603 ( 
.A(n_529),
.Y(n_603)
);

INVx6_ASAP7_75t_SL g604 ( 
.A(n_571),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_518),
.Y(n_605)
);

BUFx4_ASAP7_75t_SL g606 ( 
.A(n_576),
.Y(n_606)
);

INVx5_ASAP7_75t_SL g607 ( 
.A(n_549),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_535),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_577),
.Y(n_609)
);

BUFx12f_ASAP7_75t_L g610 ( 
.A(n_549),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_552),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_570),
.B(n_447),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_577),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_538),
.B(n_510),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_547),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_547),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_521),
.B(n_461),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_551),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_555),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_580),
.Y(n_620)
);

CKINVDCx16_ASAP7_75t_R g621 ( 
.A(n_556),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_525),
.B(n_461),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_565),
.A2(n_501),
.B1(n_464),
.B2(n_447),
.Y(n_623)
);

INVx5_ASAP7_75t_SL g624 ( 
.A(n_563),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_575),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_551),
.Y(n_626)
);

INVx3_ASAP7_75t_SL g627 ( 
.A(n_563),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_551),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_564),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_564),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_526),
.B(n_466),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_564),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_560),
.Y(n_633)
);

BUFx4f_ASAP7_75t_SL g634 ( 
.A(n_590),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_585),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_623),
.A2(n_501),
.B1(n_515),
.B2(n_445),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_598),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_594),
.A2(n_507),
.B1(n_512),
.B2(n_464),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_594),
.A2(n_507),
.B1(n_512),
.B2(n_501),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_614),
.A2(n_507),
.B1(n_512),
.B2(n_473),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_611),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_619),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_597),
.Y(n_643)
);

AOI21xp33_ASAP7_75t_L g644 ( 
.A1(n_623),
.A2(n_511),
.B(n_520),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_601),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_589),
.Y(n_646)
);

BUFx5_ASAP7_75t_L g647 ( 
.A(n_610),
.Y(n_647)
);

OAI22xp33_ASAP7_75t_L g648 ( 
.A1(n_614),
.A2(n_514),
.B1(n_445),
.B2(n_516),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_612),
.B(n_473),
.Y(n_649)
);

INVx6_ASAP7_75t_L g650 ( 
.A(n_596),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_589),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_605),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_612),
.A2(n_473),
.B1(n_445),
.B2(n_515),
.Y(n_653)
);

BUFx4f_ASAP7_75t_SL g654 ( 
.A(n_590),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_621),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_608),
.A2(n_515),
.B1(n_441),
.B2(n_516),
.Y(n_656)
);

BUFx8_ASAP7_75t_SL g657 ( 
.A(n_583),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_601),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_617),
.B(n_466),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_603),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_595),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_632),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_606),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_632),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_633),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_609),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_604),
.A2(n_441),
.B1(n_514),
.B2(n_539),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_581),
.Y(n_668)
);

CKINVDCx11_ASAP7_75t_R g669 ( 
.A(n_603),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_604),
.A2(n_539),
.B1(n_479),
.B2(n_458),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_613),
.Y(n_671)
);

INVx8_ASAP7_75t_L g672 ( 
.A(n_596),
.Y(n_672)
);

INVx4_ASAP7_75t_SL g673 ( 
.A(n_627),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_581),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_604),
.A2(n_479),
.B1(n_505),
.B2(n_504),
.Y(n_675)
);

INVx3_ASAP7_75t_SL g676 ( 
.A(n_593),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_596),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_627),
.A2(n_438),
.B1(n_506),
.B2(n_505),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_582),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_610),
.A2(n_505),
.B1(n_504),
.B2(n_524),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_582),
.B(n_466),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_600),
.A2(n_509),
.B1(n_436),
.B2(n_440),
.Y(n_682)
);

CKINVDCx11_ASAP7_75t_R g683 ( 
.A(n_587),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_587),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_643),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_645),
.Y(n_686)
);

CKINVDCx11_ASAP7_75t_R g687 ( 
.A(n_651),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_648),
.A2(n_544),
.B1(n_569),
.B2(n_559),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_655),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_671),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_638),
.A2(n_483),
.B1(n_440),
.B2(n_436),
.Y(n_691)
);

OAI222xp33_ASAP7_75t_L g692 ( 
.A1(n_639),
.A2(n_631),
.B1(n_622),
.B2(n_511),
.C1(n_485),
.C2(n_528),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_640),
.A2(n_483),
.B1(n_436),
.B2(n_440),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_SL g694 ( 
.A1(n_667),
.A2(n_670),
.B(n_636),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_678),
.A2(n_483),
.B1(n_485),
.B2(n_543),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g696 ( 
.A(n_675),
.B(n_536),
.C(n_530),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_649),
.B(n_600),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_649),
.A2(n_624),
.B1(n_607),
.B2(n_600),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_681),
.A2(n_485),
.B1(n_543),
.B2(n_541),
.Y(n_699)
);

NOR2x1_ASAP7_75t_R g700 ( 
.A(n_669),
.B(n_599),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_672),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_SL g702 ( 
.A1(n_636),
.A2(n_465),
.B1(n_541),
.B2(n_624),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_SL g703 ( 
.A1(n_634),
.A2(n_465),
.B1(n_624),
.B2(n_607),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_661),
.A2(n_471),
.B1(n_481),
.B2(n_573),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_652),
.B(n_607),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_659),
.A2(n_471),
.B1(n_481),
.B2(n_573),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_659),
.B(n_509),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_662),
.B(n_481),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_657),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_664),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_637),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_672),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_684),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_641),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_680),
.A2(n_451),
.B1(n_509),
.B2(n_542),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_643),
.Y(n_716)
);

BUFx4f_ASAP7_75t_SL g717 ( 
.A(n_676),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_666),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_679),
.B(n_451),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_653),
.A2(n_451),
.B1(n_442),
.B2(n_484),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_642),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_676),
.B(n_442),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_SL g723 ( 
.A1(n_654),
.A2(n_487),
.B1(n_444),
.B2(n_625),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_682),
.A2(n_656),
.B1(n_635),
.B2(n_660),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_658),
.B(n_442),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_665),
.B(n_629),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_644),
.A2(n_484),
.B1(n_513),
.B2(n_444),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_644),
.A2(n_484),
.B1(n_513),
.B2(n_444),
.Y(n_728)
);

INVx5_ASAP7_75t_SL g729 ( 
.A(n_643),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_647),
.A2(n_444),
.B1(n_459),
.B2(n_470),
.Y(n_730)
);

BUFx4f_ASAP7_75t_SL g731 ( 
.A(n_647),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_647),
.A2(n_444),
.B1(n_459),
.B2(n_470),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_683),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_668),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_650),
.A2(n_588),
.B1(n_625),
.B2(n_560),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_647),
.A2(n_469),
.B1(n_490),
.B2(n_492),
.Y(n_736)
);

AOI222xp33_ASAP7_75t_L g737 ( 
.A1(n_673),
.A2(n_495),
.B1(n_494),
.B2(n_487),
.C1(n_502),
.C2(n_503),
.Y(n_737)
);

BUFx8_ASAP7_75t_L g738 ( 
.A(n_647),
.Y(n_738)
);

BUFx4f_ASAP7_75t_SL g739 ( 
.A(n_647),
.Y(n_739)
);

OAI21xp33_ASAP7_75t_L g740 ( 
.A1(n_646),
.A2(n_496),
.B(n_477),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_668),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_673),
.B(n_494),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_673),
.B(n_494),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_663),
.A2(n_469),
.B1(n_490),
.B2(n_492),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_694),
.A2(n_588),
.B1(n_625),
.B2(n_579),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_711),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_688),
.A2(n_469),
.B1(n_492),
.B2(n_486),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_714),
.Y(n_748)
);

OAI222xp33_ASAP7_75t_L g749 ( 
.A1(n_702),
.A2(n_477),
.B1(n_496),
.B2(n_567),
.C1(n_566),
.C2(n_460),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_721),
.B(n_495),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_722),
.A2(n_490),
.B1(n_486),
.B2(n_588),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_696),
.A2(n_534),
.B1(n_476),
.B2(n_454),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_702),
.A2(n_476),
.B1(n_454),
.B2(n_474),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_710),
.B(n_495),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_689),
.B(n_488),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_SL g756 ( 
.A1(n_740),
.A2(n_467),
.B(n_677),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_704),
.A2(n_597),
.B1(n_650),
.B2(n_633),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_SL g758 ( 
.A(n_703),
.B(n_460),
.C(n_474),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_697),
.A2(n_454),
.B1(n_475),
.B2(n_456),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_710),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_707),
.B(n_591),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_706),
.A2(n_597),
.B1(n_650),
.B2(n_633),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_723),
.A2(n_454),
.B1(n_475),
.B2(n_456),
.Y(n_763)
);

OAI222xp33_ASAP7_75t_L g764 ( 
.A1(n_723),
.A2(n_578),
.B1(n_574),
.B2(n_557),
.C1(n_554),
.C2(n_449),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_724),
.A2(n_630),
.B1(n_602),
.B2(n_616),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_SL g766 ( 
.A1(n_698),
.A2(n_672),
.B1(n_449),
.B2(n_677),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_717),
.A2(n_602),
.B1(n_616),
.B2(n_630),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_691),
.A2(n_602),
.B1(n_616),
.B2(n_630),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_695),
.A2(n_467),
.B1(n_628),
.B2(n_591),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_693),
.A2(n_467),
.B1(n_628),
.B2(n_633),
.Y(n_770)
);

OAI22xp33_ASAP7_75t_SL g771 ( 
.A1(n_742),
.A2(n_548),
.B1(n_550),
.B2(n_531),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_SL g772 ( 
.A(n_699),
.B(n_467),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_715),
.A2(n_596),
.B1(n_584),
.B2(n_620),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_739),
.A2(n_584),
.B1(n_586),
.B2(n_620),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_720),
.A2(n_500),
.B1(n_626),
.B2(n_618),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_SL g776 ( 
.A1(n_739),
.A2(n_731),
.B1(n_719),
.B2(n_735),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_703),
.A2(n_584),
.B1(n_586),
.B2(n_620),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_730),
.A2(n_584),
.B1(n_586),
.B2(n_620),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_737),
.A2(n_472),
.B1(n_478),
.B2(n_500),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_713),
.A2(n_472),
.B1(n_478),
.B2(n_500),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_690),
.B(n_581),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_732),
.A2(n_584),
.B1(n_586),
.B2(n_620),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_743),
.A2(n_500),
.B1(n_626),
.B2(n_618),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_705),
.A2(n_478),
.B1(n_472),
.B2(n_500),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_690),
.B(n_581),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_727),
.A2(n_500),
.B1(n_626),
.B2(n_618),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_686),
.B(n_626),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_SL g788 ( 
.A1(n_738),
.A2(n_586),
.B1(n_618),
.B2(n_615),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_SL g789 ( 
.A1(n_738),
.A2(n_615),
.B1(n_592),
.B2(n_553),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_718),
.B(n_615),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_SL g791 ( 
.A1(n_718),
.A2(n_615),
.B1(n_592),
.B2(n_553),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_687),
.A2(n_592),
.B1(n_553),
.B2(n_468),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_728),
.A2(n_592),
.B1(n_468),
.B2(n_532),
.Y(n_793)
);

OAI211xp5_ASAP7_75t_SL g794 ( 
.A1(n_726),
.A2(n_488),
.B(n_533),
.C(n_562),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_744),
.A2(n_572),
.B1(n_553),
.B2(n_674),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_725),
.A2(n_517),
.B1(n_674),
.B2(n_269),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_708),
.A2(n_517),
.B1(n_269),
.B2(n_253),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_685),
.A2(n_517),
.B1(n_269),
.B2(n_253),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_SL g799 ( 
.A1(n_776),
.A2(n_692),
.B(n_712),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_748),
.B(n_741),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_755),
.B(n_733),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_748),
.B(n_734),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_746),
.B(n_716),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_760),
.B(n_685),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_790),
.B(n_685),
.Y(n_805)
);

NOR3xp33_ASAP7_75t_L g806 ( 
.A(n_794),
.B(n_700),
.C(n_701),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_790),
.B(n_716),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_745),
.A2(n_729),
.B1(n_736),
.B2(n_716),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_746),
.B(n_716),
.Y(n_809)
);

OAI211xp5_ASAP7_75t_L g810 ( 
.A1(n_758),
.A2(n_701),
.B(n_685),
.C(n_712),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_761),
.B(n_754),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_754),
.B(n_729),
.Y(n_812)
);

NAND4xp25_ASAP7_75t_L g813 ( 
.A(n_781),
.B(n_729),
.C(n_709),
.D(n_107),
.Y(n_813)
);

OAI21xp33_ASAP7_75t_L g814 ( 
.A1(n_766),
.A2(n_104),
.B(n_105),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_787),
.B(n_108),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_792),
.B(n_253),
.C(n_110),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_787),
.B(n_109),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_785),
.B(n_777),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_757),
.B(n_111),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_750),
.B(n_112),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_750),
.B(n_114),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_772),
.A2(n_253),
.B1(n_117),
.B2(n_118),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_771),
.B(n_116),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_763),
.B(n_120),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_779),
.B(n_121),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_791),
.B(n_753),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_759),
.B(n_124),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_756),
.A2(n_253),
.B(n_127),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_765),
.B(n_253),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_783),
.B(n_126),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_SL g831 ( 
.A1(n_764),
.A2(n_130),
.B(n_131),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_811),
.B(n_793),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_800),
.B(n_756),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_800),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_802),
.B(n_789),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_818),
.Y(n_836)
);

AOI221xp5_ASAP7_75t_L g837 ( 
.A1(n_831),
.A2(n_749),
.B1(n_773),
.B2(n_762),
.C(n_751),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_828),
.B(n_778),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_802),
.B(n_786),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_803),
.B(n_775),
.Y(n_840)
);

NOR3xp33_ASAP7_75t_L g841 ( 
.A(n_813),
.B(n_782),
.C(n_788),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_803),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_809),
.B(n_752),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_809),
.B(n_774),
.Y(n_844)
);

NAND3xp33_ASAP7_75t_L g845 ( 
.A(n_823),
.B(n_784),
.C(n_780),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_805),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_818),
.B(n_747),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_804),
.Y(n_848)
);

NAND4xp25_ASAP7_75t_L g849 ( 
.A(n_806),
.B(n_767),
.C(n_769),
.D(n_770),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_807),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_846),
.B(n_812),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_838),
.A2(n_814),
.B1(n_799),
.B2(n_819),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_838),
.A2(n_826),
.B1(n_816),
.B2(n_810),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_834),
.Y(n_854)
);

INVx3_ASAP7_75t_SL g855 ( 
.A(n_838),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_834),
.Y(n_856)
);

CKINVDCx16_ASAP7_75t_R g857 ( 
.A(n_844),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_838),
.A2(n_829),
.B1(n_826),
.B2(n_808),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_836),
.B(n_821),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_848),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_842),
.B(n_801),
.Y(n_861)
);

NOR4xp75_ASAP7_75t_L g862 ( 
.A(n_847),
.B(n_829),
.C(n_815),
.D(n_820),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_842),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_863),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_861),
.Y(n_865)
);

XOR2x2_ASAP7_75t_L g866 ( 
.A(n_852),
.B(n_850),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_860),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_860),
.Y(n_868)
);

XNOR2x1_ASAP7_75t_L g869 ( 
.A(n_851),
.B(n_832),
.Y(n_869)
);

XOR2x2_ASAP7_75t_L g870 ( 
.A(n_855),
.B(n_841),
.Y(n_870)
);

XNOR2xp5_ASAP7_75t_L g871 ( 
.A(n_858),
.B(n_862),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_854),
.Y(n_872)
);

OA22x2_ASAP7_75t_L g873 ( 
.A1(n_871),
.A2(n_855),
.B1(n_865),
.B2(n_868),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_866),
.B(n_857),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_867),
.Y(n_875)
);

OAI22x1_ASAP7_75t_L g876 ( 
.A1(n_867),
.A2(n_859),
.B1(n_856),
.B2(n_835),
.Y(n_876)
);

XOR2x2_ASAP7_75t_L g877 ( 
.A(n_870),
.B(n_853),
.Y(n_877)
);

OA22x2_ASAP7_75t_L g878 ( 
.A1(n_868),
.A2(n_853),
.B1(n_859),
.B2(n_835),
.Y(n_878)
);

AO22x2_ASAP7_75t_L g879 ( 
.A1(n_869),
.A2(n_848),
.B1(n_844),
.B2(n_833),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_872),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_875),
.Y(n_881)
);

OAI22x1_ASAP7_75t_L g882 ( 
.A1(n_874),
.A2(n_872),
.B1(n_864),
.B2(n_833),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_880),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_873),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_878),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_879),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_884),
.A2(n_877),
.B1(n_879),
.B2(n_876),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_881),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_883),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_887),
.A2(n_884),
.B1(n_885),
.B2(n_886),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_888),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_889),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_SL g893 ( 
.A1(n_887),
.A2(n_882),
.B1(n_845),
.B2(n_830),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_891),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_890),
.A2(n_837),
.B1(n_849),
.B2(n_843),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_892),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_893),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_891),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_890),
.A2(n_839),
.B1(n_830),
.B2(n_840),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_898),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_894),
.B(n_840),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_SL g902 ( 
.A1(n_897),
.A2(n_827),
.B1(n_817),
.B2(n_839),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_899),
.B(n_817),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_895),
.A2(n_821),
.B1(n_827),
.B2(n_822),
.Y(n_904)
);

AO22x1_ASAP7_75t_L g905 ( 
.A1(n_896),
.A2(n_824),
.B1(n_825),
.B2(n_795),
.Y(n_905)
);

OR3x2_ASAP7_75t_L g906 ( 
.A(n_900),
.B(n_132),
.C(n_133),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_901),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_903),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_905),
.Y(n_909)
);

NAND4xp75_ASAP7_75t_L g910 ( 
.A(n_904),
.B(n_134),
.C(n_135),
.D(n_136),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_907),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_906),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_908),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_909),
.B(n_902),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_910),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_911),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_913),
.Y(n_917)
);

OA22x2_ASAP7_75t_L g918 ( 
.A1(n_914),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_914),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_912),
.A2(n_772),
.B1(n_768),
.B2(n_796),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_919),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_916),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_917),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_918),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_920),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_918),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_921),
.A2(n_915),
.B1(n_797),
.B2(n_798),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_926),
.A2(n_253),
.B1(n_146),
.B2(n_147),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_927),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_928),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_930),
.A2(n_924),
.B1(n_922),
.B2(n_923),
.Y(n_931)
);

OA22x2_ASAP7_75t_L g932 ( 
.A1(n_929),
.A2(n_924),
.B1(n_925),
.B2(n_149),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_930),
.A2(n_145),
.B1(n_148),
.B2(n_151),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_931),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_932),
.Y(n_935)
);

AOI221x1_ASAP7_75t_L g936 ( 
.A1(n_934),
.A2(n_933),
.B1(n_152),
.B2(n_153),
.C(n_155),
.Y(n_936)
);

AOI211xp5_ASAP7_75t_L g937 ( 
.A1(n_936),
.A2(n_935),
.B(n_156),
.C(n_157),
.Y(n_937)
);


endmodule