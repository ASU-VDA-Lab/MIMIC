module fake_jpeg_1133_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AO22x1_ASAP7_75t_SL g17 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_7),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_2),
.C(n_3),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_20),
.C(n_7),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_21),
.B(n_15),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_10),
.A2(n_0),
.B(n_13),
.Y(n_21)
);

AOI21xp33_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_8),
.B(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_9),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_27),
.Y(n_39)
);

NOR2x1_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_29),
.C(n_34),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_33),
.B1(n_21),
.B2(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_15),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_25),
.B(n_27),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_30),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_18),
.C(n_19),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.C(n_17),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_17),
.C(n_15),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

AOI322xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_32),
.A3(n_35),
.B1(n_37),
.B2(n_38),
.C1(n_39),
.C2(n_42),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_SL g51 ( 
.A1(n_50),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_51)
);


endmodule