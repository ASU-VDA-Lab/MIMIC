module fake_jpeg_11281_n_410 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_410);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_48),
.B(n_58),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_0),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_67),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_18),
.B(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_68),
.B(n_76),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_16),
.Y(n_70)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_77),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_18),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_20),
.B(n_22),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_78),
.Y(n_133)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_81),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_2),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_3),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_85),
.Y(n_128)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_87),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_41),
.B(n_42),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_26),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_89),
.B(n_138),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_71),
.B1(n_86),
.B2(n_75),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_91),
.A2(n_137),
.B1(n_13),
.B2(n_10),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_37),
.B1(n_39),
.B2(n_16),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_95),
.A2(n_106),
.B1(n_121),
.B2(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_105),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_42),
.B1(n_41),
.B2(n_28),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_30),
.B1(n_82),
.B2(n_49),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_43),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_44),
.A2(n_16),
.B1(n_39),
.B2(n_28),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_50),
.A2(n_28),
.B1(n_36),
.B2(n_32),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_109),
.B(n_122),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_40),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_135),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_16),
.B1(n_39),
.B2(n_24),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_72),
.A2(n_39),
.B(n_24),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_60),
.A2(n_39),
.B1(n_24),
.B2(n_36),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_53),
.A2(n_40),
.B1(n_32),
.B2(n_31),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_62),
.B(n_31),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_64),
.A2(n_30),
.B1(n_4),
.B2(n_5),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_65),
.B(n_30),
.C(n_4),
.Y(n_138)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_99),
.B(n_74),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_142),
.B(n_153),
.Y(n_223)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_89),
.A2(n_66),
.B1(n_69),
.B2(n_57),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_146),
.A2(n_148),
.B1(n_174),
.B2(n_180),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_124),
.B(n_82),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_159),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_97),
.A2(n_114),
.B1(n_105),
.B2(n_104),
.Y(n_155)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_187),
.B(n_142),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_91),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_166),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_90),
.B(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_49),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_97),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_97),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_117),
.A2(n_131),
.B(n_135),
.C(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_179),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_167),
.Y(n_227)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_172),
.Y(n_215)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_126),
.B1(n_120),
.B2(n_110),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_93),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_186),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_102),
.A2(n_12),
.B(n_13),
.C(n_108),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_109),
.A2(n_126),
.B1(n_119),
.B2(n_98),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_130),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_125),
.Y(n_193)
);

NAND2x1_ASAP7_75t_SL g185 ( 
.A(n_134),
.B(n_130),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_147),
.B(n_186),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_133),
.Y(n_186)
);

INVx6_ASAP7_75t_SL g187 ( 
.A(n_115),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_125),
.C(n_133),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_226),
.C(n_162),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_193),
.B(n_140),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_194),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_149),
.B(n_139),
.CI(n_115),
.CON(n_197),
.SN(n_197)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_189),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_149),
.A2(n_94),
.B1(n_101),
.B2(n_110),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_203),
.B1(n_208),
.B2(n_211),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_101),
.B1(n_127),
.B2(n_139),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_184),
.A2(n_127),
.B1(n_180),
.B2(n_146),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_206),
.A2(n_218),
.B1(n_212),
.B2(n_189),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_176),
.A2(n_164),
.B1(n_184),
.B2(n_155),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_155),
.A2(n_169),
.B1(n_183),
.B2(n_165),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_155),
.A2(n_183),
.B1(n_142),
.B2(n_175),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_194),
.B1(n_223),
.B2(n_200),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_182),
.B(n_185),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_221),
.B(n_156),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_153),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_147),
.B(n_150),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_143),
.C(n_168),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_206),
.A2(n_178),
.B1(n_151),
.B2(n_144),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_229),
.B(n_252),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_141),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_240),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_232),
.A2(n_204),
.B(n_222),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_233),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_195),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_244),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_209),
.Y(n_283)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_162),
.B1(n_156),
.B2(n_152),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_237),
.A2(n_260),
.B1(n_261),
.B2(n_201),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_171),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_238),
.B(n_262),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_219),
.A2(n_181),
.B1(n_145),
.B2(n_167),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_201),
.B(n_224),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_198),
.A2(n_197),
.B1(n_188),
.B2(n_194),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_243),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_167),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_167),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_215),
.Y(n_244)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_245),
.Y(n_291)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_191),
.B(n_223),
.C(n_194),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_207),
.C(n_216),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_225),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_249),
.Y(n_276)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_225),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_253),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_198),
.A2(n_214),
.B1(n_193),
.B2(n_220),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_221),
.A2(n_219),
.B1(n_212),
.B2(n_203),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_205),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_257),
.Y(n_289)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_199),
.B1(n_190),
.B2(n_192),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_228),
.B1(n_231),
.B2(n_235),
.Y(n_284)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_192),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_232),
.A2(n_217),
.B(n_224),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_263),
.A2(n_268),
.B(n_269),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_273),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_262),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_279),
.Y(n_295)
);

OA22x2_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_222),
.B1(n_207),
.B2(n_216),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_283),
.C(n_242),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_285),
.B1(n_288),
.B2(n_252),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_228),
.A2(n_204),
.B1(n_209),
.B2(n_230),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_240),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_290),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_230),
.A2(n_247),
.B1(n_243),
.B2(n_248),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_259),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_234),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_254),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_294),
.A2(n_317),
.B(n_273),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_303),
.C(n_304),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_309),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_276),
.B1(n_290),
.B2(n_293),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_299),
.A2(n_301),
.B1(n_307),
.B2(n_285),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g300 ( 
.A1(n_280),
.A2(n_251),
.B(n_233),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_300),
.A2(n_316),
.B(n_266),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_289),
.A2(n_230),
.B1(n_257),
.B2(n_255),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_276),
.B(n_244),
.Y(n_302)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_302),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_238),
.C(n_233),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_242),
.C(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_255),
.B1(n_239),
.B2(n_229),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_278),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_284),
.A2(n_246),
.B1(n_250),
.B2(n_256),
.Y(n_310)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_261),
.C(n_260),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_313),
.C(n_277),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_SL g313 ( 
.A(n_280),
.B(n_245),
.C(n_236),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_286),
.B(n_245),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_314),
.B(n_319),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_292),
.Y(n_315)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_279),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_270),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_264),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_318),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_263),
.A2(n_269),
.B(n_282),
.Y(n_319)
);

AOI21xp33_ASAP7_75t_L g348 ( 
.A1(n_321),
.A2(n_298),
.B(n_314),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_277),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_329),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_325),
.A2(n_330),
.B1(n_336),
.B2(n_340),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_303),
.B(n_266),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_326),
.B(n_318),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_277),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_301),
.A2(n_282),
.B1(n_268),
.B2(n_263),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_271),
.C(n_273),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_341),
.C(n_313),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_315),
.Y(n_339)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_299),
.A2(n_273),
.B1(n_275),
.B2(n_274),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_294),
.B(n_302),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_310),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_344),
.Y(n_361)
);

AO21x1_ASAP7_75t_L g345 ( 
.A1(n_330),
.A2(n_305),
.B(n_295),
.Y(n_345)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_295),
.C(n_309),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_350),
.C(n_353),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_348),
.B(n_323),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_316),
.C(n_317),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_327),
.B(n_306),
.Y(n_351)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_351),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_334),
.A2(n_297),
.B(n_305),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_352),
.A2(n_311),
.B(n_319),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_354),
.A2(n_340),
.B1(n_338),
.B2(n_335),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_328),
.A2(n_297),
.B1(n_307),
.B2(n_311),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_357),
.A2(n_325),
.B1(n_336),
.B2(n_328),
.Y(n_369)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_358),
.Y(n_372)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_331),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_333),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_351),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_367),
.Y(n_377)
);

AO21x1_ASAP7_75t_L g364 ( 
.A1(n_357),
.A2(n_345),
.B(n_333),
.Y(n_364)
);

A2O1A1Ixp33_ASAP7_75t_SL g384 ( 
.A1(n_364),
.A2(n_352),
.B(n_342),
.C(n_341),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_369),
.Y(n_379)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_368),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_346),
.B(n_343),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_371),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_329),
.C(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_373),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_355),
.Y(n_374)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_371),
.B(n_356),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_380),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_337),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_349),
.C(n_350),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_382),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_344),
.C(n_356),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_342),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_374),
.B(n_363),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_385),
.B(n_347),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_377),
.A2(n_363),
.B(n_362),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_386),
.A2(n_389),
.B(n_367),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_369),
.C(n_364),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_387),
.B(n_391),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_380),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_362),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_392),
.A2(n_378),
.B1(n_365),
.B2(n_372),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_395),
.B(n_396),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_393),
.A2(n_365),
.B1(n_372),
.B2(n_384),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_397),
.A2(n_399),
.B(n_387),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_392),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_390),
.A2(n_388),
.B(n_389),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_401),
.A2(n_402),
.B(n_403),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_394),
.A2(n_364),
.B(n_384),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_400),
.B(n_347),
.C(n_395),
.Y(n_404)
);

O2A1O1Ixp33_ASAP7_75t_SL g406 ( 
.A1(n_404),
.A2(n_353),
.B(n_326),
.C(n_273),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_405),
.B1(n_291),
.B2(n_274),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_407),
.A2(n_272),
.B(n_265),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_272),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_265),
.Y(n_410)
);


endmodule