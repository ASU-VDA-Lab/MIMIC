module fake_jpeg_2448_n_122 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_122);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx8_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_11),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_21),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_31),
.B1(n_12),
.B2(n_13),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_34),
.B1(n_36),
.B2(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_63),
.Y(n_70)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_56),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_60),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_73),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_61),
.B1(n_39),
.B2(n_3),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_29),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_59),
.B1(n_39),
.B2(n_35),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_0),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_61),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_81),
.C(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_84),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_14),
.C(n_28),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_87),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_100),
.C(n_6),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_64),
.C(n_69),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_96),
.C(n_19),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_2),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_101),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_109),
.B1(n_9),
.B2(n_10),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_107),
.C(n_95),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_89),
.B1(n_93),
.B2(n_11),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_114),
.C(n_104),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_108),
.A2(n_92),
.B(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_113),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_115),
.B1(n_102),
.B2(n_112),
.Y(n_119)
);

OAI321xp33_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_110),
.A3(n_103),
.B1(n_105),
.B2(n_10),
.C(n_15),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_17),
.B(n_18),
.Y(n_121)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_121),
.Y(n_122)
);


endmodule