module fake_aes_5946_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_9), .B(n_4), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_3), .B(n_8), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_13), .B(n_0), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_0), .B(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_14), .B(n_1), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
OAI21x1_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_11), .B(n_15), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_20), .B(n_17), .Y(n_23) );
OAI33xp33_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_16), .A3(n_13), .B1(n_11), .B2(n_20), .B3(n_21), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_22), .B(n_20), .Y(n_25) );
OAI222xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_16), .B1(n_12), .B2(n_24), .C1(n_5), .C2(n_6), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_12), .B1(n_3), .B2(n_4), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
AOI211xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_2), .B(n_5), .C(n_6), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
INVx5_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_28), .B(n_10), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_7), .B1(n_9), .B2(n_10), .Y(n_33) );
INVx4_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
CKINVDCx20_ASAP7_75t_R g35 ( .A(n_34), .Y(n_35) );
OAI221xp5_ASAP7_75t_R g36 ( .A1(n_35), .A2(n_31), .B1(n_33), .B2(n_27), .C(n_34), .Y(n_36) );
endmodule