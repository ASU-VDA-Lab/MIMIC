module fake_jpeg_12337_n_668 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_668);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_668;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_60),
.B(n_70),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_62),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g65 ( 
.A1(n_30),
.A2(n_19),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_65),
.B(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_67),
.Y(n_175)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_68),
.Y(n_220)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_69),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_73),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g193 ( 
.A(n_77),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_79),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_81),
.B(n_84),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_19),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_85),
.B(n_90),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_86),
.Y(n_208)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_89),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_39),
.B(n_18),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_91),
.B(n_97),
.Y(n_182)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_92),
.Y(n_159)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_94),
.Y(n_217)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g170 ( 
.A(n_96),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_17),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_99),
.B(n_100),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_43),
.B(n_17),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_26),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_101),
.B(n_105),
.Y(n_209)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_43),
.B(n_16),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_119),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_35),
.Y(n_108)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_112),
.Y(n_214)
);

BUFx24_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_115),
.Y(n_199)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_35),
.Y(n_117)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_26),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_15),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_26),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_122),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_35),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_125),
.B(n_130),
.Y(n_203)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_21),
.Y(n_129)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_59),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_21),
.Y(n_131)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_21),
.B1(n_27),
.B2(n_55),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_136),
.A2(n_181),
.B1(n_195),
.B2(n_46),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_57),
.B(n_46),
.C(n_45),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_139),
.A2(n_189),
.B(n_72),
.Y(n_238)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_21),
.C(n_27),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_140),
.B(n_25),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_23),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_162),
.B(n_183),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_77),
.A2(n_23),
.B(n_56),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_165),
.B(n_194),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_27),
.B1(n_56),
.B2(n_55),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_176),
.A2(n_223),
.B1(n_9),
.B2(n_10),
.Y(n_283)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_63),
.A2(n_27),
.B1(n_80),
.B2(n_124),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_99),
.B(n_20),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_108),
.B(n_20),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_185),
.B(n_224),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_77),
.A2(n_40),
.B(n_49),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_71),
.Y(n_190)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_96),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_74),
.A2(n_22),
.B1(n_53),
.B2(n_52),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_82),
.Y(n_196)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_196),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_127),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_197),
.B(n_106),
.Y(n_245)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_69),
.Y(n_200)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_200),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_SL g201 ( 
.A1(n_78),
.A2(n_44),
.B(n_53),
.Y(n_201)
);

NAND2xp67_ASAP7_75t_SL g260 ( 
.A(n_201),
.B(n_139),
.Y(n_260)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_92),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_202),
.Y(n_293)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_215),
.Y(n_232)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_94),
.Y(n_206)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

BUFx4f_ASAP7_75t_L g210 ( 
.A(n_95),
.Y(n_210)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_98),
.Y(n_212)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_104),
.Y(n_213)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_213),
.Y(n_272)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_103),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_117),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_112),
.Y(n_222)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_222),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_114),
.A2(n_44),
.B1(n_57),
.B2(n_36),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_115),
.B(n_40),
.Y(n_224)
);

INVx11_ASAP7_75t_L g225 ( 
.A(n_73),
.Y(n_225)
);

INVx11_ASAP7_75t_L g308 ( 
.A(n_225),
.Y(n_308)
);

CKINVDCx12_ASAP7_75t_R g227 ( 
.A(n_170),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_227),
.Y(n_337)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_141),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_228),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_230),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_174),
.Y(n_230)
);

OA22x2_ASAP7_75t_SL g233 ( 
.A1(n_201),
.A2(n_64),
.B1(n_72),
.B2(n_44),
.Y(n_233)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_233),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_174),
.B(n_64),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_237),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_238),
.B(n_249),
.Y(n_317)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_141),
.Y(n_239)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_239),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_132),
.B(n_67),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_240),
.B(n_306),
.C(n_186),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_135),
.A2(n_36),
.B(n_37),
.C(n_45),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_241),
.B(n_292),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_148),
.B(n_37),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_242),
.B(n_261),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_243),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_209),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_245),
.Y(n_313)
);

CKINVDCx12_ASAP7_75t_R g246 ( 
.A(n_161),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_246),
.Y(n_310)
);

HAxp5_ASAP7_75t_SL g248 ( 
.A(n_189),
.B(n_79),
.CON(n_248),
.SN(n_248)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_178),
.A2(n_68),
.B1(n_62),
.B2(n_52),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_251),
.A2(n_274),
.B1(n_275),
.B2(n_291),
.Y(n_335)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_144),
.Y(n_253)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_253),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_209),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_254),
.B(n_276),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_155),
.A2(n_128),
.B1(n_49),
.B2(n_25),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_255),
.A2(n_283),
.B1(n_273),
.B2(n_264),
.Y(n_364)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_144),
.Y(n_256)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_256),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_258),
.B(n_260),
.Y(n_343)
);

CKINVDCx12_ASAP7_75t_R g259 ( 
.A(n_160),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_259),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_172),
.B(n_22),
.Y(n_261)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_146),
.Y(n_262)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_262),
.Y(n_339)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_146),
.Y(n_264)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_264),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_265),
.A2(n_266),
.B1(n_282),
.B2(n_239),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_177),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_266)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_149),
.Y(n_268)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_268),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_137),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_270),
.Y(n_323)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_210),
.Y(n_271)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_271),
.Y(n_325)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_149),
.Y(n_273)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_273),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_178),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_193),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_203),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_172),
.B(n_15),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_277),
.B(n_281),
.Y(n_348)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_137),
.Y(n_278)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_278),
.Y(n_351)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_156),
.Y(n_280)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_280),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_138),
.B(n_6),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_133),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_156),
.Y(n_285)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_285),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_188),
.B(n_10),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_286),
.B(n_290),
.Y(n_353)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_142),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_289),
.Y(n_334)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_142),
.Y(n_288)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_288),
.Y(n_369)
);

BUFx12f_ASAP7_75t_L g289 ( 
.A(n_219),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_188),
.B(n_10),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_191),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_167),
.B(n_12),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_193),
.A2(n_13),
.B1(n_151),
.B2(n_171),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_295),
.A2(n_303),
.B1(n_304),
.B2(n_186),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_167),
.B(n_182),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_297),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_191),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_299),
.Y(n_352)
);

BUFx4f_ASAP7_75t_SL g299 ( 
.A(n_168),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_182),
.B(n_143),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_300),
.B(n_301),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_153),
.B(n_134),
.Y(n_301)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_208),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_305),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_175),
.A2(n_150),
.B1(n_159),
.B2(n_163),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_150),
.A2(n_159),
.B1(n_220),
.B2(n_140),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_179),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_154),
.B(n_164),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_186),
.B(n_152),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_307),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_236),
.A2(n_166),
.B(n_223),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_309),
.A2(n_356),
.B(n_267),
.Y(n_403)
);

OA22x2_ASAP7_75t_L g314 ( 
.A1(n_260),
.A2(n_214),
.B1(n_177),
.B2(n_157),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_320),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_249),
.A2(n_214),
.B1(n_211),
.B2(n_145),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_315),
.A2(n_326),
.B1(n_365),
.B2(n_271),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_319),
.A2(n_328),
.B1(n_329),
.B2(n_361),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_279),
.B(n_145),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_269),
.B(n_169),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_324),
.B(n_338),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_238),
.A2(n_169),
.B1(n_226),
.B2(n_217),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_282),
.A2(n_217),
.B1(n_216),
.B2(n_199),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_248),
.A2(n_216),
.B1(n_187),
.B2(n_158),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_237),
.A2(n_233),
.B(n_240),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_332),
.A2(n_356),
.B(n_321),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_241),
.B(n_147),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_237),
.B(n_207),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_350),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_341),
.Y(n_402)
);

NOR3xp33_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_308),
.C(n_299),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_240),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_306),
.B(n_294),
.C(n_232),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_354),
.B(n_297),
.C(n_298),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_235),
.B(n_305),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_366),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_233),
.A2(n_270),
.B(n_293),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_228),
.A2(n_280),
.B1(n_302),
.B2(n_268),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_364),
.B(n_285),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_250),
.A2(n_257),
.B1(n_252),
.B2(n_234),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_293),
.B(n_247),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_231),
.B(n_272),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_267),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_231),
.A2(n_284),
.B1(n_234),
.B2(n_263),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_368),
.A2(n_272),
.B1(n_263),
.B2(n_262),
.Y(n_396)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_360),
.Y(n_370)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_370),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_372),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_373),
.A2(n_403),
.B(n_416),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_243),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_374),
.B(n_378),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_308),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_375),
.B(n_382),
.Y(n_433)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_367),
.Y(n_376)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_334),
.Y(n_377)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_377),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_318),
.B(n_253),
.Y(n_378)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_381),
.Y(n_422)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_343),
.B(n_299),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_365),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_383),
.B(n_386),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_357),
.B(n_284),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_384),
.B(n_385),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_256),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_311),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_366),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_400),
.Y(n_425)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_333),
.Y(n_388)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_388),
.Y(n_430)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_390),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_323),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_391),
.Y(n_438)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_393),
.Y(n_444)
);

INVx13_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

BUFx8_ASAP7_75t_L g445 ( 
.A(n_394),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

INVx11_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_397),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_313),
.B(n_288),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_398),
.Y(n_432)
);

AOI21xp33_ASAP7_75t_L g399 ( 
.A1(n_321),
.A2(n_229),
.B(n_289),
.Y(n_399)
);

FAx1_ASAP7_75t_SL g423 ( 
.A(n_399),
.B(n_341),
.CI(n_340),
.CON(n_423),
.SN(n_423)
);

INVx13_ASAP7_75t_L g400 ( 
.A(n_310),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_404),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_355),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_407),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_406),
.A2(n_412),
.B1(n_361),
.B2(n_328),
.Y(n_418)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_325),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_324),
.B(n_278),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_408),
.B(n_409),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_330),
.B(n_287),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_312),
.B(n_287),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_410),
.B(n_343),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_411),
.A2(n_364),
.B1(n_335),
.B2(n_347),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_336),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_320),
.B(n_291),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_415),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_414),
.B(n_329),
.C(n_314),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g415 ( 
.A(n_348),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_332),
.A2(n_289),
.B(n_317),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_338),
.B(n_316),
.Y(n_417)
);

AO22x1_ASAP7_75t_L g431 ( 
.A1(n_417),
.A2(n_403),
.B1(n_309),
.B2(n_316),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_418),
.B(n_380),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_421),
.B(n_429),
.C(n_437),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_423),
.A2(n_453),
.B(n_429),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_322),
.C(n_354),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_431),
.B(n_389),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_373),
.Y(n_460)
);

OAI32xp33_ASAP7_75t_L g436 ( 
.A1(n_379),
.A2(n_342),
.A3(n_350),
.B1(n_317),
.B2(n_346),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_448),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_379),
.B(n_317),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_371),
.A2(n_319),
.B1(n_322),
.B2(n_342),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_439),
.A2(n_442),
.B1(n_450),
.B2(n_454),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_371),
.A2(n_376),
.B1(n_387),
.B2(n_405),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_383),
.A2(n_314),
.B1(n_368),
.B2(n_347),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_402),
.B(n_314),
.C(n_353),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_414),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_408),
.A2(n_359),
.B1(n_339),
.B2(n_363),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_417),
.A2(n_352),
.B1(n_363),
.B2(n_359),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_455),
.B(n_456),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_417),
.A2(n_336),
.B1(n_344),
.B2(n_333),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_391),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_459),
.A2(n_476),
.B(n_426),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_460),
.B(n_448),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_382),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_462),
.B(n_475),
.Y(n_497)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_425),
.Y(n_463)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_463),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_457),
.B(n_384),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_465),
.B(n_472),
.Y(n_509)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_425),
.Y(n_466)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_466),
.Y(n_506)
);

O2A1O1Ixp33_ASAP7_75t_L g467 ( 
.A1(n_431),
.A2(n_397),
.B(n_416),
.C(n_375),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_467),
.A2(n_487),
.B(n_490),
.Y(n_502)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_427),
.Y(n_468)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_434),
.B(n_413),
.Y(n_469)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_469),
.Y(n_517)
);

XNOR2x1_ASAP7_75t_L g516 ( 
.A(n_470),
.B(n_423),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_427),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_434),
.Y(n_473)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_473),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_392),
.Y(n_474)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_474),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_447),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_491),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_432),
.B(n_428),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_478),
.B(n_481),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_438),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_479),
.B(n_484),
.Y(n_519)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_422),
.Y(n_480)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_480),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_390),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_310),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_482),
.B(n_483),
.Y(n_504)
);

FAx1_ASAP7_75t_SL g483 ( 
.A(n_437),
.B(n_389),
.CI(n_392),
.CON(n_483),
.SN(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_451),
.B(n_407),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_445),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_485),
.B(n_486),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_452),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_447),
.A2(n_404),
.B(n_411),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_435),
.B(n_401),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_488),
.B(n_423),
.C(n_420),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_452),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_489),
.B(n_422),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_443),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_455),
.B(n_381),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_492),
.B(n_494),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_424),
.B(n_380),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_493),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_370),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_477),
.A2(n_420),
.B(n_421),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_495),
.A2(n_490),
.B(n_487),
.Y(n_531)
);

INVxp33_ASAP7_75t_SL g496 ( 
.A(n_461),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_496),
.B(n_512),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_458),
.A2(n_466),
.B1(n_463),
.B2(n_473),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_499),
.A2(n_461),
.B1(n_464),
.B2(n_507),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_486),
.B(n_439),
.Y(n_505)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_505),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_491),
.B(n_436),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_L g532 ( 
.A(n_508),
.B(n_468),
.Y(n_532)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_510),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_451),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_472),
.B(n_454),
.Y(n_513)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_513),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_459),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_514),
.B(n_521),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_515),
.B(n_525),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_516),
.B(n_528),
.C(n_529),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_474),
.B(n_449),
.Y(n_518)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_518),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_459),
.B(n_431),
.Y(n_520)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_520),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_351),
.Y(n_521)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_523),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_469),
.B(n_449),
.Y(n_526)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_526),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_471),
.B(n_430),
.C(n_351),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_471),
.B(n_450),
.C(n_369),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_531),
.A2(n_497),
.B(n_509),
.Y(n_577)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_532),
.Y(n_564)
);

BUFx5_ASAP7_75t_L g533 ( 
.A(n_530),
.Y(n_533)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_533),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_534),
.A2(n_545),
.B1(n_557),
.B2(n_558),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_500),
.B(n_467),
.Y(n_541)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_528),
.B(n_470),
.C(n_488),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_543),
.B(n_551),
.C(n_502),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_500),
.Y(n_544)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_544),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_499),
.A2(n_475),
.B1(n_458),
.B2(n_493),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_529),
.B(n_476),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_546),
.B(n_550),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_498),
.B(n_483),
.Y(n_548)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_548),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_498),
.B(n_479),
.Y(n_549)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_549),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_516),
.B(n_464),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_495),
.B(n_492),
.C(n_493),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_505),
.A2(n_494),
.B1(n_418),
.B2(n_475),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_552),
.A2(n_560),
.B1(n_561),
.B2(n_503),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_508),
.A2(n_426),
.B1(n_462),
.B2(n_480),
.Y(n_555)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_555),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_515),
.A2(n_485),
.B1(n_406),
.B2(n_446),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_525),
.A2(n_444),
.B1(n_412),
.B2(n_395),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_502),
.B(n_400),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_559),
.B(n_558),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_523),
.A2(n_412),
.B1(n_395),
.B2(n_396),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_523),
.A2(n_388),
.B1(n_393),
.B2(n_344),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_562),
.B(n_577),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_543),
.B(n_497),
.C(n_501),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_565),
.B(n_583),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_553),
.B(n_514),
.Y(n_566)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_566),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_538),
.B(n_504),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_569),
.B(n_571),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_535),
.B(n_504),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_SL g594 ( 
.A(n_572),
.B(n_579),
.Y(n_594)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_533),
.Y(n_574)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_574),
.Y(n_590)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_554),
.Y(n_575)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_575),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_544),
.B(n_509),
.Y(n_576)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_576),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_556),
.A2(n_527),
.B1(n_517),
.B2(n_522),
.Y(n_578)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_578),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_547),
.B(n_520),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_581),
.A2(n_582),
.B1(n_534),
.B2(n_539),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_552),
.A2(n_503),
.B1(n_506),
.B2(n_501),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_542),
.B(n_527),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_537),
.B(n_506),
.C(n_522),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_585),
.B(n_524),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_565),
.B(n_559),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_589),
.B(n_567),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_585),
.B(n_537),
.C(n_546),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_595),
.B(n_599),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_570),
.B(n_519),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_597),
.B(n_575),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_SL g598 ( 
.A(n_579),
.B(n_547),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_598),
.B(n_601),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_562),
.B(n_551),
.C(n_550),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_SL g600 ( 
.A(n_577),
.B(n_541),
.C(n_524),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_600),
.A2(n_581),
.B(n_507),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_SL g601 ( 
.A(n_567),
.B(n_545),
.Y(n_601)
);

OA21x2_ASAP7_75t_L g602 ( 
.A1(n_566),
.A2(n_561),
.B(n_560),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_602),
.A2(n_603),
.B1(n_580),
.B2(n_572),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_564),
.B(n_519),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_604),
.B(n_606),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_573),
.A2(n_536),
.B(n_540),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_607),
.A2(n_518),
.B(n_526),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_600),
.A2(n_573),
.B(n_584),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_608),
.A2(n_612),
.B(n_614),
.Y(n_631)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_590),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_609),
.B(n_615),
.Y(n_630)
);

INVx11_ASAP7_75t_L g611 ( 
.A(n_607),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_611),
.A2(n_602),
.B1(n_513),
.B2(n_511),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_588),
.A2(n_576),
.B(n_568),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_605),
.A2(n_582),
.B(n_583),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_616),
.B(n_594),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_617),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_602),
.A2(n_603),
.B1(n_580),
.B2(n_596),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_618),
.A2(n_511),
.B1(n_563),
.B2(n_601),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g619 ( 
.A1(n_587),
.A2(n_586),
.B(n_557),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_619),
.B(n_530),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_593),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_620),
.B(n_621),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_SL g634 ( 
.A1(n_623),
.A2(n_563),
.B(n_599),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_592),
.B(n_574),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_624),
.B(n_625),
.Y(n_639)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_591),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_611),
.B(n_517),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_626),
.B(n_628),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_610),
.B(n_595),
.C(n_593),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_616),
.B(n_589),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_629),
.Y(n_642)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_633),
.Y(n_648)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_634),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_635),
.A2(n_615),
.B1(n_622),
.B2(n_614),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_636),
.A2(n_637),
.B(n_612),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_617),
.B(n_594),
.C(n_598),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_638),
.B(n_608),
.C(n_622),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_641),
.B(n_647),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_643),
.B(n_644),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_628),
.B(n_639),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_632),
.B(n_613),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_645),
.B(n_646),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_636),
.B(n_618),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_631),
.A2(n_400),
.B(n_445),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g652 ( 
.A(n_649),
.B(n_627),
.Y(n_652)
);

AOI322xp5_ASAP7_75t_L g651 ( 
.A1(n_650),
.A2(n_627),
.A3(n_630),
.B1(n_638),
.B2(n_637),
.C1(n_629),
.C2(n_394),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_651),
.B(n_657),
.Y(n_660)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_652),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_SL g654 ( 
.A1(n_640),
.A2(n_445),
.B(n_394),
.C(n_369),
.Y(n_654)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_654),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_642),
.B(n_331),
.C(n_327),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_653),
.B(n_648),
.Y(n_659)
);

AOI31xp33_ASAP7_75t_L g663 ( 
.A1(n_659),
.A2(n_642),
.A3(n_655),
.B(n_641),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_660),
.B(n_656),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_SL g664 ( 
.A(n_662),
.B(n_663),
.C(n_658),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_664),
.B(n_661),
.C(n_654),
.Y(n_665)
);

XNOR2xp5_ASAP7_75t_L g666 ( 
.A(n_665),
.B(n_649),
.Y(n_666)
);

XOR2xp5_ASAP7_75t_L g667 ( 
.A(n_666),
.B(n_327),
.Y(n_667)
);

OAI31xp33_ASAP7_75t_L g668 ( 
.A1(n_667),
.A2(n_331),
.A3(n_349),
.B(n_611),
.Y(n_668)
);


endmodule