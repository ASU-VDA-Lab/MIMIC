module fake_ibex_1307_n_959 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_959);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_959;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_457;
wire n_357;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_170;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_791;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_354;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_444;
wire n_200;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_927;
wire n_684;
wire n_775;
wire n_784;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g168 ( 
.A(n_64),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_47),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_3),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_31),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_19),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g177 ( 
.A(n_24),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_44),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_55),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_72),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_119),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_80),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_67),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_76),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_88),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_65),
.B(n_101),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_103),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_54),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_71),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_118),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_75),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_1),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_57),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_63),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_89),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_33),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_36),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_17),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_91),
.B(n_56),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_133),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_115),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_35),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_10),
.B(n_92),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_126),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_69),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_70),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_129),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_49),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_107),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_105),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_41),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_66),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_51),
.B(n_167),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_98),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_125),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_138),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_149),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_30),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_40),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_94),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_62),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_46),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_74),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_132),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_15),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_68),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_131),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_109),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_0),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_21),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g249 ( 
.A(n_102),
.B(n_137),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_35),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_22),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_117),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_90),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_31),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_22),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_160),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_7),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_15),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_112),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_39),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_29),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_33),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_93),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_27),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_61),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_163),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_20),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_113),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_9),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_106),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_108),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_59),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_140),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_77),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_78),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_25),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_162),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_144),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_12),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_20),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_147),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_158),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_10),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_172),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_173),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_172),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_211),
.B(n_2),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_4),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_211),
.B(n_5),
.Y(n_292)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_190),
.B(n_42),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_185),
.B(n_5),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_251),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_202),
.A2(n_257),
.B1(n_214),
.B2(n_248),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_179),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_170),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_205),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_172),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_170),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_192),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_179),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_236),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_170),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_172),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g311 ( 
.A1(n_168),
.A2(n_83),
.B(n_165),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_170),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_6),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_187),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_176),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_170),
.B(n_6),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_170),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_243),
.Y(n_320)
);

NOR2x1_ASAP7_75t_L g321 ( 
.A(n_198),
.B(n_43),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_192),
.B(n_7),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_218),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_202),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_197),
.B(n_8),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_258),
.B(n_8),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

OAI22x1_ASAP7_75t_SL g329 ( 
.A1(n_257),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_269),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_218),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_218),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_187),
.Y(n_334)
);

BUFx8_ASAP7_75t_SL g335 ( 
.A(n_175),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_218),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_280),
.Y(n_337)
);

CKINVDCx6p67_ASAP7_75t_R g338 ( 
.A(n_197),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_218),
.Y(n_339)
);

OAI21x1_ASAP7_75t_L g340 ( 
.A1(n_224),
.A2(n_237),
.B(n_231),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_218),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_177),
.B(n_14),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_238),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_177),
.A2(n_174),
.B1(n_247),
.B2(n_207),
.Y(n_344)
);

CKINVDCx6p67_ASAP7_75t_R g345 ( 
.A(n_206),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_242),
.B(n_16),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_187),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_171),
.B(n_17),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_180),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_245),
.B(n_265),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_245),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_265),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_222),
.B(n_18),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_187),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_188),
.B(n_18),
.Y(n_355)
);

INVx6_ASAP7_75t_L g356 ( 
.A(n_209),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_287),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_350),
.Y(n_359)
);

OR2x6_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_217),
.Y(n_360)
);

OR2x6_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_243),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_191),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_325),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_355),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_350),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_355),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_289),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_296),
.Y(n_370)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_322),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_306),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_289),
.Y(n_373)
);

NAND2xp33_ASAP7_75t_R g374 ( 
.A(n_303),
.B(n_250),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_299),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_R g377 ( 
.A(n_303),
.B(n_254),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_317),
.A2(n_283),
.B1(n_243),
.B2(n_204),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_264),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_322),
.B(n_189),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_291),
.B(n_314),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_291),
.B(n_267),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_326),
.B(n_194),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_323),
.A2(n_283),
.B1(n_282),
.B2(n_210),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_290),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_326),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_295),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_295),
.Y(n_389)
);

INVxp33_ASAP7_75t_SL g390 ( 
.A(n_353),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_328),
.A2(n_283),
.B1(n_215),
.B2(n_278),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_343),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_335),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_300),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_307),
.B(n_199),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_314),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_300),
.B(n_200),
.Y(n_400)
);

AND2x6_ASAP7_75t_L g401 ( 
.A(n_293),
.B(n_203),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_305),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_331),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_306),
.Y(n_404)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_311),
.A2(n_219),
.B(n_216),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_305),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_325),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_338),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_307),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_288),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_318),
.A2(n_283),
.B1(n_233),
.B2(n_277),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_309),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_309),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

BUFx10_ASAP7_75t_L g417 ( 
.A(n_292),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_345),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_301),
.Y(n_419)
);

AND3x2_ASAP7_75t_L g420 ( 
.A(n_329),
.B(n_223),
.C(n_221),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_304),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_308),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_312),
.Y(n_423)
);

BUFx4f_ASAP7_75t_L g424 ( 
.A(n_311),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_313),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_352),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_313),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_319),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_324),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_335),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_324),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_332),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_316),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_L g435 ( 
.A(n_333),
.B(n_208),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_333),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_336),
.B(n_225),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_351),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_339),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_339),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g441 ( 
.A(n_321),
.B(n_230),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_341),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_286),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_294),
.B(n_181),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_327),
.B(n_182),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_348),
.Y(n_446)
);

AOI21x1_ASAP7_75t_L g447 ( 
.A1(n_311),
.A2(n_235),
.B(n_232),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_316),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_346),
.B(n_183),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_315),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_315),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_297),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_344),
.B(n_241),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_347),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_359),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_394),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_361),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_408),
.B(n_184),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_381),
.B(n_412),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_193),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_408),
.B(n_195),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_196),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_363),
.A2(n_285),
.B1(n_239),
.B2(n_186),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_404),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_359),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_361),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_360),
.B(n_330),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_399),
.B(n_201),
.Y(n_469)
);

O2A1O1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_363),
.A2(n_259),
.B(n_270),
.C(n_266),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_361),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_409),
.B(n_226),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_382),
.B(n_178),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_409),
.B(n_212),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

A2O1A1Ixp33_ASAP7_75t_L g476 ( 
.A1(n_362),
.A2(n_367),
.B(n_365),
.C(n_383),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_418),
.B(n_220),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_416),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_403),
.B(n_227),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_372),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_390),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_398),
.B(n_271),
.Y(n_482)
);

NOR3xp33_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_274),
.C(n_273),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_387),
.A2(n_315),
.B1(n_320),
.B2(n_209),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_360),
.B(n_213),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_366),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_410),
.B(n_229),
.Y(n_487)
);

O2A1O1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_453),
.A2(n_320),
.B(n_228),
.C(n_249),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_430),
.Y(n_489)
);

AOI221xp5_ASAP7_75t_L g490 ( 
.A1(n_419),
.A2(n_422),
.B1(n_423),
.B2(n_421),
.C(n_398),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_360),
.A2(n_263),
.B1(n_240),
.B2(n_244),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_366),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_444),
.B(n_246),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_396),
.A2(n_320),
.B1(n_209),
.B2(n_356),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_379),
.B(n_252),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_426),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_374),
.A2(n_272),
.B1(n_275),
.B2(n_253),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_397),
.A2(n_368),
.B1(n_401),
.B2(n_441),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_376),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_417),
.B(n_256),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_368),
.A2(n_209),
.B1(n_356),
.B2(n_347),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_377),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_426),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_411),
.B(n_169),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_424),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_392),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_401),
.A2(n_441),
.B1(n_435),
.B2(n_384),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_405),
.A2(n_228),
.B(n_316),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_377),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_417),
.B(n_260),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_449),
.B(n_268),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_380),
.B(n_281),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_R g514 ( 
.A(n_364),
.B(n_45),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_393),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_371),
.B(n_370),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_371),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_401),
.A2(n_356),
.B1(n_354),
.B2(n_347),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_438),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_375),
.B(n_48),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_400),
.B(n_354),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_441),
.B(n_284),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_441),
.B(n_284),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_437),
.B(n_284),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_395),
.Y(n_525)
);

OAI221xp5_ASAP7_75t_L g526 ( 
.A1(n_385),
.A2(n_334),
.B1(n_310),
.B2(n_302),
.C(n_25),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_L g527 ( 
.A(n_452),
.B(n_21),
.C(n_23),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_401),
.A2(n_415),
.B1(n_402),
.B2(n_406),
.Y(n_528)
);

OAI221xp5_ASAP7_75t_L g529 ( 
.A1(n_385),
.A2(n_334),
.B1(n_310),
.B2(n_302),
.C(n_27),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_391),
.B(n_302),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_391),
.B(n_428),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_413),
.B(n_24),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_429),
.Y(n_533)
);

BUFx6f_ASAP7_75t_SL g534 ( 
.A(n_420),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_457),
.B(n_432),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_460),
.B(n_433),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_490),
.B(n_439),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_485),
.B(n_475),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_483),
.B(n_440),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_475),
.A2(n_427),
.B1(n_414),
.B2(n_415),
.Y(n_541)
);

NAND2x1_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_425),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_508),
.A2(n_427),
.B1(n_431),
.B2(n_436),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_483),
.B(n_431),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_476),
.A2(n_509),
.B(n_516),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_489),
.Y(n_546)
);

AO21x1_ASAP7_75t_L g547 ( 
.A1(n_488),
.A2(n_447),
.B(n_442),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_525),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_472),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_466),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_467),
.A2(n_378),
.B1(n_389),
.B2(n_388),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_486),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_482),
.B(n_358),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_464),
.B(n_26),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_481),
.B(n_364),
.Y(n_556)
);

NOR2x1p5_ASAP7_75t_L g557 ( 
.A(n_456),
.B(n_407),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_508),
.A2(n_378),
.B1(n_386),
.B2(n_358),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_479),
.A2(n_487),
.B(n_495),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_481),
.B(n_407),
.Y(n_560)
);

BUFx4f_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_492),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_532),
.A2(n_389),
.B1(n_369),
.B2(n_373),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_507),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_471),
.A2(n_451),
.B1(n_450),
.B2(n_448),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_517),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_510),
.B(n_26),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_510),
.B(n_28),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_515),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_463),
.A2(n_454),
.B(n_443),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_482),
.B(n_434),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_498),
.B(n_302),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_468),
.B(n_28),
.Y(n_573)
);

CKINVDCx8_ASAP7_75t_R g574 ( 
.A(n_505),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_531),
.A2(n_334),
.B(n_310),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_528),
.B(n_310),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_511),
.B(n_334),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_473),
.B(n_29),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_461),
.B(n_357),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_493),
.B(n_512),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_502),
.A2(n_357),
.B1(n_30),
.B2(n_32),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_493),
.B(n_32),
.Y(n_582)
);

O2A1O1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_469),
.A2(n_34),
.B(n_36),
.C(n_37),
.Y(n_583)
);

BUFx8_ASAP7_75t_L g584 ( 
.A(n_534),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_534),
.B(n_37),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_503),
.B(n_50),
.Y(n_586)
);

INVx11_ASAP7_75t_L g587 ( 
.A(n_514),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_504),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_491),
.A2(n_38),
.B1(n_52),
.B2(n_53),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_497),
.Y(n_590)
);

AO21x1_ASAP7_75t_L g591 ( 
.A1(n_520),
.A2(n_38),
.B(n_58),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_499),
.B(n_60),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_519),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_458),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_465),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_512),
.B(n_513),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_459),
.B(n_166),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_462),
.B(n_73),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_478),
.Y(n_599)
);

INVx11_ASAP7_75t_L g600 ( 
.A(n_477),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_530),
.A2(n_524),
.B(n_522),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_484),
.A2(n_506),
.B1(n_503),
.B2(n_494),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_500),
.B(n_79),
.Y(n_603)
);

O2A1O1Ixp33_ASAP7_75t_SL g604 ( 
.A1(n_523),
.A2(n_81),
.B(n_82),
.C(n_84),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_480),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_503),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g607 ( 
.A(n_527),
.B(n_95),
.C(n_96),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_484),
.A2(n_97),
.B1(n_100),
.B2(n_104),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_496),
.Y(n_609)
);

AO21x1_ASAP7_75t_L g610 ( 
.A1(n_524),
.A2(n_121),
.B(n_122),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_539),
.B(n_474),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_593),
.B(n_506),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_554),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_559),
.A2(n_506),
.B(n_521),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_548),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_575),
.A2(n_494),
.B(n_521),
.Y(n_616)
);

A2O1A1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_580),
.A2(n_529),
.B(n_526),
.C(n_518),
.Y(n_617)
);

OAI21xp33_ASAP7_75t_SL g618 ( 
.A1(n_553),
.A2(n_518),
.B(n_501),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_542),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_556),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_566),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_601),
.A2(n_128),
.B(n_130),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_SL g623 ( 
.A1(n_563),
.A2(n_161),
.B(n_139),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_540),
.B(n_134),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_537),
.B(n_145),
.Y(n_625)
);

A2O1A1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_596),
.A2(n_146),
.B(n_150),
.C(n_151),
.Y(n_626)
);

INVxp33_ASAP7_75t_L g627 ( 
.A(n_560),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_538),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_550),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_575),
.A2(n_152),
.B(n_156),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_549),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_590),
.B(n_574),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_566),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_597),
.B(n_598),
.Y(n_634)
);

AOI21xp33_ASAP7_75t_L g635 ( 
.A1(n_578),
.A2(n_544),
.B(n_582),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_594),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_SL g637 ( 
.A(n_546),
.B(n_587),
.Y(n_637)
);

O2A1O1Ixp5_ASAP7_75t_L g638 ( 
.A1(n_577),
.A2(n_572),
.B(n_591),
.C(n_579),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_R g639 ( 
.A(n_585),
.B(n_598),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_571),
.A2(n_570),
.B(n_563),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_584),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_588),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_595),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_573),
.B(n_555),
.Y(n_644)
);

AO32x2_ASAP7_75t_L g645 ( 
.A1(n_543),
.A2(n_558),
.A3(n_602),
.B1(n_608),
.B2(n_551),
.Y(n_645)
);

AO31x2_ASAP7_75t_L g646 ( 
.A1(n_602),
.A2(n_608),
.A3(n_606),
.B(n_567),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_552),
.B(n_541),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_568),
.B(n_562),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_609),
.Y(n_649)
);

AO32x2_ASAP7_75t_L g650 ( 
.A1(n_565),
.A2(n_583),
.A3(n_581),
.B1(n_589),
.B2(n_607),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_605),
.A2(n_592),
.B1(n_599),
.B2(n_564),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_569),
.A2(n_535),
.B(n_603),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_600),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_584),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_604),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_586),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_586),
.B(n_536),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_563),
.A2(n_390),
.B1(n_553),
.B2(n_361),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_542),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_554),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_559),
.A2(n_424),
.B(n_596),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_554),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_SL g664 ( 
.A1(n_560),
.A2(n_481),
.B(n_475),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_584),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_584),
.Y(n_666)
);

OAI22x1_ASAP7_75t_L g667 ( 
.A1(n_557),
.A2(n_464),
.B1(n_394),
.B2(n_472),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_593),
.B(n_549),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_559),
.A2(n_424),
.B(n_596),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_554),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_559),
.A2(n_424),
.B(n_596),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_536),
.B(n_381),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_539),
.B(n_475),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_542),
.Y(n_674)
);

O2A1O1Ixp5_ASAP7_75t_L g675 ( 
.A1(n_547),
.A2(n_577),
.B(n_572),
.C(n_576),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_536),
.B(n_381),
.Y(n_676)
);

CKINVDCx12_ASAP7_75t_R g677 ( 
.A(n_556),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_561),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_593),
.B(n_549),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_554),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_536),
.B(n_381),
.Y(n_681)
);

NAND2x1p5_ASAP7_75t_L g682 ( 
.A(n_561),
.B(n_546),
.Y(n_682)
);

A2O1A1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_559),
.A2(n_580),
.B(n_596),
.C(n_470),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_561),
.Y(n_684)
);

A2O1A1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_559),
.A2(n_580),
.B(n_596),
.C(n_470),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_559),
.A2(n_580),
.B(n_596),
.C(n_470),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_536),
.B(n_381),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_536),
.B(n_381),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_554),
.Y(n_689)
);

AO21x1_ASAP7_75t_L g690 ( 
.A1(n_545),
.A2(n_608),
.B(n_576),
.Y(n_690)
);

AO31x2_ASAP7_75t_L g691 ( 
.A1(n_547),
.A2(n_591),
.A3(n_610),
.B(n_545),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_561),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_546),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_542),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_536),
.B(n_381),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_546),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_554),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_549),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_554),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_539),
.B(n_475),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_554),
.Y(n_701)
);

NAND3x1_ASAP7_75t_L g702 ( 
.A(n_560),
.B(n_527),
.C(n_285),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_563),
.A2(n_390),
.B1(n_553),
.B2(n_361),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_556),
.B(n_475),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_554),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_683),
.A2(n_686),
.B(n_685),
.Y(n_706)
);

NOR2xp67_ASAP7_75t_L g707 ( 
.A(n_667),
.B(n_641),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_670),
.B(n_705),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_627),
.B(n_664),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_673),
.B(n_700),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_705),
.B(n_684),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_635),
.A2(n_659),
.B(n_703),
.C(n_634),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_680),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_665),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_692),
.B(n_678),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_612),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_672),
.B(n_676),
.Y(n_717)
);

OAI21x1_ASAP7_75t_SL g718 ( 
.A1(n_622),
.A2(n_647),
.B(n_658),
.Y(n_718)
);

NAND2x1p5_ASAP7_75t_L g719 ( 
.A(n_612),
.B(n_637),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_681),
.B(n_687),
.Y(n_720)
);

OA21x2_ASAP7_75t_L g721 ( 
.A1(n_630),
.A2(n_675),
.B(n_638),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_666),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_688),
.B(n_695),
.Y(n_723)
);

OA21x2_ASAP7_75t_L g724 ( 
.A1(n_616),
.A2(n_614),
.B(n_652),
.Y(n_724)
);

BUFx12f_ASAP7_75t_L g725 ( 
.A(n_655),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_L g726 ( 
.A1(n_618),
.A2(n_617),
.B(n_625),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_613),
.B(n_663),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_661),
.B(n_699),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_624),
.A2(n_623),
.B(n_651),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_693),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_701),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_689),
.Y(n_732)
);

AO21x2_ASAP7_75t_L g733 ( 
.A1(n_626),
.A2(n_645),
.B(n_648),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_696),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_628),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_644),
.A2(n_702),
.B1(n_697),
.B2(n_657),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_682),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_629),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_639),
.A2(n_704),
.B1(n_654),
.B2(n_657),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_620),
.B(n_611),
.Y(n_740)
);

NOR2xp67_ASAP7_75t_L g741 ( 
.A(n_653),
.B(n_632),
.Y(n_741)
);

NAND2x1p5_ASAP7_75t_L g742 ( 
.A(n_633),
.B(n_668),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_615),
.A2(n_649),
.B(n_691),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_677),
.B(n_631),
.Y(n_744)
);

AO21x2_ASAP7_75t_L g745 ( 
.A1(n_646),
.A2(n_650),
.B(n_642),
.Y(n_745)
);

OAI21x1_ASAP7_75t_L g746 ( 
.A1(n_646),
.A2(n_619),
.B(n_694),
.Y(n_746)
);

OAI21x1_ASAP7_75t_SL g747 ( 
.A1(n_633),
.A2(n_621),
.B(n_650),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_668),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_679),
.Y(n_749)
);

NAND2x1p5_ASAP7_75t_L g750 ( 
.A(n_633),
.B(n_679),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_698),
.A2(n_650),
.B(n_643),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_621),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_636),
.Y(n_753)
);

OA21x2_ASAP7_75t_L g754 ( 
.A1(n_660),
.A2(n_674),
.B(n_694),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_674),
.B(n_673),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_659),
.A2(n_703),
.B1(n_634),
.B2(n_563),
.Y(n_756)
);

AO31x2_ASAP7_75t_L g757 ( 
.A1(n_690),
.A2(n_640),
.A3(n_547),
.B(n_656),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_693),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_673),
.A2(n_700),
.B1(n_555),
.B2(n_634),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_662),
.A2(n_671),
.B(n_669),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_705),
.B(n_670),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_705),
.B(n_670),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_680),
.Y(n_763)
);

OAI21x1_ASAP7_75t_SL g764 ( 
.A1(n_622),
.A2(n_659),
.B(n_703),
.Y(n_764)
);

OAI21x1_ASAP7_75t_SL g765 ( 
.A1(n_622),
.A2(n_659),
.B(n_703),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_613),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_693),
.Y(n_767)
);

CKINVDCx14_ASAP7_75t_R g768 ( 
.A(n_641),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_664),
.B(n_468),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_613),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_683),
.A2(n_686),
.B(n_685),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_613),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_L g773 ( 
.A(n_664),
.B(n_607),
.C(n_583),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_664),
.B(n_468),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_743),
.B(n_746),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_773),
.A2(n_712),
.B(n_756),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_761),
.B(n_762),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_742),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_742),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_708),
.B(n_710),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_750),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_708),
.B(n_732),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_750),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_768),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_732),
.B(n_755),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_730),
.Y(n_786)
);

NAND2x1p5_ASAP7_75t_L g787 ( 
.A(n_753),
.B(n_754),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_713),
.B(n_763),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_717),
.B(n_720),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_734),
.Y(n_790)
);

INVx8_ASAP7_75t_L g791 ( 
.A(n_711),
.Y(n_791)
);

AO21x2_ASAP7_75t_L g792 ( 
.A1(n_706),
.A2(n_771),
.B(n_760),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_727),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_727),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_723),
.B(n_769),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_757),
.Y(n_796)
);

INVxp67_ASAP7_75t_SL g797 ( 
.A(n_728),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_754),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_728),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_711),
.Y(n_800)
);

BUFx12f_ASAP7_75t_L g801 ( 
.A(n_714),
.Y(n_801)
);

AO21x2_ASAP7_75t_L g802 ( 
.A1(n_706),
.A2(n_771),
.B(n_718),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_723),
.B(n_745),
.Y(n_803)
);

BUFx8_ASAP7_75t_L g804 ( 
.A(n_725),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_731),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_766),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_770),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_757),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_772),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_757),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_735),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_738),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_767),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_753),
.Y(n_814)
);

AOI21xp33_ASAP7_75t_L g815 ( 
.A1(n_712),
.A2(n_709),
.B(n_736),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_745),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_724),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_758),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_769),
.B(n_774),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_774),
.B(n_740),
.Y(n_820)
);

NOR2x1_ASAP7_75t_L g821 ( 
.A(n_739),
.B(n_736),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_780),
.B(n_751),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_782),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_819),
.A2(n_759),
.B1(n_740),
.B2(n_756),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_780),
.B(n_759),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_782),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_793),
.Y(n_827)
);

INVxp33_ASAP7_75t_L g828 ( 
.A(n_789),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_797),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_795),
.B(n_748),
.Y(n_830)
);

OAI322xp33_ASAP7_75t_L g831 ( 
.A1(n_820),
.A2(n_739),
.A3(n_749),
.B1(n_744),
.B2(n_719),
.C1(n_737),
.C2(n_716),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_778),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_803),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_789),
.B(n_744),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_785),
.B(n_802),
.Y(n_835)
);

INVx8_ASAP7_75t_L g836 ( 
.A(n_791),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_817),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_802),
.B(n_733),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_787),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_802),
.B(n_726),
.Y(n_840)
);

OAI221xp5_ASAP7_75t_L g841 ( 
.A1(n_776),
.A2(n_707),
.B1(n_741),
.B2(n_726),
.C(n_719),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_819),
.B(n_716),
.Y(n_842)
);

AND2x2_ASAP7_75t_SL g843 ( 
.A(n_775),
.B(n_747),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_791),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_792),
.B(n_777),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_817),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_791),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_814),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_805),
.B(n_715),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_788),
.B(n_721),
.Y(n_850)
);

AOI221xp5_ASAP7_75t_L g851 ( 
.A1(n_815),
.A2(n_765),
.B1(n_764),
.B2(n_715),
.C(n_722),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_806),
.B(n_752),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_788),
.B(n_721),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_791),
.B(n_729),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_791),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_807),
.B(n_809),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_775),
.B(n_798),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_816),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_845),
.B(n_808),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_823),
.B(n_826),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_858),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_845),
.B(n_808),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_835),
.B(n_808),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_837),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_835),
.B(n_810),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_848),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_846),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_839),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_857),
.Y(n_869)
);

INVx4_ASAP7_75t_L g870 ( 
.A(n_836),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_822),
.B(n_796),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_863),
.B(n_840),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_863),
.B(n_840),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_860),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_861),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_863),
.B(n_850),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_867),
.Y(n_877)
);

NAND2x1p5_ASAP7_75t_L g878 ( 
.A(n_870),
.B(n_847),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_864),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_860),
.B(n_833),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_859),
.B(n_853),
.Y(n_881)
);

NAND2x1_ASAP7_75t_L g882 ( 
.A(n_870),
.B(n_854),
.Y(n_882)
);

NAND2x1_ASAP7_75t_L g883 ( 
.A(n_870),
.B(n_854),
.Y(n_883)
);

CKINVDCx16_ASAP7_75t_R g884 ( 
.A(n_870),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_859),
.B(n_853),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_866),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_862),
.B(n_857),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_862),
.B(n_865),
.Y(n_888)
);

NOR2x1_ASAP7_75t_L g889 ( 
.A(n_868),
.B(n_847),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_871),
.B(n_856),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_862),
.B(n_838),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_L g892 ( 
.A(n_886),
.B(n_851),
.C(n_889),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_880),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_888),
.B(n_869),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_880),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_877),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_875),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_879),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_882),
.B(n_847),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_884),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_878),
.B(n_843),
.Y(n_901)
);

NAND2x2_ASAP7_75t_L g902 ( 
.A(n_882),
.B(n_832),
.Y(n_902)
);

OAI22xp33_ASAP7_75t_L g903 ( 
.A1(n_878),
.A2(n_829),
.B1(n_824),
.B2(n_841),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_888),
.B(n_869),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_883),
.B(n_832),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_897),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_SL g907 ( 
.A1(n_899),
.A2(n_878),
.B(n_821),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_894),
.B(n_887),
.Y(n_908)
);

NAND2x1_ASAP7_75t_L g909 ( 
.A(n_902),
.B(n_868),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_SL g910 ( 
.A1(n_899),
.A2(n_821),
.B(n_844),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_892),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_900),
.B(n_874),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_SL g913 ( 
.A1(n_901),
.A2(n_883),
.B(n_844),
.C(n_855),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_896),
.Y(n_914)
);

OAI322xp33_ASAP7_75t_L g915 ( 
.A1(n_896),
.A2(n_890),
.A3(n_825),
.B1(n_834),
.B2(n_873),
.C1(n_872),
.C2(n_875),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_898),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_893),
.B(n_872),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_895),
.B(n_873),
.Y(n_918)
);

AOI322xp5_ASAP7_75t_L g919 ( 
.A1(n_911),
.A2(n_903),
.A3(n_901),
.B1(n_904),
.B2(n_891),
.C1(n_876),
.C2(n_881),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_911),
.B(n_891),
.Y(n_920)
);

OR2x6_ASAP7_75t_L g921 ( 
.A(n_909),
.B(n_801),
.Y(n_921)
);

AOI21xp33_ASAP7_75t_L g922 ( 
.A1(n_907),
.A2(n_903),
.B(n_790),
.Y(n_922)
);

AOI211xp5_ASAP7_75t_L g923 ( 
.A1(n_913),
.A2(n_831),
.B(n_828),
.C(n_902),
.Y(n_923)
);

AOI21xp33_ASAP7_75t_L g924 ( 
.A1(n_910),
.A2(n_790),
.B(n_786),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_912),
.A2(n_887),
.B1(n_869),
.B2(n_885),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_920),
.B(n_914),
.Y(n_926)
);

NAND4xp25_ASAP7_75t_L g927 ( 
.A(n_922),
.B(n_830),
.C(n_849),
.D(n_842),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_921),
.A2(n_915),
.B(n_905),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_928),
.B(n_919),
.Y(n_929)
);

NOR2x1_ASAP7_75t_L g930 ( 
.A(n_927),
.B(n_804),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_930),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_929),
.B(n_926),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_931),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_SL g934 ( 
.A(n_932),
.B(n_784),
.Y(n_934)
);

OAI211xp5_ASAP7_75t_SL g935 ( 
.A1(n_933),
.A2(n_923),
.B(n_924),
.C(n_818),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_934),
.B(n_925),
.Y(n_936)
);

NAND4xp25_ASAP7_75t_L g937 ( 
.A(n_936),
.B(n_804),
.C(n_801),
.D(n_781),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_935),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_936),
.Y(n_939)
);

OAI22x1_ASAP7_75t_L g940 ( 
.A1(n_939),
.A2(n_804),
.B1(n_786),
.B2(n_813),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_938),
.A2(n_905),
.B1(n_813),
.B2(n_917),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_937),
.A2(n_918),
.B1(n_916),
.B2(n_906),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_939),
.B(n_916),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_939),
.B(n_804),
.Y(n_944)
);

XNOR2x1_ASAP7_75t_L g945 ( 
.A(n_940),
.B(n_778),
.Y(n_945)
);

OAI22x1_ASAP7_75t_L g946 ( 
.A1(n_944),
.A2(n_827),
.B1(n_855),
.B2(n_794),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_941),
.A2(n_783),
.B1(n_781),
.B2(n_779),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_943),
.A2(n_908),
.B(n_800),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_942),
.A2(n_781),
.B1(n_783),
.B2(n_778),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_944),
.A2(n_811),
.B(n_812),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_950),
.B(n_811),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_946),
.Y(n_952)
);

INVxp33_ASAP7_75t_L g953 ( 
.A(n_945),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_949),
.B(n_799),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_SL g955 ( 
.A1(n_953),
.A2(n_948),
.B(n_947),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_952),
.A2(n_779),
.B(n_783),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_951),
.A2(n_812),
.B(n_852),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_956),
.B(n_954),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_958),
.A2(n_955),
.B(n_957),
.Y(n_959)
);


endmodule