module real_jpeg_15965_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_0),
.B(n_150),
.Y(n_149)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_0),
.A2(n_100),
.A3(n_238),
.B1(n_240),
.B2(n_243),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_0),
.B(n_128),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_0),
.A2(n_64),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_0),
.A2(n_28),
.B1(n_359),
.B2(n_363),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_1),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_2),
.A2(n_119),
.B1(n_123),
.B2(n_127),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_2),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_2),
.A2(n_127),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_2),
.A2(n_127),
.B1(n_268),
.B2(n_272),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_2),
.A2(n_127),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_3),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_3),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_3),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_4),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_4),
.A2(n_45),
.B1(n_277),
.B2(n_436),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_4),
.A2(n_45),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_5),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_5),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_5),
.A2(n_132),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_5),
.A2(n_132),
.B1(n_341),
.B2(n_344),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_5),
.A2(n_132),
.B1(n_398),
.B2(n_400),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_6),
.A2(n_119),
.B1(n_177),
.B2(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_6),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_6),
.A2(n_180),
.B1(n_227),
.B2(n_231),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_6),
.A2(n_180),
.B1(n_281),
.B2(n_284),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_6),
.A2(n_180),
.B1(n_398),
.B2(n_449),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_7),
.A2(n_410),
.B1(n_412),
.B2(n_413),
.Y(n_409)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_7),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g485 ( 
.A1(n_7),
.A2(n_412),
.B1(n_486),
.B2(n_489),
.Y(n_485)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_8),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_8),
.Y(n_444)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_9),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_9),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_9),
.Y(n_204)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_9),
.Y(n_247)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_9),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_10),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_10),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_10),
.A2(n_141),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_10),
.A2(n_141),
.B1(n_456),
.B2(n_460),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_10),
.A2(n_141),
.B1(n_549),
.B2(n_552),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_11),
.A2(n_53),
.B1(n_56),
.B2(n_61),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_11),
.A2(n_61),
.B1(n_426),
.B2(n_428),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_11),
.A2(n_61),
.B1(n_529),
.B2(n_531),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_12),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_13),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_14),
.A2(n_183),
.B1(n_184),
.B2(n_188),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_14),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_14),
.A2(n_183),
.B1(n_251),
.B2(n_254),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_14),
.A2(n_183),
.B1(n_391),
.B2(n_393),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_14),
.A2(n_183),
.B1(n_501),
.B2(n_504),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g145 ( 
.A(n_15),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_16),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_418)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_16),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_16),
.A2(n_421),
.B1(n_539),
.B2(n_541),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g163 ( 
.A(n_17),
.Y(n_163)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_17),
.Y(n_404)
);

BUFx5_ASAP7_75t_L g452 ( 
.A(n_17),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_516),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_476),
.B(n_514),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_384),
.B(n_473),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_261),
.B(n_383),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_219),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_24),
.B(n_219),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_159),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_90),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_26),
.B(n_90),
.C(n_159),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_62),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_27),
.B(n_62),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_38),
.B1(n_50),
.B2(n_52),
.Y(n_27)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_28),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_28),
.A2(n_280),
.B1(n_286),
.B2(n_288),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_28),
.A2(n_340),
.B1(n_359),
.B2(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_28),
.A2(n_52),
.B1(n_409),
.B2(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_28),
.A2(n_368),
.B(n_418),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_31),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_31),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_32),
.Y(n_370)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_39),
.A2(n_137),
.B1(n_138),
.B2(n_146),
.Y(n_136)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_44),
.Y(n_140)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_44),
.Y(n_195)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_44),
.Y(n_197)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_44),
.Y(n_343)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_44),
.Y(n_345)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_47),
.Y(n_419)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_48),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_51),
.Y(n_287)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_54),
.Y(n_420)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_60),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_69),
.B1(n_79),
.B2(n_85),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_63),
.A2(n_64),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_64),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_64),
.B(n_320),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_SL g330 ( 
.A1(n_64),
.A2(n_319),
.B(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_64),
.B(n_355),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_64),
.B(n_218),
.Y(n_371)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_68),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_78),
.Y(n_179)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_83),
.Y(n_459)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_84),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_86),
.A2(n_151),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_87),
.Y(n_553)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_136),
.C(n_149),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_91),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_117),
.B1(n_128),
.B2(n_129),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_92),
.A2(n_128),
.B1(n_129),
.B2(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_92),
.A2(n_128),
.B1(n_526),
.B2(n_527),
.Y(n_525)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_93),
.A2(n_118),
.B1(n_297),
.B2(n_302),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_93),
.A2(n_302),
.B1(n_389),
.B2(n_390),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_93),
.A2(n_302),
.B1(n_390),
.B2(n_455),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_93),
.A2(n_302),
.B1(n_455),
.B2(n_507),
.Y(n_506)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_100),
.B(n_104),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_112),
.B2(n_114),
.Y(n_104)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_106),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_106),
.Y(n_427)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_107),
.Y(n_271)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_107),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_107),
.Y(n_333)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_128),
.Y(n_302)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_130),
.Y(n_508)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_131),
.Y(n_298)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_131),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_134),
.Y(n_393)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_134),
.Y(n_460)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_136),
.B(n_149),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_137),
.A2(n_138),
.B1(n_250),
.B2(n_257),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_137),
.A2(n_339),
.B1(n_346),
.B2(n_347),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_137),
.A2(n_408),
.B1(n_415),
.B2(n_417),
.Y(n_407)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_139),
.Y(n_285)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_140),
.Y(n_360)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_140),
.Y(n_411)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_144),
.Y(n_283)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_145),
.Y(n_256)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_145),
.Y(n_327)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_161),
.B1(n_164),
.B2(n_170),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_150),
.A2(n_164),
.B1(n_170),
.B2(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_150),
.Y(n_453)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_155),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_156),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_174),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_160),
.B(n_175),
.C(n_181),
.Y(n_467)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_163),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_164),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_181),
.Y(n_174)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_176),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_191),
.B1(n_210),
.B2(n_217),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_184),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_191),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_191),
.A2(n_217),
.B1(n_267),
.B2(n_276),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_191),
.A2(n_217),
.B1(n_226),
.B2(n_276),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_191),
.A2(n_217),
.B1(n_267),
.B2(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_191),
.B(n_434),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_191),
.A2(n_217),
.B1(n_537),
.B2(n_538),
.Y(n_536)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_202),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_205),
.B1(n_207),
.B2(n_209),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_207),
.Y(n_318)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_208),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_209),
.Y(n_436)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_209),
.Y(n_541)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_211),
.A2(n_218),
.B1(n_224),
.B2(n_435),
.Y(n_439)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_217),
.B(n_424),
.Y(n_423)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_224),
.B1(n_225),
.B2(n_234),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_218),
.A2(n_224),
.B1(n_425),
.B2(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.C(n_235),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_220),
.A2(n_221),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_223),
.A2(n_235),
.B1(n_236),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_223),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_230),
.Y(n_275)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_230),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_233),
.Y(n_432)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_248),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_237),
.A2(n_248),
.B1(n_249),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_238),
.Y(n_509)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_251),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21x1_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_376),
.B(n_382),
.Y(n_261)
);

AOI21x1_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_305),
.B(n_375),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_291),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_264),
.B(n_291),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_279),
.C(n_289),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_265),
.A2(n_266),
.B1(n_289),
.B2(n_290),
.Y(n_335)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_335),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_280),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_292),
.B(n_295),
.C(n_304),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_303),
.B2(n_304),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_336),
.B(n_374),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_334),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_307),
.B(n_334),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_328),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_308),
.A2(n_328),
.B1(n_329),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_308),
.Y(n_349)
);

OAI32xp33_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_312),
.A3(n_316),
.B1(n_319),
.B2(n_323),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_311),
.Y(n_488)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_321),
.Y(n_540)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_350),
.B(n_373),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_348),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_348),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_366),
.B(n_372),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_358),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_365),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_371),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_371),
.Y(n_372)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_381),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_381),
.Y(n_382)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_461),
.B(n_468),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_385),
.B(n_461),
.C(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_405),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_386),
.B(n_406),
.C(n_437),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_394),
.C(n_395),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_388),
.B(n_395),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_394),
.B(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_397),
.A2(n_447),
.B1(n_448),
.B2(n_453),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx8_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_403),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_404),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_437),
.Y(n_405)
);

XNOR2x2_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_422),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_407),
.A2(n_423),
.B(n_433),
.Y(n_510)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_433),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_435),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_445),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_438),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

XOR2x2_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_440),
.Y(n_465)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_454),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_446),
.Y(n_480)
);

OAI22x1_ASAP7_75t_L g499 ( 
.A1(n_447),
.A2(n_448),
.B1(n_453),
.B2(n_500),
.Y(n_499)
);

OAI22x1_ASAP7_75t_L g547 ( 
.A1(n_447),
.A2(n_453),
.B1(n_500),
.B2(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_450),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_480),
.C(n_481),
.Y(n_479)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_465),
.C(n_466),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_462),
.A2(n_463),
.B1(n_471),
.B2(n_472),
.Y(n_470)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_465),
.B(n_467),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_469),
.B(n_470),
.Y(n_475)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_471),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_478),
.B(n_513),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_478),
.B(n_513),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_479),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_483),
.A2(n_497),
.B1(n_511),
.B2(n_512),
.Y(n_482)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_483),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_483),
.B(n_512),
.C(n_519),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_484),
.A2(n_494),
.B1(n_495),
.B2(n_496),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_484),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_484),
.B(n_495),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_485),
.Y(n_537)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_494),
.A2(n_495),
.B1(n_546),
.B2(n_547),
.Y(n_545)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_497),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_510),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_506),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_510),
.C(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_506),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_507),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_515),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_556),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_520),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_518),
.B(n_520),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_523),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_543),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_525),
.A2(n_536),
.B(n_542),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_525),
.B(n_536),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_544),
.A2(n_545),
.B1(n_554),
.B2(n_555),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx6_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx6_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_554),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);


endmodule