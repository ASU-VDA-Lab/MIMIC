module real_aes_9211_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_SL g247 ( .A1(n_0), .A2(n_248), .B(n_249), .C(n_253), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_1), .B(n_242), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_2), .B(n_228), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_3), .A2(n_236), .B(n_322), .Y(n_321) );
AO21x2_ASAP7_75t_L g329 ( .A1(n_4), .A2(n_209), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g200 ( .A(n_5), .Y(n_200) );
AND2x6_ASAP7_75t_L g234 ( .A(n_5), .B(n_198), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_5), .B(n_520), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_6), .A2(n_180), .B1(n_181), .B2(n_184), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_6), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_6), .A2(n_217), .B(n_234), .C(n_300), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_7), .A2(n_39), .B1(n_182), .B2(n_183), .Y(n_181) );
INVx1_ASAP7_75t_L g183 ( .A(n_7), .Y(n_183) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_8), .A2(n_20), .B1(n_91), .B2(n_92), .Y(n_90) );
INVx1_ASAP7_75t_L g214 ( .A(n_9), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_10), .B(n_228), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_11), .A2(n_81), .B1(n_82), .B2(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_11), .Y(n_526) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_12), .A2(n_22), .B1(n_91), .B2(n_95), .Y(n_94) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_13), .A2(n_81), .B1(n_82), .B2(n_170), .Y(n_80) );
INVx1_ASAP7_75t_L g170 ( .A(n_13), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_14), .A2(n_217), .B(n_262), .C(n_269), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_15), .A2(n_217), .B(n_269), .C(n_333), .Y(n_332) );
AOI22xp5_ASAP7_75t_SL g515 ( .A1(n_15), .A2(n_81), .B1(n_82), .B2(n_516), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_15), .Y(n_516) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_16), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_17), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_18), .A2(n_236), .B(n_244), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_19), .A2(n_179), .B1(n_185), .B2(n_186), .Y(n_178) );
INVx1_ASAP7_75t_L g185 ( .A(n_19), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_19), .A2(n_232), .B(n_285), .C(n_286), .Y(n_284) );
INVx2_ASAP7_75t_L g219 ( .A(n_21), .Y(n_219) );
OAI221xp5_ASAP7_75t_L g191 ( .A1(n_22), .A2(n_41), .B1(n_52), .B2(n_192), .C(n_193), .Y(n_191) );
INVxp67_ASAP7_75t_L g194 ( .A(n_22), .Y(n_194) );
AOI22xp33_ASAP7_75t_SL g156 ( .A1(n_23), .A2(n_60), .B1(n_157), .B2(n_160), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_24), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_25), .B(n_260), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_26), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_27), .A2(n_46), .B1(n_127), .B2(n_134), .Y(n_126) );
AOI22xp33_ASAP7_75t_SL g117 ( .A1(n_28), .A2(n_36), .B1(n_118), .B2(n_122), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_29), .B(n_228), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_30), .B(n_236), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_31), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g312 ( .A1(n_32), .A2(n_232), .B(n_285), .C(n_313), .Y(n_312) );
AOI22xp33_ASAP7_75t_SL g163 ( .A1(n_33), .A2(n_53), .B1(n_164), .B2(n_167), .Y(n_163) );
AOI22xp33_ASAP7_75t_SL g138 ( .A1(n_34), .A2(n_63), .B1(n_139), .B2(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g250 ( .A(n_35), .Y(n_250) );
INVx1_ASAP7_75t_L g314 ( .A(n_37), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_38), .B(n_236), .Y(n_311) );
INVx1_ASAP7_75t_L g182 ( .A(n_39), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_40), .Y(n_274) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_41), .A2(n_65), .B1(n_91), .B2(n_95), .Y(n_98) );
INVxp67_ASAP7_75t_L g195 ( .A(n_41), .Y(n_195) );
INVx1_ASAP7_75t_L g198 ( .A(n_42), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_43), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_44), .B(n_242), .Y(n_327) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_45), .A2(n_224), .B(n_268), .C(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g213 ( .A(n_47), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_48), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_49), .B(n_228), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_50), .B(n_229), .Y(n_301) );
INVx1_ASAP7_75t_L g176 ( .A(n_51), .Y(n_176) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_52), .A2(n_70), .B1(n_91), .B2(n_92), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_54), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_55), .B(n_264), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_56), .A2(n_217), .B(n_222), .C(n_232), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g323 ( .A(n_57), .Y(n_323) );
AOI22xp33_ASAP7_75t_SL g146 ( .A1(n_58), .A2(n_59), .B1(n_147), .B2(n_151), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_61), .B(n_266), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_62), .A2(n_174), .B1(n_175), .B2(n_177), .Y(n_173) );
INVx1_ASAP7_75t_L g177 ( .A(n_62), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_64), .Y(n_291) );
INVx2_ASAP7_75t_L g211 ( .A(n_66), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_67), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_68), .B(n_252), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_69), .B(n_236), .Y(n_283) );
INVx1_ASAP7_75t_L g287 ( .A(n_71), .Y(n_287) );
INVxp67_ASAP7_75t_L g326 ( .A(n_72), .Y(n_326) );
INVx1_ASAP7_75t_L g91 ( .A(n_73), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_73), .Y(n_93) );
INVx1_ASAP7_75t_L g223 ( .A(n_74), .Y(n_223) );
INVx1_ASAP7_75t_L g297 ( .A(n_75), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_76), .Y(n_101) );
AND2x2_ASAP7_75t_L g316 ( .A(n_77), .B(n_272), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_188), .B1(n_201), .B2(n_511), .C(n_514), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_171), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NAND3xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_137), .C(n_155), .Y(n_83) );
NOR2xp33_ASAP7_75t_L g84 ( .A(n_85), .B(n_116), .Y(n_84) );
OAI222xp33_ASAP7_75t_L g85 ( .A1(n_86), .A2(n_101), .B1(n_102), .B2(n_109), .C1(n_110), .C2(n_115), .Y(n_85) );
BUFx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx4_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x6_ASAP7_75t_L g88 ( .A(n_89), .B(n_96), .Y(n_88) );
AND2x4_ASAP7_75t_L g123 ( .A(n_89), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_94), .Y(n_89) );
AND2x2_ASAP7_75t_L g108 ( .A(n_90), .B(n_98), .Y(n_108) );
INVx2_ASAP7_75t_L g133 ( .A(n_90), .Y(n_133) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g95 ( .A(n_93), .Y(n_95) );
INVx2_ASAP7_75t_L g107 ( .A(n_94), .Y(n_107) );
INVx1_ASAP7_75t_L g121 ( .A(n_94), .Y(n_121) );
OR2x2_ASAP7_75t_L g132 ( .A(n_94), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g136 ( .A(n_94), .B(n_133), .Y(n_136) );
AND2x4_ASAP7_75t_L g140 ( .A(n_96), .B(n_136), .Y(n_140) );
AND2x6_ASAP7_75t_L g159 ( .A(n_96), .B(n_131), .Y(n_159) );
AND2x2_ASAP7_75t_L g166 ( .A(n_96), .B(n_145), .Y(n_166) );
AND2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_99), .Y(n_96) );
AND2x2_ASAP7_75t_L g130 ( .A(n_97), .B(n_100), .Y(n_130) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g144 ( .A(n_98), .B(n_125), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_98), .B(n_100), .Y(n_154) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g106 ( .A(n_100), .Y(n_106) );
INVx1_ASAP7_75t_L g125 ( .A(n_100), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g114 ( .A(n_106), .Y(n_114) );
AND2x2_ASAP7_75t_L g145 ( .A(n_107), .B(n_133), .Y(n_145) );
AND2x4_ASAP7_75t_L g113 ( .A(n_108), .B(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g119 ( .A(n_108), .B(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx4f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_126), .Y(n_116) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x6_ASAP7_75t_L g153 ( .A(n_121), .B(n_154), .Y(n_153) );
BUFx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx5_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x6_ASAP7_75t_L g135 ( .A(n_130), .B(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g169 ( .A(n_130), .B(n_145), .Y(n_169) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g150 ( .A(n_136), .B(n_144), .Y(n_150) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_146), .Y(n_137) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x4_ASAP7_75t_L g161 ( .A(n_145), .B(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx8_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx6_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_163), .Y(n_155) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx11_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B1(n_178), .B2(n_187), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_178), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_179), .Y(n_186) );
INVx1_ASAP7_75t_L g184 ( .A(n_181), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
AND3x1_ASAP7_75t_SL g190 ( .A(n_191), .B(n_196), .C(n_199), .Y(n_190) );
INVxp67_ASAP7_75t_L g520 ( .A(n_191), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx1_ASAP7_75t_SL g521 ( .A(n_196), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_196), .A2(n_217), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g528 ( .A(n_196), .Y(n_528) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_197), .B(n_200), .Y(n_524) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_SL g527 ( .A(n_199), .B(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_200), .Y(n_199) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OR3x1_ASAP7_75t_L g202 ( .A(n_203), .B(n_419), .C(n_468), .Y(n_202) );
NAND5xp2_ASAP7_75t_L g203 ( .A(n_204), .B(n_353), .C(n_382), .D(n_390), .E(n_405), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_276), .B(n_292), .C(n_337), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_256), .Y(n_205) );
AND2x2_ASAP7_75t_L g348 ( .A(n_206), .B(n_345), .Y(n_348) );
AND2x2_ASAP7_75t_L g381 ( .A(n_206), .B(n_257), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_206), .B(n_280), .Y(n_474) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_241), .Y(n_206) );
INVx2_ASAP7_75t_L g279 ( .A(n_207), .Y(n_279) );
BUFx2_ASAP7_75t_L g448 ( .A(n_207), .Y(n_448) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_215), .B(n_239), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_208), .B(n_240), .Y(n_239) );
INVx3_ASAP7_75t_L g242 ( .A(n_208), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_208), .B(n_291), .Y(n_290) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_208), .A2(n_296), .B(n_306), .Y(n_295) );
INVx4_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_209), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_209), .A2(n_331), .B(n_332), .Y(n_330) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g308 ( .A(n_210), .Y(n_308) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AND2x2_ASAP7_75t_SL g272 ( .A(n_211), .B(n_212), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_235), .Y(n_215) );
INVx5_ASAP7_75t_L g246 ( .A(n_217), .Y(n_246) );
AND2x2_ASAP7_75t_L g513 ( .A(n_217), .B(n_269), .Y(n_513) );
AND2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_218), .Y(n_231) );
BUFx3_ASAP7_75t_L g254 ( .A(n_218), .Y(n_254) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g238 ( .A(n_219), .Y(n_238) );
INVx1_ASAP7_75t_L g305 ( .A(n_219), .Y(n_305) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_221), .Y(n_226) );
INVx3_ASAP7_75t_L g229 ( .A(n_221), .Y(n_229) );
AND2x2_ASAP7_75t_L g237 ( .A(n_221), .B(n_238), .Y(n_237) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_221), .Y(n_252) );
INVx1_ASAP7_75t_L g335 ( .A(n_221), .Y(n_335) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_227), .C(n_230), .Y(n_222) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g264 ( .A(n_226), .Y(n_264) );
INVx2_ASAP7_75t_L g248 ( .A(n_228), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_228), .B(n_326), .Y(n_325) );
INVx5_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g244 ( .A1(n_233), .A2(n_245), .B(n_246), .C(n_247), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_233), .A2(n_246), .B(n_323), .C(n_324), .Y(n_322) );
INVx4_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
AND2x4_ASAP7_75t_L g236 ( .A(n_234), .B(n_237), .Y(n_236) );
BUFx3_ASAP7_75t_L g269 ( .A(n_234), .Y(n_269) );
NAND2x1p5_ASAP7_75t_L g298 ( .A(n_234), .B(n_237), .Y(n_298) );
BUFx2_ASAP7_75t_L g260 ( .A(n_236), .Y(n_260) );
INVx1_ASAP7_75t_L g268 ( .A(n_238), .Y(n_268) );
AND2x2_ASAP7_75t_L g256 ( .A(n_241), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g346 ( .A(n_241), .Y(n_346) );
AND2x2_ASAP7_75t_L g432 ( .A(n_241), .B(n_345), .Y(n_432) );
AND2x2_ASAP7_75t_L g487 ( .A(n_241), .B(n_279), .Y(n_487) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_255), .Y(n_241) );
INVx2_ASAP7_75t_L g285 ( .A(n_246), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx4_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_254), .Y(n_289) );
INVx1_ASAP7_75t_L g404 ( .A(n_256), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_256), .B(n_280), .Y(n_451) );
INVx5_ASAP7_75t_L g345 ( .A(n_257), .Y(n_345) );
AND2x4_ASAP7_75t_L g366 ( .A(n_257), .B(n_346), .Y(n_366) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_257), .Y(n_388) );
AND2x2_ASAP7_75t_L g463 ( .A(n_257), .B(n_448), .Y(n_463) );
AND2x2_ASAP7_75t_L g466 ( .A(n_257), .B(n_281), .Y(n_466) );
OR2x6_ASAP7_75t_L g257 ( .A(n_258), .B(n_273), .Y(n_257) );
AOI21xp5_ASAP7_75t_SL g258 ( .A1(n_259), .A2(n_261), .B(n_270), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_265), .B(n_267), .Y(n_262) );
INVx2_ASAP7_75t_L g266 ( .A(n_264), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_266), .A2(n_287), .B(n_288), .C(n_289), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_266), .A2(n_289), .B(n_314), .C(n_315), .Y(n_313) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g275 ( .A(n_272), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_272), .A2(n_283), .B(n_284), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_272), .A2(n_311), .B(n_312), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_276), .B(n_346), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_276), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
AND2x2_ASAP7_75t_L g371 ( .A(n_278), .B(n_346), .Y(n_371) );
AND2x2_ASAP7_75t_L g389 ( .A(n_278), .B(n_281), .Y(n_389) );
INVx1_ASAP7_75t_L g409 ( .A(n_278), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_278), .B(n_345), .Y(n_454) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_278), .Y(n_496) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_279), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_280), .B(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_280), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_280), .A2(n_341), .B(n_402), .C(n_404), .Y(n_401) );
AND2x2_ASAP7_75t_L g408 ( .A(n_280), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g417 ( .A(n_280), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g421 ( .A(n_280), .B(n_345), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_280), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g436 ( .A(n_280), .B(n_346), .Y(n_436) );
AND2x2_ASAP7_75t_L g486 ( .A(n_280), .B(n_487), .Y(n_486) );
INVx5_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx2_ASAP7_75t_L g350 ( .A(n_281), .Y(n_350) );
AND2x2_ASAP7_75t_L g391 ( .A(n_281), .B(n_344), .Y(n_391) );
AND2x2_ASAP7_75t_L g403 ( .A(n_281), .B(n_378), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_281), .B(n_432), .Y(n_450) );
OR2x6_ASAP7_75t_L g281 ( .A(n_282), .B(n_290), .Y(n_281) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_317), .Y(n_292) );
INVx1_ASAP7_75t_L g339 ( .A(n_293), .Y(n_339) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_309), .Y(n_293) );
OR2x2_ASAP7_75t_L g341 ( .A(n_294), .B(n_309), .Y(n_341) );
NAND3xp33_ASAP7_75t_L g347 ( .A(n_294), .B(n_348), .C(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_294), .B(n_319), .Y(n_358) );
OR2x2_ASAP7_75t_L g373 ( .A(n_294), .B(n_361), .Y(n_373) );
AND2x2_ASAP7_75t_L g379 ( .A(n_294), .B(n_328), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_294), .B(n_510), .Y(n_509) );
INVx5_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_295), .B(n_319), .Y(n_376) );
AND2x2_ASAP7_75t_L g415 ( .A(n_295), .B(n_329), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_295), .B(n_328), .Y(n_443) );
OR2x2_ASAP7_75t_L g446 ( .A(n_295), .B(n_328), .Y(n_446) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_299), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B(n_303), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_303), .A2(n_334), .B(n_336), .Y(n_333) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx5_ASAP7_75t_SL g361 ( .A(n_309), .Y(n_361) );
OR2x2_ASAP7_75t_L g367 ( .A(n_309), .B(n_318), .Y(n_367) );
AND2x2_ASAP7_75t_L g383 ( .A(n_309), .B(n_384), .Y(n_383) );
AOI321xp33_ASAP7_75t_L g390 ( .A1(n_309), .A2(n_391), .A3(n_392), .B1(n_393), .B2(n_399), .C(n_401), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_309), .B(n_317), .Y(n_400) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_309), .Y(n_413) );
OR2x2_ASAP7_75t_L g460 ( .A(n_309), .B(n_358), .Y(n_460) );
AND2x2_ASAP7_75t_L g482 ( .A(n_309), .B(n_379), .Y(n_482) );
AND2x2_ASAP7_75t_L g501 ( .A(n_309), .B(n_319), .Y(n_501) );
OR2x6_ASAP7_75t_L g309 ( .A(n_310), .B(n_316), .Y(n_309) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_328), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_319), .B(n_328), .Y(n_342) );
AND2x2_ASAP7_75t_L g351 ( .A(n_319), .B(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g378 ( .A(n_319), .Y(n_378) );
AND2x2_ASAP7_75t_L g384 ( .A(n_319), .B(n_379), .Y(n_384) );
INVxp67_ASAP7_75t_L g414 ( .A(n_319), .Y(n_414) );
OR2x2_ASAP7_75t_L g456 ( .A(n_319), .B(n_361), .Y(n_456) );
OA21x2_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_321), .B(n_327), .Y(n_319) );
OR2x2_ASAP7_75t_L g338 ( .A(n_328), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g352 ( .A(n_328), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_328), .B(n_341), .Y(n_385) );
AND2x2_ASAP7_75t_L g434 ( .A(n_328), .B(n_378), .Y(n_434) );
AND2x2_ASAP7_75t_L g472 ( .A(n_328), .B(n_361), .Y(n_472) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_329), .B(n_361), .Y(n_360) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B(n_343), .C(n_347), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_338), .A2(n_340), .B1(n_465), .B2(n_467), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_340), .A2(n_363), .B1(n_418), .B2(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_SL g492 ( .A(n_341), .Y(n_492) );
INVx1_ASAP7_75t_SL g392 ( .A(n_342), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_344), .B(n_364), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g405 ( .A1(n_344), .A2(n_385), .B1(n_392), .B2(n_406), .C1(n_410), .C2(n_416), .Y(n_405) );
AND2x2_ASAP7_75t_L g495 ( .A(n_344), .B(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx2_ASAP7_75t_L g370 ( .A(n_345), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_345), .B(n_365), .Y(n_440) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_345), .Y(n_477) );
AND2x2_ASAP7_75t_L g480 ( .A(n_345), .B(n_389), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_345), .B(n_496), .Y(n_506) );
INVx1_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_346), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_348), .A2(n_489), .B(n_490), .C(n_493), .Y(n_488) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_350), .B(n_412), .C(n_415), .Y(n_411) );
OR2x2_ASAP7_75t_L g439 ( .A(n_350), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_350), .B(n_366), .Y(n_467) );
OR2x2_ASAP7_75t_L g372 ( .A(n_352), .B(n_373), .Y(n_372) );
AOI211xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .B(n_362), .C(n_374), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_355), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g461 ( .A(n_356), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_357), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g375 ( .A(n_360), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_361), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g429 ( .A(n_361), .B(n_379), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_361), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_361), .B(n_378), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B1(n_368), .B2(n_372), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_364), .B(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_366), .B(n_408), .Y(n_407) );
OAI221xp5_ASAP7_75t_SL g430 ( .A1(n_367), .A2(n_431), .B1(n_433), .B2(n_435), .C(n_437), .Y(n_430) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AND2x2_ASAP7_75t_L g485 ( .A(n_370), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g498 ( .A(n_370), .B(n_487), .Y(n_498) );
INVx1_ASAP7_75t_L g418 ( .A(n_371), .Y(n_418) );
INVx1_ASAP7_75t_L g489 ( .A(n_372), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_373), .A2(n_456), .B(n_479), .Y(n_478) );
AOI21xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B(n_380), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI21xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_385), .B(n_386), .Y(n_382) );
INVx1_ASAP7_75t_L g422 ( .A(n_383), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_384), .A2(n_470), .B1(n_473), .B2(n_475), .C(n_478), .Y(n_469) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_392), .A2(n_482), .B1(n_483), .B2(n_485), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g458 ( .A(n_394), .Y(n_458) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR2xp67_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g462 ( .A(n_398), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g427 ( .A(n_403), .Y(n_427) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_408), .B(n_432), .Y(n_484) );
INVxp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_414), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g500 ( .A(n_415), .B(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g507 ( .A(n_415), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI211xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_422), .B(n_423), .C(n_457), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI211xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B(n_430), .C(n_449), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g510 ( .A(n_434), .Y(n_510) );
AND2x2_ASAP7_75t_L g447 ( .A(n_436), .B(n_448), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_441), .B1(n_445), .B2(n_447), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
OR2x2_ASAP7_75t_L g455 ( .A(n_443), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g508 ( .A(n_444), .Y(n_508) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI31xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .A3(n_452), .B(n_455), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI211xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_461), .C(n_464), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
NAND5xp2_ASAP7_75t_L g468 ( .A(n_469), .B(n_481), .C(n_488), .D(n_502), .E(n_505), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_480), .A2(n_506), .B1(n_507), .B2(n_509), .Y(n_505) );
INVx1_ASAP7_75t_SL g504 ( .A(n_482), .Y(n_504) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_497), .B(n_499), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVxp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
OAI322xp33_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .A3(n_517), .B1(n_521), .B2(n_522), .C1(n_525), .C2(n_527), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
endmodule