module fake_jpeg_12504_n_391 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_391);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_391;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_74),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_4),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_60),
.B(n_67),
.Y(n_131)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_21),
.A2(n_37),
.B(n_53),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_66),
.B(n_100),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_34),
.B(n_4),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_4),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_70),
.B(n_92),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_73),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_76),
.Y(n_179)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_84),
.Y(n_139)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_5),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_86),
.B(n_89),
.Y(n_129)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_23),
.B(n_5),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_7),
.B1(n_10),
.B2(n_12),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_53),
.B1(n_52),
.B2(n_46),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_16),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_93),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_24),
.Y(n_97)
);

CKINVDCx12_ASAP7_75t_R g164 ( 
.A(n_97),
.Y(n_164)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_49),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_31),
.B(n_7),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_102),
.B(n_14),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_104),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_37),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_107),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_42),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_109),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_111),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_46),
.B(n_52),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_113),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_63),
.A2(n_44),
.B1(n_51),
.B2(n_48),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_125),
.A2(n_133),
.B1(n_141),
.B2(n_127),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_44),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_126),
.B(n_149),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_40),
.B1(n_48),
.B2(n_45),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_59),
.A2(n_40),
.B(n_45),
.C(n_43),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_143),
.A2(n_112),
.B(n_156),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_43),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_51),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_152),
.B(n_154),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_10),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_165),
.Y(n_182)
);

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_93),
.B(n_15),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_170),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_16),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_75),
.B(n_83),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_166),
.B(n_169),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_72),
.A2(n_98),
.B1(n_78),
.B2(n_83),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_168),
.A2(n_174),
.B(n_180),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_75),
.B(n_80),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_93),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_171),
.B(n_172),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_58),
.B(n_62),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_91),
.A2(n_64),
.B1(n_71),
.B2(n_76),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_88),
.B(n_81),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_156),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_101),
.B(n_65),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_180),
.Y(n_194)
);

OR2x4_ASAP7_75t_L g178 ( 
.A(n_66),
.B(n_65),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_116),
.Y(n_227)
);

NAND2x1_ASAP7_75t_L g180 ( 
.A(n_65),
.B(n_32),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_60),
.B(n_70),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_131),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_171),
.A2(n_178),
.B(n_157),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_183),
.B(n_222),
.C(n_227),
.Y(n_279)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_195),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_187),
.B(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_189),
.B(n_191),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_177),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_115),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_203),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_194),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_117),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_196),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_130),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_150),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_140),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_206),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_137),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_216),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_133),
.A2(n_174),
.B1(n_141),
.B2(n_125),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_208),
.A2(n_214),
.B1(n_225),
.B2(n_232),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_114),
.B(n_158),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_213),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_145),
.A2(n_162),
.B1(n_137),
.B2(n_116),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_223),
.B1(n_230),
.B2(n_227),
.Y(n_240)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_162),
.Y(n_211)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_211),
.Y(n_266)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_142),
.B(n_151),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_168),
.A2(n_173),
.B1(n_145),
.B2(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_148),
.Y(n_215)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_119),
.B(n_121),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_151),
.B(n_147),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_221),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_163),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_220),
.Y(n_259)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_121),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_148),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_144),
.B(n_128),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_144),
.B(n_139),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_228),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_163),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_147),
.B(n_132),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_231),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_136),
.A2(n_123),
.B1(n_134),
.B2(n_132),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_238),
.Y(n_244)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_136),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_123),
.A2(n_134),
.B1(n_179),
.B2(n_164),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_179),
.A2(n_171),
.B1(n_178),
.B2(n_133),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_233),
.A2(n_217),
.B1(n_229),
.B2(n_222),
.Y(n_275)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_124),
.Y(n_234)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_138),
.B(n_117),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_200),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_171),
.B(n_135),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_187),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_177),
.B(n_171),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_183),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

OR2x2_ASAP7_75t_SL g292 ( 
.A(n_243),
.B(n_196),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_190),
.B(n_237),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_254),
.B(n_274),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_258),
.B(n_221),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_203),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_264),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_209),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_184),
.A2(n_223),
.B1(n_226),
.B2(n_193),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_268),
.A2(n_269),
.B1(n_222),
.B2(n_199),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_218),
.A2(n_192),
.B1(n_208),
.B2(n_235),
.Y(n_269)
);

OAI32xp33_ASAP7_75t_L g271 ( 
.A1(n_238),
.A2(n_189),
.A3(n_194),
.B1(n_213),
.B2(n_182),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_212),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_194),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_278),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_276),
.B(n_277),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_188),
.B(n_198),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_204),
.B(n_211),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_280),
.B(n_284),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_277),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_285),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_220),
.C(n_215),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_299),
.C(n_304),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_259),
.Y(n_285)
);

CKINVDCx12_ASAP7_75t_R g286 ( 
.A(n_262),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_286),
.Y(n_327)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_287),
.Y(n_314)
);

AOI221xp5_ASAP7_75t_L g317 ( 
.A1(n_288),
.A2(n_292),
.B1(n_300),
.B2(n_255),
.C(n_273),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_262),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_289),
.B(n_302),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_202),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_290),
.B(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_206),
.B(n_231),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_253),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_248),
.B(n_234),
.Y(n_297)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_252),
.B(n_257),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_307),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_186),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_243),
.A2(n_254),
.B(n_241),
.Y(n_300)
);

AOI22x1_ASAP7_75t_L g301 ( 
.A1(n_268),
.A2(n_260),
.B1(n_244),
.B2(n_241),
.Y(n_301)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_301),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_278),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_260),
.A2(n_275),
.B1(n_251),
.B2(n_245),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_271),
.B1(n_255),
.B2(n_278),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_245),
.C(n_251),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_257),
.A2(n_252),
.B1(n_242),
.B2(n_244),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_247),
.B1(n_250),
.B2(n_272),
.Y(n_318)
);

NAND2xp33_ASAP7_75t_SL g307 ( 
.A(n_242),
.B(n_247),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_309),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_263),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_324),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_296),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_317),
.B(n_318),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_270),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_323),
.C(n_328),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_270),
.C(n_250),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_281),
.B(n_272),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_256),
.Y(n_325)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_300),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_256),
.Y(n_329)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_329),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_324),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_336),
.Y(n_353)
);

A2O1A1O1Ixp25_ASAP7_75t_L g333 ( 
.A1(n_326),
.A2(n_294),
.B(n_301),
.C(n_292),
.D(n_283),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_333),
.A2(n_341),
.B(n_347),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_330),
.A2(n_295),
.B(n_312),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_334),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_311),
.Y(n_336)
);

OA22x2_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_302),
.B1(n_301),
.B2(n_280),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_337),
.B(n_340),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_338),
.B(n_321),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_313),
.A2(n_295),
.B(n_296),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_339),
.B(n_342),
.Y(n_354)
);

NOR2x1_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_296),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_310),
.A2(n_293),
.B(n_307),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_315),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_343),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_285),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_322),
.C(n_319),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_351),
.C(n_357),
.Y(n_361)
);

AOI221xp5_ASAP7_75t_L g350 ( 
.A1(n_334),
.A2(n_325),
.B1(n_284),
.B2(n_329),
.C(n_328),
.Y(n_350)
);

NOR3xp33_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_345),
.C(n_340),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_322),
.C(n_310),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_335),
.A2(n_323),
.B1(n_305),
.B2(n_321),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_355),
.A2(n_332),
.B1(n_344),
.B2(n_331),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_282),
.C(n_327),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_336),
.A2(n_327),
.B(n_314),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_342),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_359),
.B(n_335),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_354),
.Y(n_362)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_362),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_332),
.C(n_338),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_370),
.C(n_359),
.Y(n_376)
);

XOR2x2_ASAP7_75t_SL g372 ( 
.A(n_364),
.B(n_365),
.Y(n_372)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_353),
.Y(n_366)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_366),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_367),
.B(n_368),
.Y(n_373)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_356),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_356),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_362),
.C(n_363),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_364),
.A2(n_360),
.B(n_352),
.C(n_339),
.Y(n_371)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_371),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_376),
.B(n_361),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_361),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_378),
.B(n_380),
.Y(n_384)
);

OAI21x1_ASAP7_75t_SL g379 ( 
.A1(n_374),
.A2(n_341),
.B(n_340),
.Y(n_379)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_379),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_348),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_372),
.C(n_351),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_383),
.B(n_381),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_387),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_384),
.B(n_375),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_386),
.A2(n_381),
.B(n_385),
.Y(n_388)
);

OAI32xp33_ASAP7_75t_L g390 ( 
.A1(n_388),
.A2(n_371),
.A3(n_372),
.B1(n_344),
.B2(n_314),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_389),
.Y(n_391)
);


endmodule