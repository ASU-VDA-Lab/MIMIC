module fake_jpeg_20926_n_107 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx8_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_25),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_14),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_26),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_17),
.B1(n_19),
.B2(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_27),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_19),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_0),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_26),
.B1(n_22),
.B2(n_21),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_46),
.B1(n_51),
.B2(n_14),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_25),
.B1(n_21),
.B2(n_27),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_48),
.B1(n_34),
.B2(n_25),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_25),
.Y(n_60)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_20),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_36),
.B1(n_33),
.B2(n_30),
.Y(n_54)
);

AO21x2_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_24),
.B(n_52),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_56),
.B1(n_50),
.B2(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_64),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_16),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_65),
.C(n_11),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_16),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_20),
.C(n_10),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_70),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_51),
.B1(n_48),
.B2(n_47),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_74),
.B(n_61),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_81),
.Y(n_91)
);

AO221x1_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_2),
.B1(n_3),
.B2(n_24),
.C(n_7),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_66),
.B1(n_74),
.B2(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_88),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_75),
.C(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_90),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_2),
.Y(n_103)
);

NOR2xp67_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_98),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_83),
.A3(n_89),
.B1(n_93),
.B2(n_65),
.C1(n_18),
.C2(n_8),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_18),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_103),
.C(n_8),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_83),
.B(n_5),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_100),
.C(n_105),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g107 ( 
.A(n_106),
.Y(n_107)
);


endmodule