module fake_jpeg_7156_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_37),
.A2(n_54),
.B1(n_26),
.B2(n_28),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_39),
.B(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_21),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_16),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_57),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_0),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_17),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_51),
.Y(n_66)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_2),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_59),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_24),
.Y(n_56)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_11),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_71),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_36),
.B1(n_31),
.B2(n_30),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_70),
.B1(n_83),
.B2(n_34),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_26),
.B1(n_36),
.B2(n_30),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_65),
.B(n_87),
.C(n_34),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_37),
.A2(n_36),
.B1(n_31),
.B2(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_86),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_51),
.B1(n_25),
.B2(n_18),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_90),
.B1(n_77),
.B2(n_82),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_84),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_35),
.B1(n_32),
.B2(n_20),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_15),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_33),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_17),
.B1(n_32),
.B2(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_89),
.Y(n_121)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_41),
.A2(n_33),
.B1(n_17),
.B2(n_35),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_33),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_76),
.Y(n_108)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_100),
.Y(n_127)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_72),
.B(n_89),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_33),
.B1(n_34),
.B2(n_32),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_68),
.B1(n_73),
.B2(n_8),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_108),
.Y(n_130)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_5),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_113),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_124),
.B1(n_20),
.B2(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_65),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

AO21x2_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_116),
.B(n_124),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_131),
.B1(n_142),
.B2(n_111),
.Y(n_152)
);

OR2x4_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_88),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_113),
.B(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_91),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_139),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_95),
.B1(n_94),
.B2(n_82),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_97),
.B1(n_100),
.B2(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_147),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_91),
.C(n_69),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_138),
.C(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_67),
.C(n_92),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_73),
.B1(n_68),
.B2(n_11),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_5),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_9),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_6),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_118),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_6),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_10),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_146),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_151),
.Y(n_174)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_126),
.B1(n_131),
.B2(n_129),
.C(n_139),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_157),
.B(n_127),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_135),
.C(n_138),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_162),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_159),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_128),
.B(n_112),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_117),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_167),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_106),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_128),
.B(n_9),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_173),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_102),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_154),
.C(n_134),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_132),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_183),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_162),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_185),
.A2(n_189),
.B(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_125),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_190),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_192),
.A2(n_195),
.B1(n_198),
.B2(n_204),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_163),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_165),
.B1(n_126),
.B2(n_153),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_165),
.B1(n_126),
.B2(n_153),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_126),
.B1(n_171),
.B2(n_164),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_199),
.A2(n_200),
.B1(n_180),
.B2(n_144),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_171),
.B1(n_125),
.B2(n_159),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_205),
.C(n_186),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_203),
.B(n_177),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_159),
.B1(n_154),
.B2(n_158),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_130),
.C(n_142),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_208),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_211),
.C(n_213),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_189),
.C(n_175),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_173),
.B(n_176),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_204),
.B(n_202),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_192),
.B(n_176),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_175),
.B1(n_174),
.B2(n_180),
.Y(n_214)
);

NAND4xp25_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_215),
.C(n_195),
.D(n_198),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_209),
.A2(n_197),
.B1(n_202),
.B2(n_196),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_217),
.A2(n_205),
.B(n_200),
.Y(n_226)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_191),
.C(n_151),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_196),
.C(n_194),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_211),
.C(n_213),
.Y(n_224)
);

OAI31xp33_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_160),
.A3(n_173),
.B(n_150),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_226),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_229),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_228),
.A2(n_218),
.B1(n_216),
.B2(n_147),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_160),
.C(n_168),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_221),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_234),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_219),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_224),
.B(n_222),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_237),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_231),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_232),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_239),
.Y(n_241)
);


endmodule