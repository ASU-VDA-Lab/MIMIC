module fake_jpeg_18692_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_15),
.B(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_55),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_67),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_43),
.B1(n_38),
.B2(n_48),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_45),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_41),
.B(n_43),
.C(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_50),
.B1(n_39),
.B2(n_2),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_64),
.B1(n_71),
.B2(n_6),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_7),
.Y(n_92)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_83),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_70),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_71),
.B1(n_64),
.B2(n_5),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_89),
.B1(n_90),
.B2(n_88),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_96),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_74),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_76),
.B(n_72),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_96),
.B(n_94),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_72),
.B1(n_82),
.B2(n_14),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_98),
.B(n_9),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_SL g103 ( 
.A(n_99),
.B(n_10),
.C(n_16),
.Y(n_103)
);

OAI322xp33_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_86),
.A3(n_93),
.B1(n_19),
.B2(n_20),
.C1(n_22),
.C2(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_101),
.C(n_26),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_103),
.B1(n_27),
.B2(n_29),
.Y(n_106)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_107)
);

AOI21x1_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_33),
.B(n_34),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_35),
.B(n_36),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_86),
.Y(n_111)
);


endmodule