module fake_jpeg_14817_n_121 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_0),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_1),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_74),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_60),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_64),
.B1(n_63),
.B2(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_80),
.Y(n_95)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_64),
.B1(n_46),
.B2(n_62),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_86),
.B(n_2),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_68),
.A2(n_46),
.B1(n_61),
.B2(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_4),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_92),
.B(n_94),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_2),
.B(n_3),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_93),
.B(n_6),
.C(n_60),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_58),
.B(n_57),
.C(n_49),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_48),
.B(n_27),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_6),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_99),
.Y(n_103)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_78),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_95),
.B1(n_96),
.B2(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_104),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_76),
.B1(n_83),
.B2(n_81),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_101),
.B(n_104),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_88),
.Y(n_110)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_105),
.B(n_53),
.CI(n_10),
.CON(n_108),
.SN(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_8),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_110),
.B1(n_108),
.B2(n_106),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_111),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_14),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_16),
.C(n_17),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_19),
.C(n_21),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_22),
.A3(n_25),
.B1(n_26),
.B2(n_31),
.C1(n_32),
.C2(n_33),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_34),
.Y(n_118)
);

AOI321xp33_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_35),
.A3(n_37),
.B1(n_38),
.B2(n_40),
.C(n_43),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_44),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_45),
.Y(n_121)
);


endmodule