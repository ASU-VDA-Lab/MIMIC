module real_aes_656_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_204;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g96 ( .A1(n_0), .A2(n_55), .B1(n_93), .B2(n_97), .Y(n_96) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_1), .A2(n_14), .B1(n_113), .B2(n_117), .Y(n_112) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_2), .A2(n_35), .B1(n_123), .B2(n_127), .Y(n_122) );
INVx1_ASAP7_75t_L g196 ( .A(n_3), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g86 ( .A1(n_4), .A2(n_72), .B1(n_87), .B2(n_107), .Y(n_86) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_5), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g267 ( .A(n_6), .Y(n_267) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_7), .A2(n_20), .B1(n_93), .B2(n_94), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_8), .Y(n_237) );
INVx2_ASAP7_75t_L g214 ( .A(n_9), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_10), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_174) );
INVx1_ASAP7_75t_L g176 ( .A(n_10), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_11), .A2(n_63), .B1(n_131), .B2(n_134), .Y(n_130) );
INVx1_ASAP7_75t_L g292 ( .A(n_12), .Y(n_292) );
INVx1_ASAP7_75t_SL g279 ( .A(n_13), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_15), .B(n_225), .Y(n_336) );
OAI22xp5_ASAP7_75t_SL g179 ( .A1(n_16), .A2(n_180), .B1(n_183), .B2(n_184), .Y(n_179) );
INVx1_ASAP7_75t_L g184 ( .A(n_16), .Y(n_184) );
AOI33xp33_ASAP7_75t_L g316 ( .A1(n_17), .A2(n_40), .A3(n_218), .B1(n_241), .B2(n_317), .B3(n_318), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_18), .A2(n_43), .B1(n_160), .B2(n_164), .Y(n_159) );
INVx1_ASAP7_75t_L g223 ( .A(n_19), .Y(n_223) );
OAI221xp5_ASAP7_75t_L g188 ( .A1(n_20), .A2(n_55), .B1(n_58), .B2(n_189), .C(n_191), .Y(n_188) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_21), .A2(n_68), .B(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g261 ( .A(n_21), .B(n_68), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_22), .B(n_245), .Y(n_276) );
INVx3_ASAP7_75t_L g93 ( .A(n_23), .Y(n_93) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_24), .A2(n_25), .B1(n_151), .B2(n_154), .Y(n_150) );
INVx1_ASAP7_75t_SL g102 ( .A(n_26), .Y(n_102) );
INVx1_ASAP7_75t_L g198 ( .A(n_27), .Y(n_198) );
AND2x2_ASAP7_75t_L g231 ( .A(n_27), .B(n_196), .Y(n_231) );
AND2x2_ASAP7_75t_L g248 ( .A(n_27), .B(n_221), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_28), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_29), .B(n_245), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_30), .A2(n_212), .B1(n_286), .B2(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_31), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_32), .B(n_225), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_33), .A2(n_70), .B1(n_181), .B2(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_33), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_34), .A2(n_81), .B1(n_82), .B2(n_169), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g169 ( .A(n_34), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_36), .B(n_264), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_37), .B(n_225), .Y(n_268) );
AO22x2_ASAP7_75t_L g105 ( .A1(n_38), .A2(n_58), .B1(n_93), .B2(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_39), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_41), .B(n_225), .Y(n_256) );
INVx1_ASAP7_75t_L g219 ( .A(n_42), .Y(n_219) );
INVx1_ASAP7_75t_L g227 ( .A(n_42), .Y(n_227) );
AND2x2_ASAP7_75t_L g258 ( .A(n_44), .B(n_259), .Y(n_258) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_45), .A2(n_59), .B1(n_239), .B2(n_245), .C(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_46), .B(n_245), .Y(n_307) );
INVx1_ASAP7_75t_L g103 ( .A(n_47), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_48), .A2(n_81), .B1(n_82), .B2(n_578), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_48), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_49), .B(n_212), .Y(n_243) );
AOI21xp5_ASAP7_75t_SL g303 ( .A1(n_50), .A2(n_239), .B(n_304), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_50), .A2(n_81), .B1(n_82), .B2(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_50), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_51), .A2(n_67), .B1(n_143), .B2(n_146), .Y(n_142) );
INVx1_ASAP7_75t_L g289 ( .A(n_52), .Y(n_289) );
INVx1_ASAP7_75t_L g255 ( .A(n_53), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_54), .A2(n_239), .B(n_254), .Y(n_253) );
INVxp33_ASAP7_75t_L g193 ( .A(n_55), .Y(n_193) );
INVx1_ASAP7_75t_L g221 ( .A(n_56), .Y(n_221) );
INVx1_ASAP7_75t_L g229 ( .A(n_56), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_57), .B(n_245), .Y(n_319) );
INVxp67_ASAP7_75t_L g192 ( .A(n_58), .Y(n_192) );
INVx1_ASAP7_75t_L g175 ( .A(n_59), .Y(n_175) );
AND2x2_ASAP7_75t_L g281 ( .A(n_60), .B(n_211), .Y(n_281) );
INVx1_ASAP7_75t_L g290 ( .A(n_61), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_62), .A2(n_239), .B(n_278), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_64), .A2(n_239), .B(n_311), .C(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_SL g301 ( .A(n_65), .B(n_211), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_66), .A2(n_239), .B1(n_314), .B2(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_69), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g182 ( .A(n_70), .Y(n_182) );
INVx1_ASAP7_75t_L g305 ( .A(n_71), .Y(n_305) );
INVx1_ASAP7_75t_L g171 ( .A(n_73), .Y(n_171) );
AND2x2_ASAP7_75t_L g320 ( .A(n_74), .B(n_211), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_75), .A2(n_216), .B(n_222), .C(n_230), .Y(n_215) );
BUFx2_ASAP7_75t_SL g190 ( .A(n_76), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_77), .B(n_225), .Y(n_306) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_185), .B1(n_199), .B2(n_565), .C(n_568), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_170), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NOR2xp33_ASAP7_75t_L g84 ( .A(n_85), .B(n_136), .Y(n_84) );
NAND4xp25_ASAP7_75t_SL g85 ( .A(n_86), .B(n_112), .C(n_122), .D(n_130), .Y(n_85) );
INVx4_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx8_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x4_ASAP7_75t_L g89 ( .A(n_90), .B(n_98), .Y(n_89) );
AND2x2_ASAP7_75t_L g115 ( .A(n_90), .B(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g132 ( .A(n_90), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g140 ( .A(n_90), .B(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g90 ( .A(n_91), .B(n_95), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x4_ASAP7_75t_L g111 ( .A(n_92), .B(n_95), .Y(n_111) );
INVx1_ASAP7_75t_L g121 ( .A(n_92), .Y(n_121) );
AND2x2_ASAP7_75t_L g129 ( .A(n_92), .B(n_96), .Y(n_129) );
INVx2_ASAP7_75t_L g94 ( .A(n_93), .Y(n_94) );
INVx1_ASAP7_75t_L g97 ( .A(n_93), .Y(n_97) );
OAI22x1_ASAP7_75t_L g100 ( .A1(n_93), .A2(n_101), .B1(n_102), .B2(n_103), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_93), .Y(n_101) );
INVx1_ASAP7_75t_L g106 ( .A(n_93), .Y(n_106) );
INVxp67_ASAP7_75t_L g149 ( .A(n_95), .Y(n_149) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g120 ( .A(n_96), .B(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g110 ( .A(n_98), .B(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g119 ( .A(n_98), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g135 ( .A(n_98), .B(n_129), .Y(n_135) );
AND2x4_ASAP7_75t_L g98 ( .A(n_99), .B(n_104), .Y(n_98) );
AND2x2_ASAP7_75t_L g116 ( .A(n_99), .B(n_105), .Y(n_116) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g133 ( .A(n_100), .B(n_104), .Y(n_133) );
AND2x2_ASAP7_75t_L g141 ( .A(n_100), .B(n_105), .Y(n_141) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_100), .Y(n_158) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_L g128 ( .A(n_105), .Y(n_128) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g145 ( .A(n_111), .B(n_116), .Y(n_145) );
AND2x2_ASAP7_75t_L g153 ( .A(n_111), .B(n_133), .Y(n_153) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g126 ( .A(n_116), .B(n_120), .Y(n_126) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx8_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g163 ( .A(n_120), .B(n_133), .Y(n_163) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_121), .Y(n_168) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x2_ASAP7_75t_L g157 ( .A(n_129), .B(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx2_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
NAND4xp25_ASAP7_75t_SL g136 ( .A(n_137), .B(n_142), .C(n_150), .D(n_159), .Y(n_136) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx6_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g148 ( .A(n_141), .B(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g166 ( .A(n_141), .B(n_167), .Y(n_166) );
BUFx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx6_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
XOR2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B1(n_178), .B2(n_179), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_SL g177 ( .A(n_175), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_176), .A2(n_292), .B1(n_293), .B2(n_295), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_180), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
AND3x1_ASAP7_75t_SL g187 ( .A(n_188), .B(n_194), .C(n_197), .Y(n_187) );
INVxp67_ASAP7_75t_L g576 ( .A(n_188), .Y(n_576) );
CKINVDCx8_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g574 ( .A(n_194), .Y(n_574) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_194), .A2(n_331), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g246 ( .A(n_195), .B(n_218), .Y(n_246) );
OR2x2_ASAP7_75t_SL g581 ( .A(n_195), .B(n_197), .Y(n_581) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g242 ( .A(n_196), .B(n_219), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_197), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2x1p5_ASAP7_75t_L g240 ( .A(n_198), .B(n_241), .Y(n_240) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND3x1_ASAP7_75t_L g202 ( .A(n_203), .B(n_444), .C(n_511), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_404), .Y(n_203) );
NOR3x1_ASAP7_75t_L g204 ( .A(n_205), .B(n_355), .C(n_384), .Y(n_204) );
OAI221xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_270), .B1(n_308), .B2(n_323), .C(n_340), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_SL g518 ( .A1(n_206), .A2(n_283), .B(n_519), .C(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_207), .A2(n_490), .B1(n_493), .B2(n_495), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_207), .B(n_309), .Y(n_564) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_249), .Y(n_207) );
BUFx2_ASAP7_75t_L g483 ( .A(n_208), .Y(n_483) );
INVx1_ASAP7_75t_SL g496 ( .A(n_208), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_208), .B(n_351), .Y(n_538) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x4_ASAP7_75t_L g321 ( .A(n_209), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g366 ( .A(n_209), .B(n_263), .Y(n_366) );
INVx1_ASAP7_75t_L g377 ( .A(n_209), .Y(n_377) );
INVx2_ASAP7_75t_L g381 ( .A(n_209), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_209), .B(n_352), .Y(n_508) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_234), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_215), .B1(n_232), .B2(n_233), .Y(n_210) );
INVx3_ASAP7_75t_L g233 ( .A(n_211), .Y(n_233) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_212), .B(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
BUFx4f_ASAP7_75t_L g264 ( .A(n_213), .Y(n_264) );
AND2x2_ASAP7_75t_SL g260 ( .A(n_214), .B(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g286 ( .A(n_214), .B(n_261), .Y(n_286) );
INVxp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_217), .A2(n_255), .B(n_256), .C(n_257), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g266 ( .A1(n_217), .A2(n_257), .B(n_267), .C(n_268), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_SL g278 ( .A1(n_217), .A2(n_257), .B(n_279), .C(n_280), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_217), .A2(n_224), .B1(n_289), .B2(n_290), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_217), .A2(n_257), .B(n_305), .C(n_306), .Y(n_304) );
INVx2_ASAP7_75t_L g338 ( .A(n_217), .Y(n_338) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
INVxp33_ASAP7_75t_L g317 ( .A(n_218), .Y(n_317) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x4_ASAP7_75t_L g296 ( .A(n_219), .B(n_228), .Y(n_296) );
INVx3_ASAP7_75t_L g241 ( .A(n_220), .Y(n_241) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x6_ASAP7_75t_L g294 ( .A(n_221), .B(n_226), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_228), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx5_ASAP7_75t_L g257 ( .A(n_231), .Y(n_257) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_233), .A2(n_251), .B(n_258), .Y(n_250) );
AO21x2_ASAP7_75t_L g352 ( .A1(n_233), .A2(n_251), .B(n_258), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_238), .B1(n_243), .B2(n_244), .Y(n_234) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVxp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
INVx1_ASAP7_75t_L g318 ( .A(n_241), .Y(n_318) );
AND2x6_ASAP7_75t_L g567 ( .A(n_242), .B(n_248), .Y(n_567) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g331 ( .A(n_246), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_247), .Y(n_332) );
BUFx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g457 ( .A(n_249), .B(n_458), .Y(n_457) );
NOR2x1_ASAP7_75t_L g249 ( .A(n_250), .B(n_262), .Y(n_249) );
INVx2_ASAP7_75t_L g360 ( .A(n_250), .Y(n_360) );
AND2x2_ASAP7_75t_L g380 ( .A(n_250), .B(n_381), .Y(n_380) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_250), .B(n_381), .Y(n_505) );
AND2x2_ASAP7_75t_L g530 ( .A(n_250), .B(n_373), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_257), .B(n_286), .Y(n_297) );
INVx1_ASAP7_75t_L g314 ( .A(n_257), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_257), .A2(n_336), .B(n_337), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_259), .Y(n_274) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g322 ( .A(n_263), .Y(n_322) );
INVx1_ASAP7_75t_L g344 ( .A(n_263), .Y(n_344) );
INVxp67_ASAP7_75t_L g383 ( .A(n_263), .Y(n_383) );
AND2x4_ASAP7_75t_L g423 ( .A(n_263), .B(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_263), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_263), .B(n_374), .Y(n_509) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B(n_269), .Y(n_263) );
INVx2_ASAP7_75t_SL g311 ( .A(n_264), .Y(n_311) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_282), .Y(n_271) );
AND2x2_ASAP7_75t_L g397 ( .A(n_272), .B(n_369), .Y(n_397) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_273), .Y(n_325) );
AND2x2_ASAP7_75t_L g353 ( .A(n_273), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g364 ( .A(n_273), .Y(n_364) );
INVx1_ASAP7_75t_L g388 ( .A(n_273), .Y(n_388) );
AND2x2_ASAP7_75t_L g391 ( .A(n_273), .B(n_284), .Y(n_391) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_273), .Y(n_413) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_275), .B(n_281), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NOR2x1_ASAP7_75t_L g282 ( .A(n_283), .B(n_298), .Y(n_282) );
AND2x2_ASAP7_75t_L g378 ( .A(n_283), .B(n_300), .Y(n_378) );
NAND2x1_ASAP7_75t_L g411 ( .A(n_283), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g514 ( .A(n_283), .Y(n_514) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g354 ( .A(n_284), .Y(n_354) );
AND2x2_ASAP7_75t_L g369 ( .A(n_284), .B(n_328), .Y(n_369) );
NOR2x1_ASAP7_75t_SL g438 ( .A(n_284), .B(n_300), .Y(n_438) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_286), .A2(n_303), .B(n_307), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_291), .B(n_297), .Y(n_287) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NOR2x1_ASAP7_75t_L g475 ( .A(n_298), .B(n_462), .Y(n_475) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g400 ( .A(n_299), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx4_ASAP7_75t_L g339 ( .A(n_300), .Y(n_339) );
AND2x4_ASAP7_75t_L g346 ( .A(n_300), .B(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_300), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_300), .B(n_363), .Y(n_463) );
AND2x2_ASAP7_75t_L g491 ( .A(n_300), .B(n_328), .Y(n_491) );
OR2x6_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
OAI222xp33_ASAP7_75t_L g568 ( .A1(n_305), .A2(n_569), .B1(n_571), .B2(n_577), .C1(n_579), .C2(n_582), .Y(n_568) );
NAND2x1_ASAP7_75t_SL g308 ( .A(n_309), .B(n_321), .Y(n_308) );
OR2x2_ASAP7_75t_L g519 ( .A(n_309), .B(n_431), .Y(n_519) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g359 ( .A(n_310), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g424 ( .A(n_310), .Y(n_424) );
AND2x2_ASAP7_75t_L g458 ( .A(n_310), .B(n_381), .Y(n_458) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_320), .Y(n_310) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_311), .A2(n_312), .B(n_320), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_313), .B(n_319), .Y(n_312) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g431 ( .A(n_321), .Y(n_431) );
AND2x2_ASAP7_75t_L g439 ( .A(n_321), .B(n_372), .Y(n_439) );
AND2x2_ASAP7_75t_L g556 ( .A(n_321), .B(n_359), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g510 ( .A(n_325), .B(n_451), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_325), .B(n_350), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_326), .A2(n_387), .B(n_390), .Y(n_386) );
AND2x2_ASAP7_75t_L g456 ( .A(n_326), .B(n_362), .Y(n_456) );
INVx2_ASAP7_75t_SL g543 ( .A(n_326), .Y(n_543) );
AND2x4_ASAP7_75t_SL g326 ( .A(n_327), .B(n_339), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g347 ( .A(n_328), .Y(n_347) );
INVx2_ASAP7_75t_L g394 ( .A(n_328), .Y(n_394) );
AND2x4_ASAP7_75t_L g401 ( .A(n_328), .B(n_354), .Y(n_401) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_334), .Y(n_328) );
NOR3xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .C(n_333), .Y(n_330) );
INVxp67_ASAP7_75t_L g584 ( .A(n_332), .Y(n_584) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_339), .Y(n_357) );
AND2x4_ASAP7_75t_L g433 ( .A(n_339), .B(n_347), .Y(n_433) );
OR2x2_ASAP7_75t_L g559 ( .A(n_339), .B(n_560), .Y(n_559) );
NAND4xp25_ASAP7_75t_L g340 ( .A(n_341), .B(n_345), .C(n_348), .D(n_353), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g406 ( .A(n_342), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g503 ( .A(n_342), .Y(n_503) );
INVx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_343), .B(n_351), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_343), .B(n_408), .Y(n_537) );
BUFx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_346), .B(n_362), .Y(n_415) );
INVx2_ASAP7_75t_L g517 ( .A(n_346), .Y(n_517) );
AND2x2_ASAP7_75t_SL g527 ( .A(n_346), .B(n_387), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_346), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g419 ( .A(n_350), .B(n_366), .Y(n_419) );
AND2x2_ASAP7_75t_L g487 ( .A(n_350), .B(n_423), .Y(n_487) );
INVx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g372 ( .A(n_351), .B(n_373), .Y(n_372) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_352), .Y(n_426) );
AND2x2_ASAP7_75t_L g477 ( .A(n_352), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_352), .B(n_374), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_353), .B(n_517), .Y(n_524) );
INVx1_ASAP7_75t_SL g560 ( .A(n_353), .Y(n_560) );
INVx1_ASAP7_75t_L g389 ( .A(n_354), .Y(n_389) );
AND2x2_ASAP7_75t_L g451 ( .A(n_354), .B(n_394), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_365), .B(n_367), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
AND2x2_ASAP7_75t_L g417 ( .A(n_359), .B(n_366), .Y(n_417) );
AND2x2_ASAP7_75t_L g525 ( .A(n_359), .B(n_376), .Y(n_525) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g399 ( .A(n_362), .Y(n_399) );
AND2x2_ASAP7_75t_L g432 ( .A(n_362), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g437 ( .A(n_362), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_362), .B(n_401), .Y(n_486) );
NOR3xp33_ASAP7_75t_L g536 ( .A(n_362), .B(n_537), .C(n_538), .Y(n_536) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B1(n_378), .B2(n_379), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx2_ASAP7_75t_L g462 ( .A(n_369), .Y(n_462) );
AND2x2_ASAP7_75t_L g396 ( .A(n_370), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g418 ( .A(n_370), .B(n_391), .Y(n_418) );
AND2x2_ASAP7_75t_SL g450 ( .A(n_370), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_375), .Y(n_371) );
INVx1_ASAP7_75t_L g429 ( .A(n_372), .Y(n_429) );
AND2x2_ASAP7_75t_L g382 ( .A(n_373), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g408 ( .A(n_373), .Y(n_408) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g471 ( .A(n_377), .B(n_423), .Y(n_471) );
INVx1_ASAP7_75t_L g529 ( .A(n_377), .Y(n_529) );
INVx1_ASAP7_75t_L g385 ( .A(n_379), .Y(n_385) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_380), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g516 ( .A(n_380), .B(n_423), .Y(n_516) );
AND2x2_ASAP7_75t_L g482 ( .A(n_382), .B(n_483), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g550 ( .A(n_382), .B(n_551), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B(n_395), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_387), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g443 ( .A(n_387), .B(n_392), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_387), .B(n_433), .Y(n_494) );
AND2x4_ASAP7_75t_SL g387 ( .A(n_388), .B(n_389), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_388), .B(n_451), .Y(n_481) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_388), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_390), .A2(n_417), .B1(n_418), .B2(n_419), .Y(n_416) );
AND2x2_ASAP7_75t_SL g390 ( .A(n_391), .B(n_392), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_391), .B(n_433), .Y(n_452) );
INVx1_ASAP7_75t_L g553 ( .A(n_391), .Y(n_553) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B(n_402), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_397), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g534 ( .A(n_400), .Y(n_534) );
INVx4_ASAP7_75t_L g436 ( .A(n_401), .Y(n_436) );
INVxp33_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g464 ( .A(n_403), .B(n_465), .Y(n_464) );
NOR2x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_420), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B(n_416), .Y(n_405) );
INVx1_ASAP7_75t_L g454 ( .A(n_407), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g459 ( .A(n_411), .Y(n_459) );
INVx1_ASAP7_75t_L g492 ( .A(n_412), .Y(n_492) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_417), .A2(n_456), .B1(n_457), .B2(n_459), .Y(n_455) );
INVx1_ASAP7_75t_L g469 ( .A(n_418), .Y(n_469) );
NAND4xp25_ASAP7_75t_SL g420 ( .A(n_421), .B(n_427), .C(n_434), .D(n_440), .Y(n_420) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g442 ( .A(n_423), .Y(n_442) );
AND2x2_ASAP7_75t_L g554 ( .A(n_423), .B(n_551), .Y(n_554) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g561 ( .A(n_431), .B(n_498), .Y(n_561) );
INVx1_ASAP7_75t_L g558 ( .A(n_432), .Y(n_558) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_433), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B(n_439), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_472), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_460), .C(n_468), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_453), .B(n_455), .Y(n_446) );
INVxp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_452), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_450), .A2(n_482), .B1(n_485), .B2(n_487), .Y(n_484) );
OAI22xp33_ASAP7_75t_L g460 ( .A1(n_453), .A2(n_461), .B1(n_464), .B2(n_466), .Y(n_460) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g465 ( .A(n_458), .Y(n_465) );
AND2x4_ASAP7_75t_L g476 ( .A(n_458), .B(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_463), .Y(n_563) );
AOI31xp33_ASAP7_75t_L g562 ( .A1(n_466), .A2(n_539), .A3(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_488), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_474), .B(n_484), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_479), .B2(n_482), .Y(n_474) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_478), .Y(n_542) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_486), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_489), .B(n_499), .Y(n_488) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AND2x2_ASAP7_75t_L g500 ( .A(n_491), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g539 ( .A(n_491), .Y(n_539) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_491), .A2(n_549), .B1(n_552), .B2(n_554), .Y(n_548) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_496), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_502), .B1(n_506), .B2(n_510), .Y(n_499) );
NOR2xp33_ASAP7_75t_SL g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVxp67_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_SL g551 ( .A(n_508), .Y(n_551) );
INVx2_ASAP7_75t_L g532 ( .A(n_509), .Y(n_532) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_546), .Y(n_511) );
AOI211xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_518), .B(n_521), .C(n_535), .Y(n_512) );
OAI21xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_517), .Y(n_513) );
INVx1_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g520 ( .A(n_517), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_522), .B(n_526), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B1(n_531), .B2(n_533), .Y(n_526) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
AND2x2_ASAP7_75t_L g531 ( .A(n_529), .B(n_532), .Y(n_531) );
AO22x1_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_539), .B1(n_540), .B2(n_544), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_557), .C(n_562), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_548), .B(n_555), .Y(n_547) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI21xp33_ASAP7_75t_R g557 ( .A1(n_558), .A2(n_559), .B(n_561), .Y(n_557) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_572), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_583), .Y(n_582) );
endmodule