module fake_jpeg_250_n_189 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_189);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_12),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_72),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_71),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_47),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_49),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_64),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_56),
.B1(n_51),
.B2(n_59),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_86),
.B1(n_88),
.B2(n_52),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_89),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_74),
.B1(n_56),
.B2(n_51),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_59),
.B1(n_64),
.B2(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_4),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_54),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_104),
.C(n_5),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_62),
.B(n_58),
.C(n_57),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_63),
.B1(n_55),
.B2(n_52),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_105),
.B1(n_22),
.B2(n_45),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_63),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_55),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_1),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_108),
.B(n_114),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_1),
.B(n_2),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_26),
.B(n_30),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_3),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_24),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_129)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_123),
.Y(n_147)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_99),
.C(n_102),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_132),
.C(n_118),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_129),
.B1(n_136),
.B2(n_139),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_27),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_29),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_135),
.Y(n_154)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_12),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_137),
.B(n_141),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_18),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_138),
.B(n_36),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_142),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_21),
.B(n_25),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_38),
.B(n_41),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_32),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_147),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_107),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_156),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_122),
.B(n_34),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_35),
.Y(n_158)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_161),
.B(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_37),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_164),
.B1(n_144),
.B2(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_128),
.B1(n_164),
.B2(n_160),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_172),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g172 ( 
.A1(n_150),
.A2(n_160),
.B1(n_153),
.B2(n_139),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_149),
.C(n_132),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_174),
.B(n_176),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_155),
.B1(n_145),
.B2(n_136),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_170),
.A2(n_156),
.B(n_154),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_167),
.B(n_169),
.Y(n_181)
);

OAI21x1_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_168),
.B(n_172),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_173),
.B1(n_172),
.B2(n_133),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_145),
.C(n_162),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_181),
.C(n_143),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_182),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_178),
.C(n_183),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_129),
.C(n_42),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_46),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);


endmodule