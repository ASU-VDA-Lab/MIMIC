module fake_jpeg_16062_n_69 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_69);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_43;
wire n_29;
wire n_50;
wire n_37;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_8),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_0),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_22),
.Y(n_29)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_2),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_2),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_17),
.B1(n_9),
.B2(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_3),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_22),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_17),
.B(n_12),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_26),
.B(n_19),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_21),
.A2(n_11),
.B1(n_12),
.B2(n_18),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_14),
.B(n_16),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_16),
.B(n_13),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_14),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_13),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_7),
.C(n_32),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_47),
.Y(n_54)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_6),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_50),
.C(n_31),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_31),
.B(n_39),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_56),
.C(n_57),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_29),
.C(n_30),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_40),
.C(n_33),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_48),
.C(n_46),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_51),
.C(n_37),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_47),
.B(n_42),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_61),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_45),
.B(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_65),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_58),
.B1(n_64),
.B2(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_66),
.Y(n_69)
);


endmodule