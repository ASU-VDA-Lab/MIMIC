module fake_jpeg_867_n_111 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_33),
.B1(n_34),
.B2(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_35),
.Y(n_48)
);

NAND2x1_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_51),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_36),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_52),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_31),
.B1(n_39),
.B2(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_54),
.B1(n_30),
.B2(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_34),
.B1(n_44),
.B2(n_38),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_61),
.B1(n_42),
.B2(n_58),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_41),
.B1(n_37),
.B2(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_64),
.Y(n_68)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_50),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_42),
.B(n_43),
.C(n_2),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_74),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_49),
.B(n_52),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_56),
.B(n_16),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_41),
.B1(n_42),
.B2(n_50),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_41),
.B1(n_42),
.B2(n_50),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_0),
.CI(n_1),
.CON(n_73),
.SN(n_73)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_62),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_14),
.B1(n_25),
.B2(n_24),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_3),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_6),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_75),
.B1(n_69),
.B2(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_95),
.Y(n_98)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_75),
.B(n_17),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_96),
.A2(n_77),
.B(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_100),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_91),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_94),
.C(n_89),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_102),
.B(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_87),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_96),
.B(n_88),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_81),
.A3(n_99),
.B1(n_95),
.B2(n_93),
.C1(n_19),
.C2(n_20),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_99),
.A3(n_21),
.B1(n_11),
.B2(n_12),
.C1(n_10),
.C2(n_7),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_12),
.Y(n_111)
);


endmodule