module fake_jpeg_17865_n_362 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_362);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_362;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_44),
.B(n_45),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_52),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_49),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_14),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_29),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_59),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_62),
.Y(n_82)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_13),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_68),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_17),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_4),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_71),
.B(n_115),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_33),
.B1(n_37),
.B2(n_22),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_77),
.B1(n_80),
.B2(n_88),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_37),
.B1(n_20),
.B2(n_22),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_76),
.A2(n_78),
.B1(n_91),
.B2(n_96),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_20),
.B1(n_28),
.B2(n_24),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_60),
.B1(n_39),
.B2(n_46),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_81),
.B(n_95),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_45),
.B(n_54),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_90),
.C(n_103),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_29),
.B1(n_21),
.B2(n_27),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_40),
.B(n_19),
.C(n_27),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_68),
.B1(n_59),
.B2(n_58),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_21),
.B1(n_27),
.B2(n_23),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_99),
.B1(n_100),
.B2(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_19),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_23),
.B1(n_9),
.B2(n_10),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_41),
.A2(n_23),
.B1(n_9),
.B2(n_10),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_101),
.B1(n_96),
.B2(n_81),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_42),
.A2(n_19),
.B1(n_13),
.B2(n_12),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_43),
.A2(n_19),
.B1(n_13),
.B2(n_12),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_48),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_40),
.B(n_1),
.C(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_40),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_106),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_2),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_2),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_3),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

HAxp5_ASAP7_75t_SL g118 ( 
.A(n_67),
.B(n_4),
.CON(n_118),
.SN(n_118)
);

OR2x2_ASAP7_75t_SL g164 ( 
.A(n_118),
.B(n_102),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_63),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_6),
.B1(n_76),
.B2(n_119),
.Y(n_121)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_6),
.Y(n_123)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_6),
.Y(n_127)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

CKINVDCx12_ASAP7_75t_R g133 ( 
.A(n_82),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_164),
.B1(n_137),
.B2(n_167),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_135),
.Y(n_200)
);

OR2x4_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_85),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_170),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_87),
.A2(n_104),
.B1(n_98),
.B2(n_89),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_111),
.B1(n_109),
.B2(n_95),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_142),
.A2(n_161),
.B1(n_169),
.B2(n_157),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_85),
.B(n_117),
.C(n_71),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_143),
.B(n_146),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_105),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_147),
.B(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_103),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_170),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_113),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_87),
.A2(n_104),
.B1(n_86),
.B2(n_98),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

CKINVDCx12_ASAP7_75t_R g159 ( 
.A(n_84),
.Y(n_159)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_92),
.B(n_90),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_160),
.B(n_162),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_74),
.B1(n_94),
.B2(n_108),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_114),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_163),
.B(n_167),
.Y(n_208)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_115),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_117),
.B(n_73),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_168),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_96),
.A2(n_37),
.B1(n_30),
.B2(n_33),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_109),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_177),
.A2(n_194),
.B(n_151),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_150),
.C(n_125),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_190),
.C(n_202),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_184),
.B(n_126),
.Y(n_230)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_186),
.A2(n_188),
.B1(n_199),
.B2(n_175),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_187),
.A2(n_131),
.B(n_155),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_130),
.A2(n_169),
.B1(n_125),
.B2(n_136),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_190),
.A2(n_213),
.B1(n_149),
.B2(n_151),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_142),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_202),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_164),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_124),
.A2(n_122),
.B1(n_148),
.B2(n_134),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_135),
.B1(n_152),
.B2(n_154),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_144),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g205 ( 
.A(n_132),
.B(n_121),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_205),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_141),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_146),
.Y(n_218)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_158),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_132),
.A2(n_121),
.B1(n_129),
.B2(n_165),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_228),
.Y(n_264)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_249),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_219),
.B(n_225),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_140),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_222),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_238),
.B1(n_198),
.B2(n_185),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_135),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_138),
.B(n_149),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_242),
.B(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_138),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_224),
.B(n_226),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_138),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_231),
.C(n_234),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_207),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_232),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_230),
.A2(n_246),
.B(n_248),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_182),
.B(n_191),
.C(n_197),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_172),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_205),
.A2(n_171),
.B1(n_212),
.B2(n_184),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_233),
.A2(n_250),
.B1(n_198),
.B2(n_185),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_194),
.C(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_171),
.A2(n_212),
.B1(n_193),
.B2(n_178),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_173),
.Y(n_240)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_200),
.B(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_200),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_186),
.B(n_204),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_176),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_247),
.A2(n_180),
.B(n_250),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_176),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_174),
.B(n_193),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_188),
.A2(n_199),
.B1(n_211),
.B2(n_175),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_251),
.A2(n_257),
.B1(n_258),
.B2(n_260),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_221),
.A2(n_180),
.B1(n_244),
.B2(n_224),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_223),
.B(n_225),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_251),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_215),
.A2(n_230),
.B1(n_229),
.B2(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_215),
.A2(n_238),
.B1(n_222),
.B2(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_219),
.A2(n_218),
.B(n_220),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_239),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_227),
.B(n_231),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_279),
.C(n_226),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_249),
.A2(n_242),
.B(n_245),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_236),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_240),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_278),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_235),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_234),
.B(n_241),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_287),
.C(n_293),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_232),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_214),
.Y(n_284)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_217),
.Y(n_286)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_216),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_296),
.Y(n_308)
);

BUFx12_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_SL g291 ( 
.A(n_253),
.B(n_243),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_299),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_292),
.A2(n_280),
.B1(n_277),
.B2(n_271),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_279),
.C(n_256),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_252),
.B(n_246),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_301),
.Y(n_312)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_295),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_248),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_297),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_298),
.A2(n_273),
.B(n_275),
.Y(n_316)
);

A2O1A1O1Ixp25_ASAP7_75t_L g299 ( 
.A1(n_253),
.A2(n_256),
.B(n_272),
.C(n_266),
.D(n_267),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_265),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_277),
.Y(n_301)
);

INVx13_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_304),
.Y(n_321)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_303),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_268),
.B(n_260),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_309),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_310),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_281),
.A2(n_261),
.B1(n_273),
.B2(n_257),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_311),
.A2(n_319),
.B1(n_285),
.B2(n_300),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_316),
.A2(n_314),
.B(n_310),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_298),
.A2(n_261),
.B1(n_262),
.B2(n_255),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_262),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_322),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_288),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_324),
.Y(n_345)
);

XNOR2x1_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_299),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_326),
.B(n_330),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_287),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_313),
.A2(n_302),
.B1(n_304),
.B2(n_298),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_293),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_319),
.A2(n_305),
.B1(n_286),
.B2(n_291),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_332),
.A2(n_333),
.B(n_314),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_313),
.A2(n_315),
.B1(n_322),
.B2(n_321),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_307),
.B(n_289),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_312),
.Y(n_339)
);

AOI31xp33_ASAP7_75t_L g336 ( 
.A1(n_315),
.A2(n_255),
.A3(n_282),
.B(n_269),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_337),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_339),
.B(n_343),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_323),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_344),
.C(n_328),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_332),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_326),
.B(n_290),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_323),
.Y(n_344)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_346),
.Y(n_354)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_348),
.B(n_349),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_327),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_350),
.A2(n_306),
.B1(n_317),
.B2(n_329),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_331),
.C(n_324),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_351),
.A2(n_335),
.B1(n_325),
.B2(n_329),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_338),
.C(n_340),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_355),
.Y(n_357)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_356),
.A2(n_352),
.B(n_351),
.Y(n_358)
);

AOI322xp5_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_354),
.A3(n_348),
.B1(n_347),
.B2(n_353),
.C1(n_333),
.C2(n_349),
.Y(n_359)
);

FAx1_ASAP7_75t_SL g360 ( 
.A(n_359),
.B(n_355),
.CI(n_346),
.CON(n_360),
.SN(n_360)
);

AOI322xp5_ASAP7_75t_L g361 ( 
.A1(n_360),
.A2(n_335),
.A3(n_357),
.B1(n_338),
.B2(n_318),
.C1(n_306),
.C2(n_317),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_360),
.Y(n_362)
);


endmodule