module fake_jpeg_30434_n_266 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_266);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_266;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_149;
wire n_35;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_63),
.Y(n_70)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_59),
.Y(n_86)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_20),
.B(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_29),
.B(n_0),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_27),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_12),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_19),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_37),
.B1(n_27),
.B2(n_23),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_77),
.B1(n_49),
.B2(n_25),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_37),
.B1(n_38),
.B2(n_31),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_89),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_19),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_44),
.A2(n_50),
.B1(n_61),
.B2(n_55),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_53),
.B1(n_46),
.B2(n_48),
.Y(n_94)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_86),
.A3(n_71),
.B1(n_80),
.B2(n_28),
.Y(n_140)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_38),
.B1(n_23),
.B2(n_31),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_64),
.B1(n_59),
.B2(n_37),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_99),
.A2(n_109),
.B1(n_110),
.B2(n_119),
.Y(n_148)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_73),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_38),
.B1(n_31),
.B2(n_45),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_57),
.B1(n_60),
.B2(n_25),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_108),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_111),
.B(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_114),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_30),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_70),
.B(n_41),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_122),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_68),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

BUFx2_ASAP7_75t_SL g120 ( 
.A(n_86),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_121),
.B(n_80),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_26),
.C(n_36),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_41),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_89),
.B1(n_72),
.B2(n_90),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_86),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_132),
.A2(n_105),
.B1(n_97),
.B2(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_142),
.B1(n_100),
.B2(n_110),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_94),
.A2(n_69),
.B1(n_28),
.B2(n_30),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_135),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_42),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_115),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_80),
.B(n_96),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_154),
.B(n_165),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_158),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_151),
.A2(n_141),
.B(n_129),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_99),
.B1(n_121),
.B2(n_94),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_140),
.A2(n_111),
.B1(n_117),
.B2(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_164),
.B1(n_148),
.B2(n_128),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_129),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_93),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_69),
.B1(n_109),
.B2(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_42),
.B1(n_40),
.B2(n_35),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_32),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_147),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_40),
.B1(n_35),
.B2(n_2),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_32),
.B1(n_108),
.B2(n_98),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_108),
.B(n_98),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_147),
.B(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_169),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_161),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_153),
.B1(n_160),
.B2(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_179),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_135),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_175),
.C(n_139),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_130),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_134),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_180),
.Y(n_185)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_163),
.C(n_150),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_186),
.A2(n_188),
.B1(n_189),
.B2(n_175),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_174),
.B1(n_183),
.B2(n_181),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_154),
.B1(n_156),
.B2(n_162),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_181),
.A2(n_164),
.B1(n_165),
.B2(n_144),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_198),
.B1(n_178),
.B2(n_169),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_172),
.C(n_173),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_184),
.A2(n_177),
.B1(n_176),
.B2(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_188),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_191),
.B(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_212),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_193),
.C(n_185),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_189),
.B1(n_191),
.B2(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_209),
.A2(n_210),
.B1(n_197),
.B2(n_194),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_171),
.B1(n_144),
.B2(n_139),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_199),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_194),
.B(n_190),
.Y(n_214)
);

AOI221xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_137),
.B1(n_131),
.B2(n_130),
.C(n_144),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_196),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_220),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_218),
.B1(n_205),
.B2(n_211),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_208),
.C(n_185),
.Y(n_226)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_190),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_0),
.C(n_1),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_229),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_201),
.B(n_210),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_204),
.C(n_207),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_233),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_213),
.B(n_0),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_217),
.B1(n_225),
.B2(n_214),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_137),
.C(n_130),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_236),
.C(n_1),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

OAI22x1_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_218),
.B1(n_220),
.B2(n_216),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_238),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_224),
.B1(n_2),
.B2(n_4),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_241),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_12),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_236),
.C(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_250),
.Y(n_255)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_5),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_246),
.A2(n_238),
.B(n_244),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_240),
.C(n_239),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_5),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_247),
.A2(n_240),
.B1(n_6),
.B2(n_7),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_SL g257 ( 
.A1(n_254),
.A2(n_247),
.B(n_6),
.C(n_8),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_257),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_258),
.A2(n_253),
.B(n_255),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_256),
.C(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_SL g264 ( 
.A1(n_263),
.A2(n_261),
.B(n_9),
.C(n_11),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_9),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_265),
.A2(n_9),
.B(n_11),
.Y(n_266)
);


endmodule