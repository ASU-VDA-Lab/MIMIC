module fake_jpeg_1145_n_686 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_686);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_686;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_612;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_1),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_59),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_60),
.Y(n_163)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g164 ( 
.A(n_63),
.Y(n_164)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_66),
.B(n_72),
.Y(n_132)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_68),
.Y(n_199)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_70),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_73),
.B(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_30),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_80),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_76),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_81),
.B(n_89),
.Y(n_145)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_83),
.B(n_45),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_24),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g155 ( 
.A(n_86),
.Y(n_155)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_2),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_93),
.Y(n_204)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_94),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_98),
.Y(n_222)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_99),
.Y(n_208)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_57),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_102),
.B(n_114),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_51),
.B(n_2),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_36),
.B(n_2),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_33),
.B(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_117),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_26),
.Y(n_109)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_110),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_28),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_22),
.Y(n_112)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_40),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_115),
.Y(n_214)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_4),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_41),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_128),
.Y(n_180)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_39),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_42),
.Y(n_125)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_39),
.Y(n_126)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_42),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_47),
.Y(n_129)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_129),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_43),
.B(n_4),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_130),
.B(n_44),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_73),
.A2(n_48),
.B1(n_47),
.B2(n_56),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_139),
.A2(n_170),
.B1(n_191),
.B2(n_164),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_141),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_147),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_71),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_149),
.B(n_162),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_71),
.B(n_43),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_158),
.B(n_190),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_63),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_161),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_87),
.Y(n_162)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_166),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_120),
.A2(n_47),
.B1(n_48),
.B2(n_33),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_110),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_172),
.B(n_189),
.Y(n_264)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_75),
.Y(n_173)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_193),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_82),
.B(n_45),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_182),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_77),
.Y(n_184)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_68),
.Y(n_187)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_62),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_99),
.B(n_53),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_95),
.A2(n_48),
.B1(n_53),
.B2(n_44),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_92),
.Y(n_198)
);

CKINVDCx9p33_ASAP7_75t_R g256 ( 
.A(n_198),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_90),
.Y(n_200)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_200),
.Y(n_282)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_98),
.B(n_37),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_220),
.Y(n_238)
);

INVx6_ASAP7_75t_SL g210 ( 
.A(n_59),
.Y(n_210)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_97),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_212),
.B(n_213),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_111),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g216 ( 
.A1(n_70),
.A2(n_50),
.B(n_49),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_5),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_107),
.B(n_37),
.Y(n_220)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_115),
.Y(n_224)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

BUFx12_ASAP7_75t_L g225 ( 
.A(n_92),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_155),
.A2(n_113),
.B1(n_94),
.B2(n_107),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_227),
.A2(n_237),
.B1(n_251),
.B2(n_252),
.Y(n_325)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_141),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_228),
.Y(n_318)
);

CKINVDCx12_ASAP7_75t_R g231 ( 
.A(n_136),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_231),
.Y(n_322)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_232),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_146),
.B(n_49),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g368 ( 
.A(n_233),
.B(n_236),
.C(n_246),
.Y(n_368)
);

CKINVDCx12_ASAP7_75t_R g236 ( 
.A(n_136),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_204),
.A2(n_119),
.B1(n_109),
.B2(n_50),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_34),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_243),
.B(n_247),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_170),
.A2(n_211),
.B1(n_195),
.B2(n_34),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_244),
.A2(n_248),
.B1(n_284),
.B2(n_217),
.Y(n_315)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_245),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_163),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_133),
.B(n_119),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_145),
.B(n_5),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_250),
.B(n_272),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_204),
.A2(n_109),
.B1(n_127),
.B2(n_125),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_202),
.A2(n_129),
.B1(n_121),
.B2(n_93),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_152),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_253),
.Y(n_348)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_176),
.Y(n_254)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_160),
.A2(n_182),
.B(n_132),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_258),
.A2(n_268),
.B(n_279),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_186),
.A2(n_32),
.B1(n_31),
.B2(n_24),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_260),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_152),
.Y(n_261)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_197),
.A2(n_32),
.B1(n_31),
.B2(n_24),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_262),
.Y(n_351)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_159),
.Y(n_263)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_267),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_198),
.A2(n_24),
.B(n_32),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_269),
.A2(n_221),
.B(n_171),
.Y(n_331)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_201),
.Y(n_270)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_270),
.Y(n_334)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_165),
.Y(n_271)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_271),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_142),
.B(n_7),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_174),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_273),
.B(n_274),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_180),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_143),
.B(n_7),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_289),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_144),
.B(n_7),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_276),
.B(n_278),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_176),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_148),
.B(n_8),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_167),
.Y(n_280)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_280),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_150),
.B(n_8),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g362 ( 
.A1(n_281),
.A2(n_293),
.B(n_297),
.Y(n_362)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_201),
.Y(n_283)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_283),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_153),
.A2(n_31),
.B1(n_9),
.B2(n_10),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_181),
.Y(n_285)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_285),
.Y(n_341)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_183),
.Y(n_286)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_286),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_208),
.Y(n_287)
);

BUFx2_ASAP7_75t_SL g327 ( 
.A(n_287),
.Y(n_327)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_147),
.Y(n_288)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_288),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_156),
.B(n_8),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_178),
.Y(n_290)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_199),
.Y(n_292)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_292),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_138),
.B(n_10),
.Y(n_293)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_168),
.Y(n_295)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_295),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_135),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_269),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_151),
.B(n_11),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_217),
.Y(n_298)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_298),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_157),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_299),
.A2(n_196),
.B1(n_188),
.B2(n_214),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_199),
.B(n_12),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g365 ( 
.A1(n_301),
.A2(n_305),
.B(n_14),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_188),
.Y(n_302)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_302),
.Y(n_346)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_208),
.Y(n_303)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_303),
.Y(n_349)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_219),
.Y(n_304)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_304),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_154),
.B(n_12),
.Y(n_305)
);

OA22x2_ASAP7_75t_L g306 ( 
.A1(n_219),
.A2(n_14),
.B1(n_209),
.B2(n_207),
.Y(n_306)
);

AO22x1_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_209),
.B1(n_137),
.B2(n_223),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_235),
.B(n_222),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_308),
.B(n_309),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_242),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_238),
.B(n_137),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_310),
.B(n_330),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_315),
.A2(n_257),
.B1(n_265),
.B2(n_267),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_316),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_229),
.A2(n_135),
.B1(n_131),
.B2(n_184),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_319),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_264),
.B(n_185),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_323),
.B(n_335),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_248),
.A2(n_134),
.B1(n_205),
.B2(n_140),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_324),
.A2(n_326),
.B1(n_332),
.B2(n_333),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_256),
.A2(n_218),
.B1(n_214),
.B2(n_196),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_328),
.A2(n_234),
.B1(n_228),
.B2(n_291),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_266),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_331),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_299),
.A2(n_157),
.B1(n_192),
.B2(n_218),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_192),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_256),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_337),
.B(n_358),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_306),
.A2(n_200),
.B1(n_164),
.B2(n_131),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_344),
.A2(n_359),
.B1(n_319),
.B2(n_227),
.Y(n_406)
);

NAND2x1_ASAP7_75t_L g350 ( 
.A(n_226),
.B(n_169),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_350),
.A2(n_352),
.B(n_356),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_226),
.B(n_225),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_286),
.B(n_241),
.Y(n_353)
);

AND2x2_ASAP7_75t_SL g402 ( 
.A(n_353),
.B(n_282),
.Y(n_402)
);

NAND2xp33_ASAP7_75t_SL g356 ( 
.A(n_234),
.B(n_221),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_300),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_258),
.A2(n_134),
.B1(n_140),
.B2(n_205),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_306),
.B(n_169),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_361),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_255),
.B(n_169),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_300),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_365),
.Y(n_394)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_353),
.Y(n_372)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_364),
.Y(n_373)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_373),
.Y(n_443)
);

OAI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_376),
.A2(n_377),
.B1(n_342),
.B2(n_311),
.Y(n_429)
);

INVx13_ASAP7_75t_L g378 ( 
.A(n_322),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_378),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_379),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_354),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_380),
.B(n_396),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_316),
.A2(n_261),
.B1(n_302),
.B2(n_253),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_382),
.A2(n_401),
.B1(n_311),
.B2(n_342),
.Y(n_428)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_384),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_294),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_398),
.Y(n_438)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_386),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g387 ( 
.A1(n_316),
.A2(n_245),
.B(n_288),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_387),
.A2(n_361),
.B(n_350),
.Y(n_424)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_SL g450 ( 
.A1(n_388),
.A2(n_393),
.B1(n_395),
.B2(n_404),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_310),
.B(n_295),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_391),
.B(n_397),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_343),
.Y(n_393)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_338),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_323),
.B(n_259),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_346),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_357),
.B(n_240),
.Y(n_398)
);

OA22x2_ASAP7_75t_L g399 ( 
.A1(n_351),
.A2(n_252),
.B1(n_251),
.B2(n_262),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g451 ( 
.A1(n_399),
.A2(n_291),
.B(n_343),
.Y(n_451)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_403),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_360),
.A2(n_303),
.B1(n_230),
.B2(n_254),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_402),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_308),
.B(n_335),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_338),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_406),
.A2(n_351),
.B1(n_340),
.B2(n_325),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_333),
.A2(n_260),
.B1(n_296),
.B2(n_237),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_407),
.A2(n_340),
.B1(n_328),
.B2(n_332),
.Y(n_420)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_346),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_409),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_362),
.B(n_230),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_412),
.Y(n_427)
);

INVx6_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_414),
.Y(n_448)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_317),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_336),
.B(n_239),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_413),
.B(n_314),
.Y(n_431)
);

INVx5_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_318),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_415),
.B(n_416),
.Y(n_456)
);

INVx3_ASAP7_75t_SL g416 ( 
.A(n_329),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_419),
.A2(n_420),
.B1(n_422),
.B2(n_435),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_390),
.A2(n_328),
.B1(n_320),
.B2(n_314),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_371),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_423),
.B(n_434),
.C(n_449),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_424),
.A2(n_451),
.B(n_455),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_428),
.B(n_429),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_431),
.B(n_433),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_383),
.B(n_321),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_374),
.B(n_350),
.C(n_317),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_390),
.A2(n_345),
.B1(n_348),
.B2(n_318),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_375),
.Y(n_437)
);

INVx13_ASAP7_75t_L g465 ( 
.A(n_437),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_405),
.A2(n_271),
.B1(n_307),
.B2(n_341),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_440),
.A2(n_369),
.B1(n_376),
.B2(n_384),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_383),
.B(n_345),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_442),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_339),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_402),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_444),
.B(n_453),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_413),
.B(n_379),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_446),
.B(n_452),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_389),
.B(n_339),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_366),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_402),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_389),
.A2(n_307),
.B1(n_366),
.B2(n_313),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_454),
.A2(n_386),
.B1(n_388),
.B2(n_397),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_381),
.A2(n_294),
.B(n_367),
.Y(n_455)
);

MAJx2_ASAP7_75t_L g457 ( 
.A(n_392),
.B(n_368),
.C(n_313),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_457),
.B(n_400),
.C(n_240),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_409),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_458),
.B(n_472),
.Y(n_507)
);

BUFx12f_ASAP7_75t_L g460 ( 
.A(n_436),
.Y(n_460)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_460),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_452),
.A2(n_387),
.B(n_392),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_462),
.B(n_488),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_427),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_463),
.A2(n_467),
.B1(n_480),
.B2(n_481),
.Y(n_515)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_427),
.Y(n_466)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_466),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_436),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_468),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_470),
.A2(n_471),
.B1(n_473),
.B2(n_475),
.Y(n_521)
);

OAI21xp33_ASAP7_75t_L g471 ( 
.A1(n_431),
.A2(n_394),
.B(n_387),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_418),
.B(n_334),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_440),
.A2(n_381),
.B1(n_407),
.B2(n_399),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_443),
.Y(n_474)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_474),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_451),
.A2(n_382),
.B1(n_401),
.B2(n_370),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_423),
.B(n_385),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_477),
.B(n_434),
.C(n_457),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_433),
.B(n_373),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_478),
.B(n_483),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_436),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_447),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_422),
.B(n_334),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_489),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_439),
.A2(n_399),
.B(n_372),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_486),
.A2(n_439),
.B(n_455),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_441),
.B(n_412),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_487),
.B(n_454),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_444),
.B(n_399),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_447),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_417),
.B(n_410),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_491),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_438),
.B(n_378),
.Y(n_491)
);

CKINVDCx14_ASAP7_75t_R g492 ( 
.A(n_424),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_492),
.Y(n_503)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_445),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_493),
.B(n_417),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_494),
.A2(n_428),
.B1(n_430),
.B2(n_453),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_435),
.Y(n_516)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_496),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_490),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_497),
.B(n_498),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_485),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_461),
.B(n_393),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_500),
.B(n_504),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_501),
.A2(n_518),
.B(n_511),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_502),
.A2(n_530),
.B1(n_479),
.B2(n_475),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_425),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_505),
.B(n_516),
.Y(n_550)
);

XNOR2x2_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_425),
.Y(n_508)
);

OAI21xp33_ASAP7_75t_L g561 ( 
.A1(n_508),
.A2(n_480),
.B(n_397),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_449),
.C(n_442),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_512),
.B(n_522),
.C(n_462),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_464),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_513),
.B(n_528),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_476),
.B(n_477),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_517),
.B(n_519),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_459),
.A2(n_446),
.B(n_451),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_421),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_460),
.Y(n_520)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_520),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_466),
.B(n_421),
.C(n_430),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_470),
.A2(n_420),
.B1(n_451),
.B2(n_426),
.Y(n_523)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_523),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_487),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_524),
.B(n_525),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_464),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_469),
.B(n_426),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_526),
.B(n_465),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_481),
.B(n_367),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_529),
.B(n_531),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_482),
.A2(n_432),
.B1(n_448),
.B2(n_456),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_469),
.B(n_463),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_499),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_534),
.B(n_554),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_535),
.A2(n_542),
.B1(n_530),
.B2(n_511),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_521),
.A2(n_482),
.B1(n_488),
.B2(n_479),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_536),
.A2(n_460),
.B1(n_411),
.B2(n_298),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_537),
.B(n_526),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_525),
.A2(n_479),
.B1(n_488),
.B2(n_489),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_538),
.A2(n_551),
.B1(n_502),
.B2(n_515),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_432),
.C(n_486),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_539),
.B(n_541),
.C(n_519),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_493),
.C(n_484),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_518),
.A2(n_459),
.B1(n_491),
.B2(n_465),
.Y(n_542)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_499),
.Y(n_547)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_547),
.Y(n_575)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_522),
.Y(n_549)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_549),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_506),
.A2(n_494),
.B1(n_474),
.B2(n_468),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_503),
.B(n_414),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_552),
.B(n_555),
.Y(n_580)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_527),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_503),
.B(n_312),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_520),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_556),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_507),
.B(n_312),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_557),
.B(n_558),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_501),
.A2(n_465),
.B(n_467),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_559),
.B(n_560),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_509),
.B(n_347),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_561),
.B(n_562),
.Y(n_592)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_527),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_524),
.B(n_347),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_563),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_564),
.B(n_511),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_566),
.A2(n_571),
.B1(n_538),
.B2(n_545),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_567),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_569),
.B(n_570),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_505),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_545),
.A2(n_514),
.B1(n_506),
.B2(n_516),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_572),
.B(n_544),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_553),
.B(n_508),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_573),
.B(n_578),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g579 ( 
.A(n_548),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_579),
.B(n_582),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_SL g581 ( 
.A(n_550),
.B(n_514),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_SL g593 ( 
.A(n_581),
.B(n_535),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_537),
.B(n_532),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_550),
.B(n_532),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_583),
.B(n_586),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_548),
.A2(n_510),
.B1(n_450),
.B2(n_460),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_584),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_541),
.B(n_395),
.C(n_404),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_585),
.B(n_588),
.C(n_589),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_549),
.B(n_416),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_539),
.B(n_408),
.C(n_239),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_558),
.B(n_510),
.C(n_283),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_591),
.A2(n_559),
.B1(n_547),
.B2(n_542),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_SL g618 ( 
.A(n_593),
.B(n_569),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_582),
.B(n_546),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_594),
.B(n_282),
.Y(n_629)
);

NAND2x1p5_ASAP7_75t_R g597 ( 
.A(n_566),
.B(n_564),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_597),
.B(n_611),
.Y(n_633)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_599),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_572),
.B(n_583),
.C(n_585),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_600),
.B(n_612),
.C(n_589),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_603),
.B(n_613),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_573),
.B(n_536),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_604),
.B(n_574),
.Y(n_622)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_568),
.Y(n_605)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_605),
.Y(n_627)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_587),
.Y(n_606)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_606),
.Y(n_628)
);

XNOR2x1_ASAP7_75t_L g634 ( 
.A(n_607),
.B(n_608),
.Y(n_634)
);

OA22x2_ASAP7_75t_L g608 ( 
.A1(n_571),
.A2(n_551),
.B1(n_565),
.B2(n_556),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_575),
.Y(n_609)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_609),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_592),
.A2(n_540),
.B(n_543),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_590),
.B(n_533),
.C(n_562),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_580),
.Y(n_613)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_577),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_615),
.B(n_577),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_611),
.A2(n_588),
.B(n_586),
.Y(n_616)
);

OAI21x1_ASAP7_75t_SL g639 ( 
.A1(n_616),
.A2(n_601),
.B(n_596),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_602),
.A2(n_581),
.B1(n_533),
.B2(n_576),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_617),
.A2(n_604),
.B1(n_608),
.B2(n_595),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_618),
.B(n_623),
.Y(n_649)
);

OAI22x1_ASAP7_75t_L g619 ( 
.A1(n_602),
.A2(n_599),
.B1(n_597),
.B2(n_608),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_619),
.B(n_622),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_621),
.B(n_625),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_595),
.B(n_570),
.Y(n_623)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_624),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_600),
.B(n_565),
.C(n_554),
.Y(n_625)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_629),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_603),
.B(n_249),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_631),
.B(n_632),
.Y(n_647)
);

FAx1_ASAP7_75t_L g632 ( 
.A(n_593),
.B(n_327),
.CI(n_166),
.CON(n_632),
.SN(n_632)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_632),
.A2(n_612),
.B(n_610),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g651 ( 
.A(n_637),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g659 ( 
.A1(n_639),
.A2(n_645),
.B(n_626),
.Y(n_659)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_625),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_640),
.B(n_641),
.Y(n_653)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_630),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_620),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_642),
.B(n_643),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_621),
.B(n_614),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_633),
.A2(n_614),
.B(n_607),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_617),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_646),
.B(n_647),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_648),
.B(n_650),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_627),
.B(n_608),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_644),
.B(n_623),
.Y(n_652)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_652),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_636),
.B(n_628),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_654),
.B(n_659),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_649),
.B(n_633),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_655),
.A2(n_658),
.B(n_637),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_645),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_657),
.B(n_661),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_649),
.B(n_622),
.Y(n_658)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_648),
.B(n_598),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_663),
.A2(n_666),
.B(n_670),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_656),
.B(n_638),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_664),
.B(n_665),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_653),
.B(n_635),
.C(n_634),
.Y(n_665)
);

INVxp33_ASAP7_75t_L g666 ( 
.A(n_662),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_SL g669 ( 
.A1(n_660),
.A2(n_635),
.B(n_654),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_669),
.A2(n_270),
.B(n_249),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g670 ( 
.A(n_651),
.B(n_634),
.C(n_619),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_667),
.B(n_651),
.C(n_618),
.Y(n_672)
);

XNOR2xp5_ASAP7_75t_L g679 ( 
.A(n_672),
.B(n_674),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_SL g673 ( 
.A1(n_668),
.A2(n_632),
.B(n_598),
.Y(n_673)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_673),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_666),
.B(n_277),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_676),
.B(n_671),
.C(n_232),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g682 ( 
.A(n_680),
.B(n_675),
.C(n_671),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_679),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_681),
.B(n_682),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g684 ( 
.A(n_683),
.B(n_678),
.C(n_677),
.Y(n_684)
);

XOR2xp5_ASAP7_75t_L g685 ( 
.A(n_684),
.B(n_277),
.Y(n_685)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_685),
.B(n_277),
.C(n_215),
.Y(n_686)
);


endmodule