module fake_jpeg_9375_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_22),
.Y(n_52)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_39),
.B1(n_32),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_32),
.B1(n_22),
.B2(n_27),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_32),
.B1(n_18),
.B2(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_27),
.B1(n_29),
.B2(n_33),
.Y(n_85)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_21),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_33),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_63),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_62),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_71),
.Y(n_97)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_26),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_34),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_19),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_83),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_91),
.B1(n_92),
.B2(n_109),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_55),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_78),
.B(n_24),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_32),
.B(n_29),
.C(n_35),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_85),
.A2(n_95),
.B1(n_54),
.B2(n_16),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_27),
.B1(n_26),
.B2(n_28),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_29),
.C(n_35),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_94),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_88),
.B(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_27),
.B1(n_35),
.B2(n_31),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_34),
.B1(n_31),
.B2(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_93),
.B(n_96),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_28),
.B1(n_31),
.B2(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_30),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_28),
.B1(n_30),
.B2(n_16),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_69),
.B1(n_61),
.B2(n_54),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_24),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_62),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_30),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_66),
.CI(n_60),
.CON(n_117),
.SN(n_117)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVxp67_ASAP7_75t_SL g127 ( 
.A(n_104),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_1),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_106),
.B(n_20),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_1),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_49),
.A2(n_34),
.B1(n_23),
.B2(n_20),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_49),
.A2(n_23),
.B1(n_20),
.B2(n_30),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_23),
.B1(n_51),
.B2(n_61),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_114),
.B(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_118),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_126),
.B1(n_91),
.B2(n_81),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_78),
.A2(n_51),
.A3(n_62),
.B1(n_60),
.B2(n_47),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_123),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_78),
.B(n_75),
.C(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_135),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_134),
.A2(n_93),
.B1(n_80),
.B2(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_62),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_96),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_140),
.A2(n_76),
.B1(n_81),
.B2(n_90),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_144),
.B(n_145),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_74),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_149),
.B(n_151),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_150),
.A2(n_113),
.B(n_112),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_162),
.B1(n_167),
.B2(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_124),
.B1(n_132),
.B2(n_112),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_94),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_164),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_115),
.A2(n_100),
.B1(n_106),
.B2(n_105),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_94),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_168),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_115),
.A2(n_106),
.B1(n_105),
.B2(n_87),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_103),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_102),
.C(n_110),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_130),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_90),
.B1(n_76),
.B2(n_92),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_77),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_175),
.Y(n_204)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_77),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_136),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_176),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_124),
.B1(n_131),
.B2(n_129),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_177),
.A2(n_150),
.B1(n_65),
.B2(n_24),
.Y(n_233)
);

XNOR2x2_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_120),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_178),
.A2(n_180),
.B(n_189),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_136),
.B(n_141),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_207),
.C(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_187),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

AOI21x1_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_141),
.B(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_197),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_113),
.C(n_136),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_192),
.B(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_202),
.B(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_117),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_149),
.A2(n_127),
.B(n_104),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_143),
.B(n_102),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_203),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_154),
.B(n_110),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_24),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_72),
.B1(n_56),
.B2(n_57),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_158),
.B1(n_173),
.B2(n_174),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_189),
.A2(n_155),
.B1(n_144),
.B2(n_170),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_210),
.A2(n_226),
.B(n_202),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_212),
.B(n_214),
.C(n_218),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_159),
.C(n_164),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_215),
.B(n_224),
.Y(n_253)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_228),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_167),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_153),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_148),
.Y(n_223)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_151),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_162),
.C(n_163),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_230),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_221),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_249),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_198),
.B1(n_201),
.B2(n_193),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_242),
.B1(n_257),
.B2(n_227),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_234),
.B1(n_225),
.B2(n_219),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_213),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_196),
.B(n_197),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_244),
.Y(n_263)
);

INVxp33_ASAP7_75t_SL g246 ( 
.A(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

OAI32xp33_ASAP7_75t_L g248 ( 
.A1(n_236),
.A2(n_199),
.A3(n_191),
.B1(n_183),
.B2(n_186),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_213),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_187),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_182),
.B(n_186),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_259),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_206),
.B1(n_190),
.B2(n_184),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_261),
.A2(n_269),
.B(n_255),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_259),
.A2(n_228),
.B1(n_217),
.B2(n_210),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_264),
.A2(n_274),
.B1(n_279),
.B2(n_239),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_265),
.B(n_244),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_212),
.C(n_214),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_267),
.C(n_272),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_223),
.C(n_218),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_270),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_241),
.A2(n_217),
.B1(n_232),
.B2(n_211),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_183),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_207),
.C(n_232),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_65),
.B1(n_72),
.B2(n_57),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_99),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_277),
.C(n_278),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_242),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_99),
.C(n_108),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_122),
.B1(n_108),
.B2(n_56),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_287),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_252),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_296),
.C(n_272),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_277),
.B(n_258),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_289),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_245),
.B(n_240),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_245),
.B(n_251),
.Y(n_288)
);

OAI321xp33_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_279),
.A3(n_278),
.B1(n_10),
.B2(n_11),
.C(n_14),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_239),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_257),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_295),
.B1(n_273),
.B2(n_265),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_255),
.C(n_248),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_12),
.C(n_11),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_247),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_303),
.B(n_304),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_267),
.C(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_306),
.Y(n_310)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_268),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_307),
.C(n_282),
.Y(n_312)
);

OAI221xp5_ASAP7_75t_L g304 ( 
.A1(n_287),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.C(n_12),
.Y(n_304)
);

OA21x2_ASAP7_75t_L g305 ( 
.A1(n_283),
.A2(n_2),
.B(n_3),
.Y(n_305)
);

O2A1O1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_13),
.C(n_12),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_294),
.B1(n_284),
.B2(n_296),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_312),
.C(n_315),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_291),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_314),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_291),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_10),
.B(n_9),
.Y(n_315)
);

AOI221xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_298),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_319),
.A2(n_9),
.B(n_4),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_317),
.A2(n_298),
.B1(n_305),
.B2(n_302),
.Y(n_320)
);

AOI31xp67_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_325),
.A3(n_326),
.B(n_316),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_305),
.C(n_310),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_324),
.Y(n_329)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_3),
.C(n_4),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_327),
.A2(n_326),
.B(n_7),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_319),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_330),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_24),
.Y(n_330)
);

NAND3xp33_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_329),
.C(n_7),
.Y(n_333)
);

NOR3xp33_ASAP7_75t_SL g334 ( 
.A(n_333),
.B(n_5),
.C(n_8),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_5),
.C(n_8),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_332),
.Y(n_336)
);


endmodule