module real_jpeg_13184_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_3),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_3),
.B(n_34),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_3),
.B(n_29),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_3),
.B(n_86),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_4),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_4),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_4),
.B(n_69),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_4),
.B(n_27),
.Y(n_155)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_7),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_7),
.B(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_8),
.B(n_34),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_8),
.B(n_69),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_8),
.B(n_54),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_11),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_11),
.B(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_11),
.B(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_11),
.B(n_54),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_11),
.B(n_29),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_11),
.B(n_86),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_11),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_13),
.B(n_29),
.Y(n_107)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_14),
.B(n_38),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_14),
.B(n_86),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_14),
.B(n_27),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_15),
.B(n_29),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_15),
.B(n_54),
.Y(n_126)
);

HAxp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_138),
.CON(n_16),
.SN(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_100),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_20),
.B(n_100),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_64),
.C(n_87),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_21),
.A2(n_22),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_22),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_39),
.CI(n_47),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_23),
.B(n_39),
.C(n_47),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.C(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_24),
.A2(n_25),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_26),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_26),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_26),
.A2(n_28),
.B1(n_108),
.B2(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_28),
.Y(n_168)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_30),
.B(n_42),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_30),
.B(n_63),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_32),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B(n_46),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_42),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_44),
.B(n_84),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_44),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_46),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_58),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_SL g86 ( 
.A(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_51),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_51),
.B(n_63),
.Y(n_185)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_53),
.B(n_56),
.C(n_58),
.Y(n_134)
);

INVx5_ASAP7_75t_SL g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_64),
.A2(n_65),
.B1(n_87),
.B2(n_88),
.Y(n_219)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_73),
.B2(n_74),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_66),
.B(n_75),
.C(n_79),
.Y(n_135)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_67),
.Y(n_224)
);

FAx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.CI(n_72),
.CON(n_67),
.SN(n_67)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_71),
.C(n_72),
.Y(n_111)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_93),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.C(n_85),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_91),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.C(n_94),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_89),
.B(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_92),
.B(n_94),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_97),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_116),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_114),
.B2(n_115),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_110),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_107),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_111),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_135),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_127),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_125),
.B2(n_126),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_121),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_122),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_215),
.B(n_220),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_200),
.B(n_214),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_170),
.B(n_199),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_156),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_142),
.B(n_156),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.C(n_151),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_196),
.Y(n_195)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_145),
.CI(n_146),
.CON(n_143),
.SN(n_143)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_152),
.B(n_155),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_163),
.B2(n_169),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_162),
.C(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_193),
.B(n_198),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_183),
.B(n_192),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_178),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_181),
.C(n_182),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_187),
.B(n_191),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_185),
.B(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_201),
.B(n_202),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_208),
.C(n_213),
.Y(n_216)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);


endmodule