module fake_jpeg_9417_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_40),
.Y(n_49)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_28),
.B1(n_17),
.B2(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_50),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_51),
.B1(n_56),
.B2(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_63),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_28),
.B1(n_17),
.B2(n_27),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_24),
.B1(n_18),
.B2(n_26),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_42),
.B1(n_37),
.B2(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_1),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_68),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_36),
.B(n_26),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_60),
.B1(n_50),
.B2(n_52),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_85),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_81),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_42),
.B1(n_35),
.B2(n_40),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_83),
.B1(n_90),
.B2(n_34),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_33),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_82),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_43),
.B1(n_39),
.B2(n_35),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_53),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_34),
.B1(n_39),
.B2(n_22),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_106),
.B1(n_108),
.B2(n_85),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_100),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_98),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_71),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_86),
.B(n_80),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_105),
.C(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_77),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_30),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_70),
.B(n_81),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_66),
.B(n_47),
.C(n_33),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_112),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_74),
.A2(n_53),
.B1(n_46),
.B2(n_47),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_65),
.C(n_55),
.Y(n_110)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_124),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_106),
.B(n_108),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_127),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_70),
.B1(n_69),
.B2(n_66),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_135),
.B1(n_107),
.B2(n_96),
.Y(n_137)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_95),
.C(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_134),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_69),
.C(n_66),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_93),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_109),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_97),
.B(n_92),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_143),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_137),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_99),
.B(n_105),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_142),
.B(n_147),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_97),
.B(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_94),
.Y(n_144)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_96),
.B1(n_101),
.B2(n_106),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_135),
.B1(n_96),
.B2(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_150),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_129),
.B1(n_118),
.B2(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_154),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_153),
.B(n_155),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_119),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_112),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_144),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_132),
.B1(n_130),
.B2(n_128),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_139),
.B(n_143),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_116),
.C(n_126),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_154),
.B(n_153),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_161),
.A2(n_167),
.B(n_148),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_166),
.B1(n_30),
.B2(n_3),
.Y(n_187)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_168),
.Y(n_177)
);

OAI22x1_ASAP7_75t_SL g166 ( 
.A1(n_147),
.A2(n_134),
.B1(n_121),
.B2(n_21),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_137),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_121),
.B1(n_113),
.B2(n_25),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_150),
.B1(n_25),
.B2(n_30),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_25),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_151),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_179),
.B(n_182),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_152),
.B1(n_148),
.B2(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_171),
.A2(n_142),
.B(n_140),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_183),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_184),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_188),
.Y(n_191)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_186),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_13),
.B1(n_25),
.B2(n_30),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_187),
.B(n_6),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_2),
.B(n_3),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_195),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_157),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_178),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_157),
.C(n_158),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_175),
.C(n_177),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_183),
.B1(n_162),
.B2(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_206),
.C(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_167),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_208),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_6),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_194),
.A2(n_176),
.B1(n_160),
.B2(n_185),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_190),
.B1(n_199),
.B2(n_172),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_168),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_188),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_204),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_198),
.A2(n_186),
.B(n_189),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_190),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_214),
.B(n_216),
.Y(n_221)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_215),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_196),
.B(n_8),
.Y(n_214)
);

AOI21x1_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_205),
.B(n_215),
.Y(n_217)
);

O2A1O1Ixp5_ASAP7_75t_SL g224 ( 
.A1(n_217),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_211),
.A2(n_201),
.B(n_206),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_210),
.C(n_9),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_6),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_11),
.B(n_12),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_220),
.B1(n_221),
.B2(n_225),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_12),
.Y(n_229)
);


endmodule