module real_jpeg_23415_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_354, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_354;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_2),
.A2(n_61),
.B1(n_65),
.B2(n_68),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_61),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_2),
.A2(n_61),
.B1(n_80),
.B2(n_83),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g87 ( 
.A(n_4),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_5),
.A2(n_65),
.B1(n_68),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_5),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_76),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_76),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_5),
.A2(n_76),
.B1(n_80),
.B2(n_83),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_6),
.A2(n_51),
.B1(n_65),
.B2(n_68),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_6),
.A2(n_51),
.B1(n_80),
.B2(n_83),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_7),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_7),
.A2(n_67),
.B1(n_80),
.B2(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_67),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_8),
.B(n_91),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_8),
.B(n_30),
.C(n_46),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_81),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_8),
.B(n_74),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_27),
.B1(n_170),
.B2(n_173),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_10),
.A2(n_83),
.B1(n_90),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_10),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_10),
.A2(n_65),
.B1(n_68),
.B2(n_94),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_94),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_94),
.Y(n_170)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_12),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_12),
.A2(n_35),
.B1(n_65),
.B2(n_68),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_12),
.A2(n_35),
.B1(n_322),
.B2(n_324),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_14),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_14),
.A2(n_38),
.B1(n_65),
.B2(n_68),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_14),
.A2(n_38),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_346),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_333),
.B(n_345),
.Y(n_17)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_296),
.A3(n_326),
.B1(n_331),
.B2(n_332),
.C(n_354),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_268),
.B(n_295),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_239),
.B(n_267),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_132),
.B(n_218),
.C(n_238),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_116),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_23),
.B(n_116),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_95),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_58),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_25),
.B(n_58),
.C(n_95),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_26),
.B(n_43),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_36),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_27),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_27),
.A2(n_40),
.B1(n_163),
.B2(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_27),
.A2(n_36),
.B(n_152),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_27),
.A2(n_152),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_28),
.A2(n_34),
.B1(n_39),
.B2(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_28),
.B(n_37),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_28),
.A2(n_150),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_29),
.B(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_31),
.Y(n_173)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_32),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_32),
.B(n_81),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_42),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B(n_52),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_57),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_44),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_44),
.A2(n_54),
.B1(n_145),
.B2(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_44),
.B(n_81),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_44),
.A2(n_54),
.B(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_45),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_47),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_49),
.B1(n_71),
.B2(n_72),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_48),
.A2(n_72),
.B(n_184),
.C(n_186),
.Y(n_183)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_49),
.B(n_140),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g186 ( 
.A(n_49),
.B(n_68),
.C(n_71),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_52),
.B(n_208),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_60),
.B(n_62),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_53),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_53),
.A2(n_143),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_53),
.A2(n_143),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_54),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_54),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_77),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_59),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_60),
.B(n_143),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_60),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_62),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_63)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_68),
.B1(n_86),
.B2(n_88),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_65),
.A2(n_82),
.B(n_86),
.C(n_114),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g185 ( 
.A(n_65),
.B(n_81),
.CON(n_185),
.SN(n_185)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_83),
.C(n_88),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_69),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_69),
.A2(n_74),
.B1(n_130),
.B2(n_185),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_69),
.A2(n_107),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_69),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_69),
.A2(n_74),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_69),
.A2(n_235),
.B(n_275),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_69),
.A2(n_74),
.B(n_107),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_73),
.A2(n_105),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_73),
.B(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_73),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_74),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_91),
.B2(n_92),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B(n_82),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_79),
.Y(n_288)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_80),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_84),
.A2(n_91),
.B1(n_101),
.B2(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_84),
.B(n_286),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_84),
.A2(n_91),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_84),
.A2(n_321),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_85),
.A2(n_301),
.B(n_302),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_91),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_91),
.B(n_286),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_108),
.B2(n_115),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_98),
.B(n_103),
.C(n_115),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_99),
.A2(n_255),
.B(n_256),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_99),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g323 ( 
.A(n_102),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B(n_106),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_106),
.B(n_261),
.Y(n_318)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_123),
.B(n_125),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.C(n_121),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_117),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_119),
.B(n_121),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_128),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_125),
.B(n_149),
.Y(n_224)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_128),
.B(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_217),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_212),
.B(n_216),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_196),
.B(n_211),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_179),
.B(n_195),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_159),
.B(n_178),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_146),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_146),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_141),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_147),
.B(n_154),
.C(n_157),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_166),
.B(n_177),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_165),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_171),
.B(n_176),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_194),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_194),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_190),
.C(n_191),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_187),
.B2(n_188),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_193),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_198),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_206),
.C(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_215),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_220),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_237),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_229),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_229),
.C(n_237),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_228),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_228),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_227),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_232),
.C(n_234),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_240),
.B(n_241),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_266),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_251),
.B1(n_264),
.B2(n_265),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_265),
.C(n_266),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_250),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_244),
.A2(n_245),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_244),
.A2(n_279),
.B(n_283),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_258),
.C(n_263),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_258),
.B1(n_259),
.B2(n_263),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_256),
.B(n_302),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_257),
.Y(n_284)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_260),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_269),
.B(n_270),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_270)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_278),
.B1(n_290),
.B2(n_291),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_276),
.B(n_277),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_276),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_277),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_277),
.A2(n_298),
.B1(n_310),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_290),
.C(n_294),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_289),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_285),
.Y(n_340)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_292),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_312),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_312),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_310),
.C(n_311),
.Y(n_297)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_303),
.B2(n_304),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_300),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_305),
.C(n_309),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_315),
.C(n_325),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_301),
.Y(n_320)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_306),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_317),
.C(n_319),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_325),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_335),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_343),
.B2(n_344),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_341),
.B2(n_342),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_338),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_339),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_341),
.C(n_343),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_351),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_348),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_352),
.Y(n_351)
);


endmodule