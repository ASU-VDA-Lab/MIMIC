module fake_jpeg_8258_n_334 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_16),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_34),
.B1(n_29),
.B2(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_63),
.B1(n_36),
.B2(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_36),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_18),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_25),
.B1(n_19),
.B2(n_23),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_20),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_20),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_39),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_73),
.B(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_84),
.Y(n_112)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_81),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_31),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_26),
.B(n_17),
.C(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_89),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_39),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_25),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_56),
.B1(n_46),
.B2(n_38),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_108),
.B(n_110),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_50),
.B1(n_59),
.B2(n_66),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_115),
.B1(n_121),
.B2(n_86),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_71),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_25),
.B(n_41),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_50),
.B1(n_47),
.B2(n_66),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_48),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_118),
.B(n_123),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_124),
.B1(n_94),
.B2(n_26),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_18),
.B1(n_46),
.B2(n_38),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_86),
.B1(n_24),
.B2(n_30),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_72),
.A2(n_48),
.B1(n_38),
.B2(n_46),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_62),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_127),
.A2(n_132),
.B1(n_137),
.B2(n_142),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_134),
.B(n_141),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_76),
.CI(n_82),
.CON(n_130),
.SN(n_130)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_118),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_82),
.C(n_77),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_124),
.C(n_104),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_40),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_62),
.B1(n_92),
.B2(n_81),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_139),
.B1(n_145),
.B2(n_147),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_SL g138 ( 
.A(n_114),
.B(n_77),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_114),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_79),
.B1(n_89),
.B2(n_63),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_143),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_41),
.B1(n_80),
.B2(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_17),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_113),
.B(n_28),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_24),
.B(n_41),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_113),
.B(n_112),
.Y(n_159)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_160),
.Y(n_197)
);

HAxp5_ASAP7_75t_SL g208 ( 
.A(n_159),
.B(n_164),
.CON(n_208),
.SN(n_208)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_168),
.B(n_171),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_169),
.A2(n_28),
.B(n_21),
.Y(n_211)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_172),
.B(n_175),
.Y(n_201)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_114),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_106),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_102),
.C(n_103),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_179),
.B(n_180),
.Y(n_205)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_102),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_182),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_98),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_98),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_154),
.B1(n_148),
.B2(n_136),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_185),
.A2(n_187),
.B1(n_190),
.B2(n_193),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_142),
.B1(n_131),
.B2(n_137),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_174),
.A2(n_139),
.B1(n_127),
.B2(n_147),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_188),
.A2(n_200),
.B1(n_203),
.B2(n_198),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_132),
.B1(n_141),
.B2(n_149),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_192),
.Y(n_222)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_129),
.B1(n_133),
.B2(n_151),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_134),
.B1(n_146),
.B2(n_130),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_199),
.B1(n_204),
.B2(n_99),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_170),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_202),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_150),
.B1(n_126),
.B2(n_128),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_173),
.A2(n_128),
.B1(n_150),
.B2(n_116),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_158),
.A2(n_116),
.B1(n_111),
.B2(n_122),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_158),
.A2(n_107),
.B1(n_99),
.B2(n_117),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_207),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_11),
.B(n_16),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_176),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_220),
.C(n_224),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_196),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_215),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_183),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_161),
.B1(n_160),
.B2(n_159),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_216),
.A2(n_219),
.B1(n_227),
.B2(n_231),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_218),
.B(n_211),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_162),
.B1(n_157),
.B2(n_169),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_178),
.C(n_122),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_230),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_107),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_208),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_96),
.C(n_80),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_229),
.C(n_234),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_96),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_205),
.B1(n_184),
.B2(n_192),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_235),
.B1(n_221),
.B2(n_228),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_96),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_184),
.A2(n_33),
.B1(n_23),
.B2(n_27),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_0),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_27),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_33),
.C(n_23),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_242),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_209),
.B1(n_206),
.B2(n_201),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_244),
.B1(n_257),
.B2(n_220),
.Y(n_268)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_247),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_191),
.B1(n_208),
.B2(n_187),
.Y(n_244)
);

INVx13_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_226),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_10),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_251),
.B(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_253),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_212),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_SL g255 ( 
.A1(n_237),
.A2(n_33),
.B(n_23),
.C(n_3),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_255),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_27),
.C(n_33),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_260),
.C(n_229),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_9),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_258),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_1),
.C(n_2),
.Y(n_260)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_224),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_270),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_265),
.A2(n_254),
.B1(n_255),
.B2(n_260),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_249),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_1),
.C(n_2),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_273),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_4),
.C(n_5),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_11),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_275),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g279 ( 
.A(n_276),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_240),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_282),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_286),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_245),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_245),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_255),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_291),
.C(n_293),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_256),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_12),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_289),
.A2(n_267),
.B1(n_278),
.B2(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_295),
.B(n_302),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_289),
.A2(n_278),
.B1(n_276),
.B2(n_263),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_6),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_270),
.C(n_269),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_298),
.B(n_6),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_274),
.C(n_273),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_277),
.C(n_265),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_8),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_284),
.A2(n_255),
.B1(n_5),
.B2(n_7),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_5),
.B1(n_13),
.B2(n_14),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_12),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_283),
.Y(n_307)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_280),
.B1(n_285),
.B2(n_8),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_314),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_313),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_315),
.B(n_15),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_8),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_10),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_316),
.A2(n_305),
.B1(n_304),
.B2(n_301),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_299),
.C(n_297),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_320),
.Y(n_326)
);

OA21x2_ASAP7_75t_SL g321 ( 
.A1(n_307),
.A2(n_306),
.B(n_15),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_321),
.B(n_15),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_316),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_325),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_311),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_328),
.C(n_319),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_323),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_324),
.B(n_326),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_329),
.C(n_318),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_5),
.Y(n_334)
);


endmodule