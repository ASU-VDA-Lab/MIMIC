module fake_netlist_6_867_n_1561 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1561);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1561;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1558;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_1159;
wire n_995;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_1045;
wire n_706;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_329),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_318),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_162),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_245),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_128),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_175),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_18),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_334),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_144),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_324),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_159),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_332),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_326),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_51),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_130),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_312),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_196),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_140),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_233),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_96),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_290),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_145),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_202),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_8),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_293),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_157),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_246),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_44),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_230),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_248),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_208),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_127),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_73),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_261),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_272),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_243),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_139),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_235),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_176),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_20),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_224),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_274),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_21),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_276),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_153),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_288),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_189),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_80),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_22),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_44),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_242),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_118),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_240),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_19),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_103),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_109),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_3),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_41),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_260),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_119),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_165),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_24),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_94),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_126),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_11),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_309),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_84),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_46),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_84),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_308),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_61),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_194),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_207),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_41),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_249),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_89),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_78),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_95),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_234),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_164),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_184),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_170),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_232),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_10),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_20),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_297),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_268),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_163),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_200),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_201),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_124),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_215),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_85),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_147),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_273),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_244),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_228),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_173),
.Y(n_435)
);

BUFx10_ASAP7_75t_L g436 ( 
.A(n_198),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_148),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_18),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_38),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_313),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_295),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_285),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_40),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_229),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_307),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_160),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_73),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_89),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_289),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_169),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_65),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_16),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_158),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_120),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_32),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_315),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_52),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_180),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_331),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_193),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_83),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_281),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_92),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_252),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_287),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_117),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_271),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_104),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_24),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_333),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_12),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_27),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_116),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_320),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_66),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_236),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_129),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_282),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_108),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_174),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_36),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_300),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_150),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_106),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_79),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_76),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_143),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_283),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_97),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_294),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_166),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_155),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_278),
.Y(n_493)
);

BUFx5_ASAP7_75t_L g494 ( 
.A(n_185),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_74),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_29),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_77),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_183),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_99),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_133),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_15),
.Y(n_501)
);

BUFx10_ASAP7_75t_L g502 ( 
.A(n_112),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_152),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_269),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_78),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_34),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_188),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_266),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_137),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_86),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_227),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_23),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_146),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_75),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_330),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_6),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_179),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g518 ( 
.A(n_284),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_26),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_4),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_132),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_32),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_31),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_327),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_265),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_98),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_34),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_204),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_85),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_182),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_45),
.Y(n_531)
);

CKINVDCx14_ASAP7_75t_R g532 ( 
.A(n_53),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_5),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_161),
.Y(n_534)
);

BUFx8_ASAP7_75t_SL g535 ( 
.A(n_251),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_72),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_68),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_61),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_167),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_304),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_1),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_115),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_214),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_205),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_0),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_238),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_51),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_186),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_219),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_280),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_141),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_53),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_199),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_195),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_257),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_30),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_80),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_302),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_226),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_66),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_114),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_125),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_56),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_154),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_250),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_149),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_473),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_351),
.B(n_0),
.Y(n_568)
);

CKINVDCx11_ASAP7_75t_R g569 ( 
.A(n_448),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_439),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_473),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_528),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_532),
.B(n_1),
.Y(n_573)
);

INVx6_ASAP7_75t_L g574 ( 
.A(n_340),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_366),
.B(n_2),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_343),
.B(n_2),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_343),
.B(n_3),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_473),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_470),
.B(n_4),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_363),
.B(n_547),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_473),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_384),
.B(n_5),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_386),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_503),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_503),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_470),
.B(n_6),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_483),
.B(n_7),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_528),
.B(n_7),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_503),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_503),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_402),
.B(n_8),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_511),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_386),
.B(n_9),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_485),
.B(n_9),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_544),
.B(n_553),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_441),
.B(n_10),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_487),
.B(n_11),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_439),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_544),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_553),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_439),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_439),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_511),
.B(n_12),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_443),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_483),
.B(n_13),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_443),
.B(n_13),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_447),
.B(n_14),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_447),
.B(n_14),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_455),
.B(n_15),
.Y(n_609)
);

BUFx8_ASAP7_75t_SL g610 ( 
.A(n_535),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_455),
.B(n_16),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_472),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_472),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_511),
.B(n_17),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_485),
.B(n_17),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_472),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_472),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_350),
.B(n_19),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_350),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_388),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_340),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_494),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_388),
.B(n_434),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_434),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_477),
.B(n_21),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_340),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_380),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_411),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_436),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_436),
.Y(n_630)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_436),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_371),
.B(n_22),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_477),
.B(n_23),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_438),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_502),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_365),
.B(n_25),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_494),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_509),
.B(n_25),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_481),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_502),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_518),
.B(n_26),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_502),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_494),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_341),
.B(n_27),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_369),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_538),
.B(n_342),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_562),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_391),
.B(n_28),
.Y(n_648)
);

INVx5_ASAP7_75t_L g649 ( 
.A(n_562),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_562),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_505),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_347),
.B(n_28),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_541),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_344),
.B(n_29),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_383),
.B(n_30),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_557),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_415),
.B(n_31),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_535),
.Y(n_658)
);

BUFx12f_ASAP7_75t_L g659 ( 
.A(n_349),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_372),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_425),
.B(n_33),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_457),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_378),
.B(n_33),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_382),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_482),
.B(n_35),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_389),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_400),
.B(n_35),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_410),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_412),
.B(n_36),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_416),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_546),
.B(n_37),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_494),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_423),
.B(n_37),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_336),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_368),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_424),
.B(n_38),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_359),
.B(n_377),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_494),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_426),
.B(n_39),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_427),
.B(n_39),
.Y(n_680)
);

BUFx12f_ASAP7_75t_L g681 ( 
.A(n_385),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_442),
.B(n_40),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_494),
.Y(n_683)
);

BUFx8_ASAP7_75t_SL g684 ( 
.A(n_448),
.Y(n_684)
);

AND2x6_ASAP7_75t_L g685 ( 
.A(n_432),
.B(n_93),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_437),
.B(n_42),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_453),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_460),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_464),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_494),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_467),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_491),
.B(n_42),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_387),
.B(n_43),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_504),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_338),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g696 ( 
.A(n_394),
.B(n_43),
.C(n_45),
.Y(n_696)
);

BUFx8_ASAP7_75t_SL g697 ( 
.A(n_469),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_507),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_517),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_524),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_534),
.B(n_46),
.Y(n_701)
);

NOR2x1_ASAP7_75t_L g702 ( 
.A(n_549),
.B(n_100),
.Y(n_702)
);

INVx5_ASAP7_75t_L g703 ( 
.A(n_395),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_456),
.B(n_47),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_551),
.B(n_47),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_554),
.Y(n_706)
);

BUFx12f_ASAP7_75t_L g707 ( 
.A(n_399),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_558),
.B(n_559),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_565),
.Y(n_709)
);

INVx5_ASAP7_75t_L g710 ( 
.A(n_404),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_498),
.B(n_48),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_405),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_339),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_406),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_408),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_345),
.B(n_48),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_413),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_346),
.B(n_49),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_414),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_348),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_421),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_352),
.B(n_354),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_355),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_422),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_357),
.B(n_49),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_430),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_601),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_598),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_601),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_677),
.B(n_358),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_610),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_591),
.A2(n_522),
.B1(n_560),
.B2(n_469),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_613),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_601),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_662),
.A2(n_452),
.B1(n_461),
.B2(n_451),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_570),
.Y(n_736)
);

OAI22xp33_ASAP7_75t_SL g737 ( 
.A1(n_629),
.A2(n_475),
.B1(n_486),
.B2(n_471),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_626),
.B(n_337),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_654),
.A2(n_353),
.B1(n_356),
.B2(n_337),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_661),
.A2(n_356),
.B1(n_398),
.B2(n_353),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_570),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_583),
.B(n_495),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_665),
.A2(n_403),
.B1(n_429),
.B2(n_398),
.Y(n_743)
);

AO22x2_ASAP7_75t_L g744 ( 
.A1(n_696),
.A2(n_54),
.B1(n_50),
.B2(n_52),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_717),
.B(n_360),
.Y(n_745)
);

OA22x2_ASAP7_75t_L g746 ( 
.A1(n_580),
.A2(n_497),
.B1(n_501),
.B2(n_496),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_671),
.A2(n_429),
.B1(n_431),
.B2(n_403),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_632),
.A2(n_476),
.B1(n_484),
.B2(n_431),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_674),
.B(n_566),
.Y(n_749)
);

OAI22xp33_ASAP7_75t_L g750 ( 
.A1(n_662),
.A2(n_510),
.B1(n_512),
.B2(n_506),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_602),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_602),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_612),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_573),
.A2(n_516),
.B1(n_519),
.B2(n_514),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_724),
.B(n_361),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_629),
.B(n_362),
.Y(n_756)
);

AO22x2_ASAP7_75t_L g757 ( 
.A1(n_696),
.A2(n_57),
.B1(n_50),
.B2(n_55),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_641),
.A2(n_484),
.B1(n_515),
.B2(n_476),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_568),
.A2(n_582),
.B1(n_596),
.B2(n_575),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_612),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_640),
.B(n_364),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_SL g762 ( 
.A1(n_626),
.A2(n_522),
.B1(n_560),
.B2(n_515),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_597),
.A2(n_523),
.B1(n_527),
.B2(n_520),
.Y(n_763)
);

AO22x2_ASAP7_75t_L g764 ( 
.A1(n_603),
.A2(n_58),
.B1(n_55),
.B2(n_57),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_616),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_640),
.B(n_367),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_635),
.B(n_370),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_571),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_642),
.B(n_373),
.Y(n_769)
);

BUFx10_ASAP7_75t_L g770 ( 
.A(n_574),
.Y(n_770)
);

XNOR2xp5_ASAP7_75t_L g771 ( 
.A(n_647),
.B(n_529),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_617),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_659),
.B(n_531),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_652),
.A2(n_536),
.B1(n_537),
.B2(n_533),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_655),
.A2(n_552),
.B1(n_556),
.B2(n_545),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_571),
.Y(n_776)
);

OA22x2_ASAP7_75t_L g777 ( 
.A1(n_646),
.A2(n_563),
.B1(n_375),
.B2(n_376),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_713),
.B(n_374),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_635),
.A2(n_381),
.B1(n_390),
.B2(n_379),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_712),
.B(n_58),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_571),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_578),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_642),
.B(n_392),
.Y(n_783)
);

AO22x2_ASAP7_75t_L g784 ( 
.A1(n_603),
.A2(n_62),
.B1(n_59),
.B2(n_60),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_657),
.A2(n_396),
.B1(n_397),
.B2(n_393),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_574),
.A2(n_407),
.B1(n_409),
.B2(n_401),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_712),
.B(n_59),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_682),
.A2(n_478),
.B1(n_561),
.B2(n_555),
.Y(n_788)
);

OAI22xp33_ASAP7_75t_SL g789 ( 
.A1(n_576),
.A2(n_564),
.B1(n_550),
.B2(n_548),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_715),
.B(n_417),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_715),
.B(n_418),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_721),
.B(n_419),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_704),
.A2(n_543),
.B1(n_542),
.B2(n_540),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_684),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_711),
.A2(n_466),
.B1(n_530),
.B2(n_526),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_714),
.A2(n_539),
.B1(n_525),
.B2(n_521),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_SL g797 ( 
.A(n_650),
.B(n_420),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_711),
.A2(n_513),
.B1(n_508),
.B2(n_500),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_681),
.A2(n_499),
.B1(n_493),
.B2(n_492),
.Y(n_799)
);

AO22x2_ASAP7_75t_L g800 ( 
.A1(n_614),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_726),
.B(n_428),
.Y(n_801)
);

OAI22xp33_ASAP7_75t_L g802 ( 
.A1(n_576),
.A2(n_490),
.B1(n_489),
.B2(n_488),
.Y(n_802)
);

AO22x2_ASAP7_75t_L g803 ( 
.A1(n_614),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_577),
.A2(n_480),
.B1(n_479),
.B2(n_474),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_719),
.B(n_572),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_621),
.B(n_433),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_578),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_578),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_577),
.A2(n_468),
.B1(n_465),
.B2(n_463),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_707),
.A2(n_462),
.B1(n_459),
.B2(n_458),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_713),
.B(n_435),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_579),
.A2(n_454),
.B1(n_450),
.B2(n_449),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_693),
.A2(n_445),
.B1(n_444),
.B2(n_440),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_579),
.A2(n_586),
.B1(n_605),
.B2(n_638),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_604),
.B(n_67),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_718),
.A2(n_446),
.B1(n_68),
.B2(n_69),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_713),
.B(n_67),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_604),
.B(n_69),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_581),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_586),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_587),
.A2(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_581),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_725),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_621),
.B(n_81),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_675),
.B(n_599),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_587),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_621),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_581),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_805),
.B(n_658),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_756),
.B(n_720),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_761),
.B(n_658),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_781),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_742),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_781),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_822),
.Y(n_835)
);

XNOR2xp5_ASAP7_75t_L g836 ( 
.A(n_732),
.B(n_739),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_822),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_732),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_728),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_825),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_766),
.B(n_658),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_794),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_814),
.B(n_759),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_768),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_770),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_768),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_740),
.Y(n_847)
);

XOR2xp5_ASAP7_75t_L g848 ( 
.A(n_743),
.B(n_722),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_828),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_828),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_776),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_745),
.B(n_720),
.Y(n_852)
);

OR2x6_ASAP7_75t_L g853 ( 
.A(n_764),
.B(n_606),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_755),
.B(n_720),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_769),
.B(n_723),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_783),
.B(n_630),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_782),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_807),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_729),
.Y(n_859)
);

INVxp33_ASAP7_75t_L g860 ( 
.A(n_771),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_808),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_819),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_790),
.B(n_595),
.Y(n_863)
);

INVxp33_ASAP7_75t_L g864 ( 
.A(n_747),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_748),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_762),
.Y(n_866)
);

XOR2x2_ASAP7_75t_L g867 ( 
.A(n_758),
.B(n_697),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_727),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_727),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_734),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_733),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_772),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_729),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_741),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_791),
.B(n_595),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_751),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_752),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_770),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_753),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_760),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_778),
.A2(n_623),
.B(n_590),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_736),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_736),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_765),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_754),
.B(n_722),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_765),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_817),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_749),
.B(n_723),
.Y(n_888)
);

NOR2xp67_ASAP7_75t_L g889 ( 
.A(n_785),
.B(n_630),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_730),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_792),
.B(n_630),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_815),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_818),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_801),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_777),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_797),
.B(n_723),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_780),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_811),
.B(n_695),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_821),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_806),
.B(n_567),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_787),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_R g902 ( 
.A(n_773),
.B(n_588),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_746),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_824),
.Y(n_904)
);

XOR2xp5_ASAP7_75t_L g905 ( 
.A(n_731),
.B(n_675),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_788),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_826),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_764),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_827),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_784),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_800),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_767),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_800),
.Y(n_913)
);

XOR2xp5_ASAP7_75t_L g914 ( 
.A(n_799),
.B(n_716),
.Y(n_914)
);

CKINVDCx16_ASAP7_75t_R g915 ( 
.A(n_798),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_803),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_803),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_796),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_802),
.A2(n_623),
.B(n_590),
.Y(n_919)
);

INVxp33_ASAP7_75t_L g920 ( 
.A(n_738),
.Y(n_920)
);

NAND2x1p5_ASAP7_75t_L g921 ( 
.A(n_863),
.B(n_702),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_884),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_859),
.Y(n_923)
);

AND2x2_ASAP7_75t_SL g924 ( 
.A(n_843),
.B(n_821),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_863),
.B(n_798),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_886),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_884),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_888),
.B(n_793),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_839),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_875),
.B(n_708),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_840),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_888),
.B(n_804),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_839),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_912),
.B(n_795),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_871),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_875),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_843),
.B(n_708),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_830),
.A2(n_813),
.B(n_812),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_833),
.B(n_779),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_895),
.B(n_588),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_896),
.B(n_890),
.Y(n_941)
);

BUFx4f_ASAP7_75t_L g942 ( 
.A(n_885),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_887),
.B(n_763),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_894),
.B(n_593),
.Y(n_944)
);

AND2x2_ASAP7_75t_SL g945 ( 
.A(n_915),
.B(n_618),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_882),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_871),
.Y(n_947)
);

AND2x2_ASAP7_75t_SL g948 ( 
.A(n_906),
.B(n_618),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_883),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_872),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_859),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_892),
.B(n_594),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_852),
.B(n_685),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_903),
.B(n_644),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_852),
.B(n_685),
.Y(n_955)
);

BUFx4f_ASAP7_75t_L g956 ( 
.A(n_918),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_855),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_832),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_834),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_904),
.B(n_644),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_835),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_909),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_854),
.B(n_685),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_893),
.B(n_615),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_837),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_909),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_854),
.B(n_685),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_897),
.B(n_679),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_840),
.B(n_774),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_874),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_898),
.A2(n_809),
.B(n_789),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_901),
.B(n_679),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_856),
.B(n_636),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_868),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_899),
.B(n_680),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_907),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_908),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_878),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_891),
.B(n_896),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_831),
.B(n_636),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_869),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_899),
.B(n_680),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_841),
.B(n_775),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_910),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_853),
.B(n_627),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_876),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_851),
.B(n_633),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_842),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_853),
.B(n_627),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_857),
.B(n_633),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_905),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_909),
.Y(n_992)
);

BUFx4_ASAP7_75t_SL g993 ( 
.A(n_838),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_914),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_909),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_919),
.A2(n_605),
.B(n_638),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_877),
.Y(n_997)
);

INVxp67_ASAP7_75t_SL g998 ( 
.A(n_879),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_920),
.B(n_810),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_853),
.B(n_656),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_829),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_848),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_889),
.B(n_786),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_845),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_920),
.B(n_656),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_900),
.B(n_619),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_880),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_858),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_861),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_862),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_881),
.B(n_619),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_870),
.B(n_620),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_844),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_846),
.B(n_620),
.Y(n_1014)
);

AND2x6_ASAP7_75t_L g1015 ( 
.A(n_911),
.B(n_823),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_925),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_957),
.B(n_913),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_957),
.B(n_916),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_922),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_928),
.B(n_864),
.Y(n_1020)
);

AND2x2_ASAP7_75t_SL g1021 ( 
.A(n_924),
.B(n_865),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_925),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1005),
.B(n_864),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_SL g1024 ( 
.A(n_924),
.B(n_866),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_957),
.B(n_937),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_957),
.B(n_917),
.Y(n_1026)
);

BUFx8_ASAP7_75t_L g1027 ( 
.A(n_985),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_922),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_936),
.B(n_849),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_SL g1030 ( 
.A(n_948),
.B(n_866),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_936),
.B(n_773),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_923),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_931),
.B(n_969),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_934),
.B(n_860),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_988),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_922),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_948),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_927),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1005),
.B(n_860),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_975),
.B(n_850),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_939),
.B(n_847),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_976),
.B(n_847),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_975),
.B(n_873),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_SL g1044 ( 
.A(n_945),
.B(n_942),
.Y(n_1044)
);

INVx5_ASAP7_75t_L g1045 ( 
.A(n_992),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_957),
.B(n_744),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_988),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_923),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_927),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_927),
.Y(n_1050)
);

NAND2x1p5_ASAP7_75t_L g1051 ( 
.A(n_962),
.B(n_599),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_929),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_929),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_945),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_1015),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_982),
.B(n_628),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_933),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_937),
.B(n_744),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_1015),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_933),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_992),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_969),
.B(n_836),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_935),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_982),
.B(n_634),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_992),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_1015),
.Y(n_1066)
);

NAND2x1_ASAP7_75t_SL g1067 ( 
.A(n_999),
.B(n_816),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_935),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_932),
.B(n_757),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_1001),
.B(n_639),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_956),
.B(n_569),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_923),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_947),
.Y(n_1073)
);

INVx6_ASAP7_75t_L g1074 ( 
.A(n_954),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_943),
.B(n_631),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_SL g1076 ( 
.A(n_942),
.B(n_820),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_979),
.B(n_757),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_962),
.B(n_599),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_1001),
.B(n_651),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_977),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_996),
.B(n_737),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_1001),
.B(n_653),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_956),
.B(n_735),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_943),
.B(n_620),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_952),
.B(n_631),
.Y(n_1085)
);

NAND2x1_ASAP7_75t_L g1086 ( 
.A(n_992),
.B(n_622),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_1015),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_984),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_923),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_968),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_949),
.B(n_624),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_968),
.Y(n_1092)
);

BUFx12f_ASAP7_75t_L g1093 ( 
.A(n_1015),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1008),
.B(n_653),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_947),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_966),
.B(n_923),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_951),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_952),
.B(n_649),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_978),
.B(n_867),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_992),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1008),
.B(n_606),
.Y(n_1101)
);

INVx5_ASAP7_75t_L g1102 ( 
.A(n_1045),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1057),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_1080),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1073),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_1045),
.Y(n_1106)
);

CKINVDCx11_ASAP7_75t_R g1107 ( 
.A(n_1035),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1097),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_1039),
.Y(n_1109)
);

INVx3_ASAP7_75t_SL g1110 ( 
.A(n_1031),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_1074),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1047),
.Y(n_1112)
);

CKINVDCx16_ASAP7_75t_R g1113 ( 
.A(n_1030),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_1027),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1095),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_1054),
.Y(n_1116)
);

INVx6_ASAP7_75t_L g1117 ( 
.A(n_1032),
.Y(n_1117)
);

INVx8_ASAP7_75t_L g1118 ( 
.A(n_1045),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1052),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1053),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1060),
.Y(n_1121)
);

BUFx12f_ASAP7_75t_L g1122 ( 
.A(n_1031),
.Y(n_1122)
);

BUFx2_ASAP7_75t_SL g1123 ( 
.A(n_1094),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_1061),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1061),
.Y(n_1125)
);

INVx3_ASAP7_75t_SL g1126 ( 
.A(n_1031),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_1033),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1097),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1063),
.Y(n_1129)
);

BUFx2_ASAP7_75t_SL g1130 ( 
.A(n_1082),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1023),
.B(n_944),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_1088),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_1061),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1093),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1055),
.B(n_921),
.Y(n_1135)
);

BUFx5_ASAP7_75t_L g1136 ( 
.A(n_1019),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_1032),
.Y(n_1137)
);

BUFx12f_ASAP7_75t_L g1138 ( 
.A(n_1062),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_1099),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1068),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1049),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1016),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1050),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1028),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1032),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1059),
.B(n_926),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1017),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1048),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1048),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1020),
.B(n_1069),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1022),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1017),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1018),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_1066),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1048),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_1072),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1072),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1087),
.Y(n_1158)
);

BUFx12f_ASAP7_75t_L g1159 ( 
.A(n_1082),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1018),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_1072),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1089),
.Y(n_1162)
);

INVx5_ASAP7_75t_L g1163 ( 
.A(n_1089),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1021),
.A2(n_942),
.B1(n_983),
.B2(n_941),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1026),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1089),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_1065),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_1074),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1026),
.Y(n_1169)
);

INVx6_ASAP7_75t_SL g1170 ( 
.A(n_1056),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1046),
.Y(n_1171)
);

CKINVDCx16_ASAP7_75t_R g1172 ( 
.A(n_1112),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1129),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1129),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1150),
.A2(n_1041),
.B1(n_1024),
.B2(n_1030),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1140),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1119),
.Y(n_1177)
);

BUFx8_ASAP7_75t_L g1178 ( 
.A(n_1159),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1120),
.Y(n_1179)
);

CKINVDCx11_ASAP7_75t_R g1180 ( 
.A(n_1107),
.Y(n_1180)
);

BUFx8_ASAP7_75t_L g1181 ( 
.A(n_1159),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1113),
.A2(n_1139),
.B1(n_1034),
.B2(n_1042),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1104),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_1109),
.B(n_1077),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1121),
.Y(n_1185)
);

INVx5_ASAP7_75t_L g1186 ( 
.A(n_1118),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1125),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1134),
.B(n_1090),
.Y(n_1188)
);

CKINVDCx11_ASAP7_75t_R g1189 ( 
.A(n_1107),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1103),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1150),
.A2(n_1024),
.B1(n_1076),
.B2(n_1037),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1164),
.A2(n_1069),
.B1(n_1058),
.B2(n_1077),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1171),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1131),
.A2(n_1076),
.B1(n_1037),
.B2(n_1083),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1138),
.A2(n_1044),
.B1(n_1071),
.B2(n_956),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1146),
.A2(n_1015),
.B1(n_938),
.B2(n_1064),
.Y(n_1196)
);

OAI22xp33_ASAP7_75t_R g1197 ( 
.A1(n_1127),
.A2(n_991),
.B1(n_1132),
.B2(n_902),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1146),
.A2(n_1064),
.B1(n_1044),
.B2(n_1092),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_1116),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1147),
.A2(n_1025),
.B1(n_1046),
.B2(n_1084),
.Y(n_1200)
);

CKINVDCx11_ASAP7_75t_R g1201 ( 
.A(n_1114),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1138),
.A2(n_994),
.B1(n_1081),
.B2(n_971),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1125),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1139),
.A2(n_1075),
.B1(n_1067),
.B2(n_985),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1152),
.A2(n_1025),
.B1(n_1084),
.B2(n_1101),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1103),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1151),
.Y(n_1207)
);

INVx11_ASAP7_75t_L g1208 ( 
.A(n_1154),
.Y(n_1208)
);

BUFx8_ASAP7_75t_L g1209 ( 
.A(n_1114),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1151),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1105),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1153),
.A2(n_1101),
.B1(n_1043),
.B2(n_1040),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1105),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1115),
.Y(n_1214)
);

CKINVDCx11_ASAP7_75t_R g1215 ( 
.A(n_1122),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1160),
.B(n_1165),
.Y(n_1216)
);

OAI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1142),
.A2(n_1002),
.B1(n_902),
.B2(n_1004),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1115),
.Y(n_1218)
);

BUFx12f_ASAP7_75t_L g1219 ( 
.A(n_1104),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1130),
.A2(n_989),
.B1(n_1000),
.B2(n_1085),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1169),
.A2(n_1135),
.B1(n_1158),
.B2(n_1102),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1142),
.A2(n_1079),
.B1(n_1070),
.B2(n_1043),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1158),
.A2(n_1070),
.B1(n_1040),
.B2(n_989),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1116),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1144),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1123),
.A2(n_1000),
.B1(n_972),
.B2(n_980),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1154),
.Y(n_1227)
);

INVx5_ASAP7_75t_L g1228 ( 
.A(n_1118),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1170),
.A2(n_1098),
.B1(n_930),
.B2(n_940),
.Y(n_1229)
);

CKINVDCx11_ASAP7_75t_R g1230 ( 
.A(n_1122),
.Y(n_1230)
);

CKINVDCx11_ASAP7_75t_R g1231 ( 
.A(n_1110),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_1134),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1110),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1135),
.A2(n_973),
.B1(n_1096),
.B2(n_955),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1126),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1170),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1144),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1111),
.B(n_964),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1175),
.A2(n_607),
.B1(n_609),
.B2(n_608),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1182),
.A2(n_607),
.B1(n_609),
.B2(n_608),
.Y(n_1240)
);

BUFx12f_ASAP7_75t_L g1241 ( 
.A(n_1180),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1177),
.Y(n_1242)
);

BUFx4f_ASAP7_75t_SL g1243 ( 
.A(n_1219),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1182),
.A2(n_611),
.B1(n_667),
.B2(n_663),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1207),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1191),
.A2(n_611),
.B1(n_667),
.B2(n_663),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1202),
.A2(n_750),
.B(n_1003),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1194),
.A2(n_669),
.B1(n_676),
.B2(n_673),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1197),
.A2(n_669),
.B1(n_676),
.B2(n_673),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1210),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1192),
.A2(n_686),
.B1(n_701),
.B2(n_692),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1192),
.A2(n_686),
.B1(n_701),
.B2(n_692),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1204),
.A2(n_705),
.B1(n_648),
.B2(n_625),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1179),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1226),
.A2(n_1126),
.B1(n_649),
.B2(n_1135),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_SL g1256 ( 
.A1(n_1195),
.A2(n_648),
.B(n_930),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1196),
.A2(n_1135),
.B1(n_1010),
.B2(n_946),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1186),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1186),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1212),
.A2(n_1170),
.B1(n_1168),
.B2(n_1111),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1178),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1220),
.A2(n_1168),
.B1(n_960),
.B2(n_964),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1198),
.A2(n_1010),
.B1(n_949),
.B2(n_1007),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1208),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1222),
.A2(n_921),
.B1(n_1102),
.B2(n_981),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1217),
.B(n_1102),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1216),
.B(n_972),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1190),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1199),
.A2(n_649),
.B1(n_993),
.B2(n_1118),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1223),
.A2(n_921),
.B1(n_1102),
.B2(n_981),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1224),
.A2(n_1118),
.B1(n_716),
.B2(n_1136),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1189),
.Y(n_1272)
);

NOR2x1_ASAP7_75t_SL g1273 ( 
.A(n_1186),
.B(n_1102),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1187),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1185),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1184),
.B(n_997),
.Y(n_1276)
);

AOI222xp33_ASAP7_75t_L g1277 ( 
.A1(n_1238),
.A2(n_940),
.B1(n_954),
.B2(n_960),
.C1(n_691),
.C2(n_709),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1229),
.A2(n_965),
.B1(n_953),
.B2(n_963),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1193),
.B(n_940),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_L g1280 ( 
.A(n_1205),
.B(n_970),
.C(n_997),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1214),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1183),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1200),
.A2(n_986),
.B1(n_990),
.B2(n_987),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1231),
.A2(n_1235),
.B1(n_1221),
.B2(n_1233),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1173),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1174),
.A2(n_600),
.B1(n_959),
.B2(n_958),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1227),
.A2(n_960),
.B(n_954),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1172),
.B(n_1029),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1176),
.B(n_1029),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1225),
.B(n_998),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1237),
.A2(n_1206),
.B1(n_1213),
.B2(n_1211),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1218),
.A2(n_600),
.B1(n_959),
.B2(n_958),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1187),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1187),
.Y(n_1294)
);

OAI21xp33_ASAP7_75t_L g1295 ( 
.A1(n_1188),
.A2(n_986),
.B(n_1091),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1203),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1221),
.A2(n_967),
.B1(n_951),
.B2(n_1051),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1188),
.B(n_987),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1178),
.A2(n_1136),
.B1(n_1167),
.B2(n_1125),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1236),
.B(n_987),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1234),
.A2(n_600),
.B1(n_974),
.B2(n_961),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1228),
.A2(n_951),
.B1(n_1078),
.B2(n_1167),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1228),
.A2(n_1167),
.B1(n_961),
.B2(n_974),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1215),
.A2(n_1009),
.B1(n_664),
.B2(n_698),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1244),
.A2(n_1230),
.B1(n_1232),
.B2(n_1201),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1270),
.A2(n_1181),
.B1(n_1209),
.B2(n_1228),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1285),
.B(n_1141),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1276),
.B(n_1141),
.Y(n_1308)
);

OAI222xp33_ASAP7_75t_L g1309 ( 
.A1(n_1240),
.A2(n_1143),
.B1(n_1128),
.B2(n_1108),
.C1(n_950),
.C2(n_1006),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1242),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1254),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1265),
.A2(n_1136),
.B1(n_1203),
.B2(n_1125),
.Y(n_1312)
);

NAND3xp33_ASAP7_75t_L g1313 ( 
.A(n_1247),
.B(n_1252),
.C(n_1251),
.Y(n_1313)
);

OAI21xp33_ASAP7_75t_L g1314 ( 
.A1(n_1240),
.A2(n_990),
.B(n_1012),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1253),
.A2(n_1251),
.B1(n_1252),
.B2(n_1248),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1260),
.A2(n_1136),
.B1(n_1203),
.B2(n_1125),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_SL g1317 ( 
.A1(n_1267),
.A2(n_1136),
.B1(n_592),
.B2(n_1163),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1249),
.B(n_1239),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_L g1319 ( 
.A(n_1246),
.B(n_660),
.C(n_645),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1249),
.A2(n_1013),
.B1(n_1128),
.B2(n_1136),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1239),
.A2(n_1013),
.B1(n_1136),
.B2(n_966),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1271),
.A2(n_1117),
.B1(n_1106),
.B2(n_1133),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1245),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1255),
.A2(n_700),
.B1(n_694),
.B2(n_699),
.Y(n_1324)
);

NOR3xp33_ASAP7_75t_L g1325 ( 
.A(n_1287),
.B(n_1011),
.C(n_1156),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1284),
.A2(n_1117),
.B1(n_1106),
.B2(n_1124),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1275),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1262),
.A2(n_1156),
.B1(n_1163),
.B2(n_1161),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1268),
.B(n_1145),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1281),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1266),
.A2(n_1036),
.B1(n_1038),
.B2(n_1014),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1256),
.A2(n_660),
.B(n_645),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1277),
.A2(n_1166),
.B1(n_1145),
.B2(n_1155),
.Y(n_1333)
);

AOI221xp5_ASAP7_75t_L g1334 ( 
.A1(n_1304),
.A2(n_668),
.B1(n_689),
.B2(n_688),
.C(n_687),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1280),
.A2(n_592),
.B1(n_1163),
.B2(n_1161),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1288),
.A2(n_592),
.B1(n_1163),
.B2(n_1161),
.Y(n_1336)
);

AOI221xp5_ASAP7_75t_L g1337 ( 
.A1(n_1304),
.A2(n_670),
.B1(n_687),
.B2(n_706),
.C(n_689),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1300),
.A2(n_703),
.B1(n_710),
.B2(n_1117),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1257),
.A2(n_1166),
.B1(n_1155),
.B2(n_660),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1283),
.A2(n_666),
.B1(n_706),
.B2(n_688),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1295),
.A2(n_666),
.B1(n_706),
.B2(n_688),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1291),
.B(n_1137),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1250),
.A2(n_1163),
.B1(n_1161),
.B2(n_1162),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1269),
.A2(n_1117),
.B1(n_1124),
.B2(n_1106),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1289),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1261),
.A2(n_670),
.B1(n_687),
.B2(n_689),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_L g1347 ( 
.A(n_1263),
.B(n_1298),
.C(n_1279),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1291),
.B(n_1137),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1278),
.A2(n_1301),
.B1(n_1282),
.B2(n_1243),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1243),
.A2(n_703),
.B1(n_710),
.B2(n_995),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1290),
.B(n_1137),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1293),
.B(n_1294),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1241),
.A2(n_995),
.B1(n_1162),
.B2(n_1157),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1297),
.A2(n_1161),
.B1(n_1162),
.B2(n_1157),
.Y(n_1354)
);

AO22x1_ASAP7_75t_L g1355 ( 
.A1(n_1258),
.A2(n_1162),
.B1(n_1157),
.B2(n_1149),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1296),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1286),
.A2(n_1124),
.B1(n_1133),
.B2(n_1100),
.Y(n_1357)
);

OAI222xp33_ASAP7_75t_L g1358 ( 
.A1(n_1299),
.A2(n_1086),
.B1(n_683),
.B2(n_690),
.C1(n_637),
.C2(n_643),
.Y(n_1358)
);

OAI221xp5_ASAP7_75t_L g1359 ( 
.A1(n_1286),
.A2(n_1133),
.B1(n_1065),
.B2(n_1100),
.C(n_624),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1292),
.A2(n_995),
.B1(n_1162),
.B2(n_1149),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1274),
.B(n_1148),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1273),
.A2(n_1157),
.B1(n_1149),
.B2(n_1148),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1303),
.A2(n_1157),
.B1(n_1149),
.B2(n_1148),
.Y(n_1363)
);

AOI221xp5_ASAP7_75t_L g1364 ( 
.A1(n_1313),
.A2(n_624),
.B1(n_1292),
.B2(n_1302),
.C(n_1272),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_L g1365 ( 
.A(n_1315),
.B(n_1259),
.C(n_1258),
.Y(n_1365)
);

OAI221xp5_ASAP7_75t_L g1366 ( 
.A1(n_1305),
.A2(n_1264),
.B1(n_1259),
.B2(n_1274),
.C(n_1149),
.Y(n_1366)
);

AND2x2_ASAP7_75t_SL g1367 ( 
.A(n_1318),
.B(n_1274),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1310),
.B(n_1274),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1310),
.B(n_82),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1345),
.B(n_86),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1345),
.B(n_87),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1311),
.B(n_1327),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1323),
.B(n_87),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1359),
.A2(n_1148),
.B(n_678),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1311),
.B(n_88),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1332),
.A2(n_678),
.B(n_672),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1347),
.B(n_88),
.Y(n_1377)
);

AND2x2_ASAP7_75t_SL g1378 ( 
.A(n_1349),
.B(n_584),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1330),
.B(n_90),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1314),
.A2(n_678),
.B1(n_672),
.B2(n_90),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1327),
.B(n_91),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1352),
.B(n_91),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1342),
.B(n_585),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1342),
.B(n_585),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1330),
.B(n_589),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1308),
.B(n_589),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1307),
.B(n_101),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1307),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1356),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1319),
.A2(n_590),
.B1(n_567),
.B2(n_107),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1348),
.B(n_102),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1329),
.B(n_105),
.Y(n_1393)
);

OAI221xp5_ASAP7_75t_L g1394 ( 
.A1(n_1338),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.C(n_121),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1329),
.B(n_122),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1348),
.B(n_123),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1312),
.B(n_1306),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1350),
.B(n_567),
.C(n_134),
.Y(n_1398)
);

NOR3xp33_ASAP7_75t_L g1399 ( 
.A(n_1326),
.B(n_131),
.C(n_135),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1316),
.B(n_136),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1354),
.B(n_1320),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1317),
.B(n_138),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1346),
.A2(n_142),
.B(n_151),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1361),
.B(n_156),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1336),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1322),
.A2(n_177),
.B1(n_178),
.B2(n_181),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1324),
.B(n_187),
.C(n_190),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1363),
.B(n_191),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1325),
.A2(n_192),
.B(n_197),
.Y(n_1409)
);

NOR3xp33_ASAP7_75t_L g1410 ( 
.A(n_1377),
.B(n_1344),
.C(n_1309),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1372),
.Y(n_1411)
);

NOR3xp33_ASAP7_75t_L g1412 ( 
.A(n_1377),
.B(n_1328),
.C(n_1337),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1390),
.B(n_1388),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1388),
.B(n_1362),
.Y(n_1414)
);

NAND4xp75_ASAP7_75t_L g1415 ( 
.A(n_1409),
.B(n_1334),
.C(n_1353),
.D(n_1343),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1368),
.B(n_1355),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1380),
.A2(n_1340),
.B1(n_1339),
.B2(n_1335),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1368),
.B(n_1355),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1389),
.B(n_1321),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_L g1420 ( 
.A(n_1365),
.B(n_1333),
.C(n_1341),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1367),
.B(n_1360),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1383),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1397),
.A2(n_1331),
.B1(n_1357),
.B2(n_1358),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1385),
.A2(n_203),
.B(n_206),
.Y(n_1424)
);

NOR3xp33_ASAP7_75t_L g1425 ( 
.A(n_1366),
.B(n_209),
.C(n_210),
.Y(n_1425)
);

NOR3xp33_ASAP7_75t_L g1426 ( 
.A(n_1394),
.B(n_211),
.C(n_212),
.Y(n_1426)
);

AND2x4_ASAP7_75t_SL g1427 ( 
.A(n_1383),
.B(n_335),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1399),
.A2(n_213),
.B1(n_216),
.B2(n_217),
.Y(n_1428)
);

NOR3xp33_ASAP7_75t_L g1429 ( 
.A(n_1398),
.B(n_218),
.C(n_220),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1367),
.B(n_221),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1384),
.B(n_1369),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1384),
.B(n_222),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1381),
.B(n_223),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1381),
.B(n_225),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1392),
.B(n_231),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1373),
.B(n_237),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1379),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1375),
.Y(n_1438)
);

NOR2x1_ASAP7_75t_L g1439 ( 
.A(n_1370),
.B(n_239),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1371),
.B(n_1382),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1386),
.B(n_241),
.Y(n_1441)
);

NAND4xp75_ASAP7_75t_L g1442 ( 
.A(n_1378),
.B(n_247),
.C(n_253),
.D(n_254),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1401),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1443),
.B(n_1431),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1411),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1413),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1413),
.B(n_1396),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1422),
.B(n_1392),
.Y(n_1448)
);

NAND4xp75_ASAP7_75t_L g1449 ( 
.A(n_1439),
.B(n_1400),
.C(n_1408),
.D(n_1402),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1427),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1437),
.Y(n_1451)
);

NOR3xp33_ASAP7_75t_L g1452 ( 
.A(n_1442),
.B(n_1412),
.C(n_1415),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1440),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1416),
.B(n_1401),
.Y(n_1454)
);

XOR2x2_ASAP7_75t_L g1455 ( 
.A(n_1443),
.B(n_1378),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1440),
.Y(n_1456)
);

NAND4xp75_ASAP7_75t_L g1457 ( 
.A(n_1430),
.B(n_1400),
.C(n_1408),
.D(n_1402),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1437),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1416),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1431),
.B(n_1387),
.Y(n_1460)
);

NAND4xp75_ASAP7_75t_L g1461 ( 
.A(n_1430),
.B(n_1364),
.C(n_1376),
.D(n_1393),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1438),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1418),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1418),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1414),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1423),
.A2(n_1406),
.B1(n_1391),
.B2(n_1403),
.Y(n_1466)
);

NAND4xp75_ASAP7_75t_L g1467 ( 
.A(n_1421),
.B(n_1376),
.C(n_1395),
.D(n_1404),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1436),
.B(n_1376),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1414),
.Y(n_1469)
);

XNOR2xp5_ASAP7_75t_L g1470 ( 
.A(n_1435),
.B(n_1405),
.Y(n_1470)
);

XOR2x2_ASAP7_75t_L g1471 ( 
.A(n_1457),
.B(n_1442),
.Y(n_1471)
);

AO22x2_ASAP7_75t_L g1472 ( 
.A1(n_1452),
.A2(n_1415),
.B1(n_1410),
.B2(n_1425),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1454),
.Y(n_1473)
);

OA22x2_ASAP7_75t_L g1474 ( 
.A1(n_1454),
.A2(n_1427),
.B1(n_1433),
.B2(n_1434),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1465),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1458),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1462),
.Y(n_1477)
);

XNOR2xp5_ASAP7_75t_L g1478 ( 
.A(n_1455),
.B(n_1470),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1465),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1451),
.Y(n_1480)
);

INVxp33_ASAP7_75t_L g1481 ( 
.A(n_1468),
.Y(n_1481)
);

XOR2x2_ASAP7_75t_L g1482 ( 
.A(n_1452),
.B(n_1420),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_1469),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1459),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1459),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1466),
.A2(n_1426),
.B1(n_1429),
.B2(n_1421),
.Y(n_1486)
);

XNOR2x2_ASAP7_75t_L g1487 ( 
.A(n_1449),
.B(n_1432),
.Y(n_1487)
);

XNOR2x1_ASAP7_75t_L g1488 ( 
.A(n_1466),
.B(n_1435),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1445),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1463),
.B(n_1419),
.Y(n_1490)
);

OA22x2_ASAP7_75t_L g1491 ( 
.A1(n_1478),
.A2(n_1464),
.B1(n_1463),
.B2(n_1453),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1473),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1471),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1477),
.Y(n_1494)
);

INVxp33_ASAP7_75t_SL g1495 ( 
.A(n_1486),
.Y(n_1495)
);

XOR2x2_ASAP7_75t_L g1496 ( 
.A(n_1482),
.B(n_1456),
.Y(n_1496)
);

AOI22x1_ASAP7_75t_L g1497 ( 
.A1(n_1472),
.A2(n_1487),
.B1(n_1484),
.B2(n_1479),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1472),
.A2(n_1468),
.B1(n_1461),
.B2(n_1467),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1489),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1483),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1472),
.A2(n_1464),
.B1(n_1450),
.B2(n_1419),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1483),
.Y(n_1502)
);

OA22x2_ASAP7_75t_L g1503 ( 
.A1(n_1475),
.A2(n_1450),
.B1(n_1444),
.B2(n_1446),
.Y(n_1503)
);

AOI22x1_ASAP7_75t_L g1504 ( 
.A1(n_1484),
.A2(n_1432),
.B1(n_1441),
.B2(n_1460),
.Y(n_1504)
);

XNOR2x1_ASAP7_75t_L g1505 ( 
.A(n_1488),
.B(n_1447),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1474),
.A2(n_1448),
.B1(n_1417),
.B2(n_1441),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1490),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1492),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1497),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1494),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1497),
.Y(n_1511)
);

OAI322xp33_ASAP7_75t_L g1512 ( 
.A1(n_1498),
.A2(n_1485),
.A3(n_1474),
.B1(n_1476),
.B2(n_1481),
.C1(n_1480),
.C2(n_1374),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1507),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1500),
.Y(n_1514)
);

INVxp67_ASAP7_75t_SL g1515 ( 
.A(n_1496),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1499),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1502),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1504),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1508),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1513),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1510),
.Y(n_1521)
);

NAND4xp25_ASAP7_75t_L g1522 ( 
.A(n_1509),
.B(n_1495),
.C(n_1501),
.D(n_1506),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1509),
.A2(n_1493),
.B1(n_1491),
.B2(n_1503),
.Y(n_1523)
);

BUFx4_ASAP7_75t_R g1524 ( 
.A(n_1511),
.Y(n_1524)
);

OAI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1522),
.A2(n_1515),
.B1(n_1511),
.B2(n_1518),
.C(n_1505),
.Y(n_1525)
);

O2A1O1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1520),
.A2(n_1518),
.B(n_1512),
.C(n_1514),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1519),
.Y(n_1527)
);

OAI22x1_ASAP7_75t_L g1528 ( 
.A1(n_1523),
.A2(n_1504),
.B1(n_1517),
.B2(n_1516),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1521),
.Y(n_1529)
);

NOR4xp25_ASAP7_75t_L g1530 ( 
.A(n_1525),
.B(n_1524),
.C(n_1428),
.D(n_1407),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1526),
.Y(n_1531)
);

NOR2x1_ASAP7_75t_L g1532 ( 
.A(n_1527),
.B(n_1424),
.Y(n_1532)
);

NOR2x1_ASAP7_75t_L g1533 ( 
.A(n_1529),
.B(n_1424),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1528),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1534),
.B(n_255),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1531),
.B(n_256),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1530),
.A2(n_258),
.B1(n_259),
.B2(n_262),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1537),
.A2(n_1532),
.B1(n_1533),
.B2(n_267),
.Y(n_1538)
);

NAND4xp25_ASAP7_75t_L g1539 ( 
.A(n_1536),
.B(n_263),
.C(n_264),
.D(n_270),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1535),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1538),
.A2(n_275),
.B1(n_277),
.B2(n_279),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1539),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1540),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1540),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1542),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1543),
.A2(n_286),
.B1(n_291),
.B2(n_292),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1544),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1541),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1547),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1548),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1545),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1551),
.A2(n_1546),
.B1(n_298),
.B2(n_299),
.Y(n_1552)
);

AOI221xp5_ASAP7_75t_L g1553 ( 
.A1(n_1550),
.A2(n_296),
.B1(n_303),
.B2(n_305),
.C(n_306),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1552),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1553),
.Y(n_1555)
);

AOI22x1_ASAP7_75t_L g1556 ( 
.A1(n_1554),
.A2(n_1549),
.B1(n_310),
.B2(n_311),
.Y(n_1556)
);

AOI22x1_ASAP7_75t_L g1557 ( 
.A1(n_1555),
.A2(n_1549),
.B1(n_314),
.B2(n_316),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1557),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1556),
.Y(n_1559)
);

OAI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1559),
.A2(n_317),
.B1(n_319),
.B2(n_321),
.C(n_322),
.Y(n_1560)
);

AOI211xp5_ASAP7_75t_L g1561 ( 
.A1(n_1560),
.A2(n_1558),
.B(n_325),
.C(n_328),
.Y(n_1561)
);


endmodule