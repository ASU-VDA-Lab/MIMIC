module fake_ibex_220_n_1139 (n_151, n_147, n_85, n_167, n_128, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1139);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1139;

wire n_1084;
wire n_599;
wire n_822;
wire n_778;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_418;
wire n_256;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_991;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_457;
wire n_412;
wire n_357;
wire n_494;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1044;
wire n_1018;
wire n_1106;
wire n_1129;
wire n_449;
wire n_1131;
wire n_547;
wire n_1134;
wire n_727;
wire n_1138;
wire n_1077;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_375;
wire n_280;
wire n_340;
wire n_317;
wire n_708;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_327;
wire n_326;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_339;
wire n_470;
wire n_276;
wire n_770;
wire n_965;
wire n_348;
wire n_1109;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_497;
wire n_711;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1112;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_1055;
wire n_732;
wire n_673;
wire n_832;
wire n_798;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1057;
wire n_1068;
wire n_325;
wire n_496;
wire n_301;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_787;
wire n_694;
wire n_977;
wire n_1075;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_569;
wire n_321;
wire n_600;
wire n_907;
wire n_933;
wire n_1081;
wire n_279;
wire n_1037;
wire n_374;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1101;
wire n_518;
wire n_367;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_1082;
wire n_1137;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_759;
wire n_917;
wire n_388;
wire n_968;
wire n_625;
wire n_953;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1028;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_300;
wire n_1135;
wire n_973;
wire n_358;
wire n_771;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1092;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_433;
wire n_262;
wire n_299;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_1054;
wire n_918;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_721;
wire n_365;
wire n_651;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1049;
wire n_1086;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_444;
wire n_564;
wire n_562;
wire n_506;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_1118;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_744;
wire n_817;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_597;
wire n_415;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_1128;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_440;
wire n_268;
wire n_858;
wire n_385;
wire n_729;
wire n_342;
wire n_430;
wire n_414;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_805;
wire n_820;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_1016;
wire n_482;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1119;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_1136;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_513;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_737;
wire n_606;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_890;
wire n_921;
wire n_874;
wire n_912;
wire n_1058;
wire n_1105;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_503;
wire n_292;
wire n_807;
wire n_1000;
wire n_394;
wire n_984;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_298;
wire n_1035;
wire n_587;
wire n_760;
wire n_1038;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_220),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_137),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_211),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_90),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_77),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_52),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_25),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_94),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_112),
.Y(n_255)
);

BUFx8_ASAP7_75t_SL g256 ( 
.A(n_97),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_59),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_68),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_172),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_114),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_188),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_192),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_50),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_140),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_239),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_144),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_138),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_65),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_33),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_81),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_117),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_196),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_85),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_201),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_241),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_33),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_31),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_197),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_175),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_132),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_96),
.Y(n_286)
);

BUFx2_ASAP7_75t_SL g287 ( 
.A(n_128),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_45),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_208),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_213),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_202),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_150),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_229),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_2),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_153),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_34),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_122),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_88),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_131),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_178),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_101),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_43),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_215),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_100),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_20),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_118),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_154),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_133),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_104),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_98),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_189),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_183),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_210),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_63),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_34),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_219),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_199),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_82),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_170),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_24),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_110),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_65),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_186),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_48),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_145),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_84),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_224),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_55),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_226),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_20),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_44),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_237),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_222),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_111),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_181),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_198),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_205),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_134),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_194),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_120),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_142),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_179),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_160),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_92),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_212),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_232),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_9),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_195),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_234),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_109),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_116),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_193),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_216),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_227),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_207),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_91),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_76),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_127),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_135),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_203),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_146),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_99),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_99),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_149),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_90),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_171),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_113),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_200),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_165),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_228),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_173),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_66),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_209),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_89),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_57),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_218),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_123),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_107),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_206),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_230),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_47),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_221),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_74),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_148),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_143),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_243),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_76),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_86),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_12),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_204),
.Y(n_392)
);

BUFx10_ASAP7_75t_L g393 ( 
.A(n_141),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_32),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_217),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_152),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_242),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_2),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_49),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_106),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_32),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_130),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_108),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_161),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_214),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_139),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_11),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_136),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_129),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_100),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_59),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_40),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_30),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_164),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_10),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_115),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_158),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_235),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_37),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_35),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_147),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_420),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_279),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_327),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_364),
.B(n_0),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_260),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_394),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_261),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_271),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_263),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_372),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_295),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_256),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_274),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_322),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_256),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_254),
.B(n_0),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_303),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_254),
.B(n_1),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_334),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_406),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_339),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_339),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_372),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_315),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_264),
.B(n_1),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_417),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_266),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_323),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_316),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_285),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_248),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_333),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_416),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_269),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_333),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_269),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_340),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_385),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_340),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_385),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_257),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_360),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_257),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_252),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_259),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_360),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_362),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_362),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_370),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_370),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_266),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_375),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_257),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_273),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_277),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_326),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_330),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_375),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_378),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_378),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_395),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_395),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_368),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_294),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_294),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_368),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_431),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_444),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_444),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_426),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_445),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_429),
.Y(n_496)
);

CKINVDCx14_ASAP7_75t_R g497 ( 
.A(n_486),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_434),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_432),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_437),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_454),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_445),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_442),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_489),
.B(n_267),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_443),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_450),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_433),
.B(n_318),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_474),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_446),
.B(n_354),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_446),
.B(n_267),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_449),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_464),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_466),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_457),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_474),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_487),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_455),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_439),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_487),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_459),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_460),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_488),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_430),
.B(n_267),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g526 ( 
.A1(n_488),
.A2(n_325),
.B(n_308),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_470),
.B(n_249),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_423),
.B(n_390),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_486),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_470),
.B(n_250),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_465),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_467),
.B(n_400),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_458),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_461),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_463),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_468),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_477),
.B(n_308),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_469),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_478),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_456),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_479),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_471),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_472),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_475),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_422),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_480),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_424),
.B(n_393),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_471),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_427),
.B(n_411),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_481),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_473),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_436),
.B(n_413),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_473),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_448),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_425),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_485),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_484),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_462),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_R g560 ( 
.A(n_435),
.B(n_245),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_438),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_482),
.B(n_419),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_483),
.B(n_325),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_R g564 ( 
.A(n_440),
.B(n_247),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_447),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_451),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_431),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_476),
.B(n_287),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_431),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_444),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_450),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_426),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_444),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_426),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_431),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_450),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_431),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_426),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_426),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_444),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_454),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_426),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_431),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_426),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_R g585 ( 
.A(n_453),
.B(n_258),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_444),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_444),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_450),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_446),
.B(n_265),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_431),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_454),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_431),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_431),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_454),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_431),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_431),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_444),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_486),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_431),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_431),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_426),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_490),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_526),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_518),
.B(n_281),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_591),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_490),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_492),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_555),
.B(n_255),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_513),
.B(n_253),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_515),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_589),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_495),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_568),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_594),
.B(n_501),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_512),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_517),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_516),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_529),
.B(n_550),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_519),
.A2(n_399),
.B1(n_251),
.B2(n_270),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_541),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_568),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_580),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_524),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_510),
.B(n_345),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_581),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_507),
.B(n_268),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_570),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_568),
.B(n_399),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_573),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_520),
.B(n_537),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_524),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_524),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_548),
.B(n_246),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_571),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_525),
.B(n_275),
.Y(n_636)
);

NOR2x1p5_ASAP7_75t_L g637 ( 
.A(n_561),
.B(n_494),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_586),
.Y(n_638)
);

INVx6_ASAP7_75t_L g639 ( 
.A(n_502),
.Y(n_639)
);

INVx6_ASAP7_75t_L g640 ( 
.A(n_502),
.Y(n_640)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_542),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_571),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_587),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_576),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_597),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_546),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_553),
.B(n_276),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_547),
.B(n_563),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_535),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_564),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_540),
.B(n_278),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_588),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_588),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_508),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_538),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_504),
.B(n_289),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_521),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_533),
.B(n_280),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_491),
.A2(n_399),
.B1(n_262),
.B2(n_284),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_562),
.B(n_288),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_530),
.B(n_399),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_498),
.B(n_283),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_496),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_557),
.B(n_300),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_536),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_558),
.A2(n_299),
.B1(n_305),
.B2(n_297),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_536),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_567),
.B(n_309),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_565),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_569),
.B(n_329),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_598),
.B(n_272),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_575),
.B(n_577),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_583),
.A2(n_291),
.B1(n_292),
.B2(n_290),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_590),
.B(n_369),
.Y(n_674)
);

NAND3xp33_ASAP7_75t_L g675 ( 
.A(n_585),
.B(n_311),
.C(n_306),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_493),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_592),
.B(n_593),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_595),
.B(n_321),
.C(n_319),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_493),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_596),
.B(n_403),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_599),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_600),
.Y(n_682)
);

AND2x2_ASAP7_75t_SL g683 ( 
.A(n_562),
.B(n_298),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_506),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_534),
.B(n_296),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_499),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_514),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_500),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_497),
.B(n_302),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_560),
.B(n_328),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_528),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_522),
.B(n_304),
.Y(n_692)
);

XNOR2xp5_ASAP7_75t_L g693 ( 
.A(n_543),
.B(n_332),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_523),
.B(n_307),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_532),
.B(n_310),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_539),
.A2(n_349),
.B1(n_358),
.B2(n_346),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_544),
.B(n_312),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_545),
.B(n_282),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_551),
.B(n_503),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_505),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_511),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_572),
.A2(n_365),
.B1(n_367),
.B2(n_359),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_601),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_566),
.B(n_314),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_574),
.B(n_313),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_561),
.B(n_320),
.Y(n_706)
);

INVxp33_ASAP7_75t_L g707 ( 
.A(n_531),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_578),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_579),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_582),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_584),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_559),
.B(n_286),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_549),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_552),
.B(n_374),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_554),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_568),
.B(n_376),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_509),
.B(n_317),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_512),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_556),
.B(n_324),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_565),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_526),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_565),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_548),
.A2(n_377),
.B1(n_391),
.B2(n_383),
.Y(n_723)
);

OR2x6_ASAP7_75t_L g724 ( 
.A(n_512),
.B(n_336),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_518),
.B(n_398),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_512),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_526),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_526),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_591),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_518),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_490),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_526),
.Y(n_732)
);

INVx4_ASAP7_75t_SL g733 ( 
.A(n_568),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_556),
.B(n_331),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_518),
.B(n_401),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_490),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_591),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_730),
.B(n_407),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_605),
.B(n_410),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_729),
.B(n_335),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_737),
.Y(n_741)
);

CKINVDCx11_ASAP7_75t_R g742 ( 
.A(n_663),
.Y(n_742)
);

BUFx8_ASAP7_75t_L g743 ( 
.A(n_650),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_655),
.A2(n_338),
.B(n_341),
.C(n_337),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_625),
.B(n_412),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_616),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_649),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_613),
.B(n_343),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_613),
.B(n_344),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_648),
.B(n_415),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_665),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_657),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_620),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_614),
.B(n_604),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_631),
.B(n_356),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_618),
.B(n_347),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_733),
.B(n_342),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_657),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_654),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_641),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_688),
.B(n_621),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_611),
.B(n_348),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_683),
.A2(n_352),
.B1(n_353),
.B2(n_351),
.Y(n_763)
);

BUFx12f_ASAP7_75t_L g764 ( 
.A(n_663),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_716),
.B(n_350),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_716),
.B(n_355),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_681),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_682),
.A2(n_361),
.B1(n_363),
.B2(n_357),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_626),
.B(n_366),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_667),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_684),
.Y(n_771)
);

INVx5_ASAP7_75t_L g772 ( 
.A(n_629),
.Y(n_772)
);

BUFx8_ASAP7_75t_L g773 ( 
.A(n_699),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_629),
.A2(n_382),
.B1(n_384),
.B2(n_371),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_634),
.A2(n_388),
.B1(n_392),
.B2(n_386),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_677),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_725),
.B(n_3),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_634),
.A2(n_402),
.B1(n_404),
.B2(n_396),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_615),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_669),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_634),
.A2(n_409),
.B1(n_414),
.B2(n_405),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_735),
.B(n_4),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_607),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_672),
.B(n_421),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_607),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_661),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_603),
.B(n_397),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_733),
.B(n_418),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_612),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_612),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_622),
.B(n_380),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_636),
.B(n_381),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_721),
.B(n_397),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_717),
.B(n_387),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_718),
.Y(n_795)
);

BUFx6f_ASAP7_75t_SL g796 ( 
.A(n_711),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_727),
.B(n_728),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_726),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_732),
.A2(n_408),
.B(n_293),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_SL g800 ( 
.A(n_720),
.B(n_722),
.C(n_712),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_646),
.B(n_647),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_628),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_630),
.Y(n_803)
);

INVx5_ASAP7_75t_L g804 ( 
.A(n_610),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_630),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_668),
.B(n_5),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_670),
.B(n_5),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_638),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_674),
.B(n_6),
.Y(n_809)
);

AND2x4_ASAP7_75t_SL g810 ( 
.A(n_711),
.B(n_301),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_680),
.B(n_6),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_638),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_723),
.B(n_7),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_691),
.B(n_7),
.C(n_8),
.Y(n_814)
);

AOI221xp5_ASAP7_75t_L g815 ( 
.A1(n_660),
.A2(n_379),
.B1(n_14),
.B2(n_10),
.C(n_13),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_698),
.B(n_13),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_724),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_643),
.Y(n_818)
);

AND2x6_ASAP7_75t_SL g819 ( 
.A(n_714),
.B(n_15),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_645),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_679),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_645),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_678),
.A2(n_379),
.B1(n_18),
.B2(n_16),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_632),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_624),
.A2(n_379),
.B1(n_19),
.B2(n_17),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_698),
.B(n_18),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_676),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_679),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_609),
.B(n_21),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_664),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_666),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_831)
);

BUFx12f_ASAP7_75t_L g832 ( 
.A(n_637),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_686),
.B(n_26),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_619),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_675),
.B(n_27),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_673),
.B(n_28),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_679),
.B(n_29),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_L g838 ( 
.A1(n_671),
.A2(n_703),
.B1(n_704),
.B2(n_700),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_651),
.B(n_30),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_696),
.A2(n_36),
.B(n_31),
.C(n_35),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_656),
.B(n_36),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_719),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_659),
.B(n_39),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_690),
.B(n_40),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_658),
.B(n_41),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_701),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_734),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_744),
.A2(n_830),
.B(n_840),
.C(n_836),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_741),
.A2(n_714),
.B1(n_708),
.B2(n_709),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_772),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_797),
.A2(n_608),
.B(n_662),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_754),
.B(n_713),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_776),
.A2(n_708),
.B1(n_710),
.B2(n_709),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_746),
.Y(n_854)
);

BUFx4f_ASAP7_75t_L g855 ( 
.A(n_764),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_767),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_752),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_799),
.A2(n_606),
.B(n_602),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_838),
.B(n_715),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_758),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_772),
.A2(n_671),
.B1(n_704),
.B2(n_687),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_761),
.B(n_706),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_817),
.B(n_707),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_787),
.A2(n_736),
.B(n_617),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_800),
.B(n_689),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_783),
.Y(n_866)
);

O2A1O1Ixp5_ASAP7_75t_L g867 ( 
.A1(n_841),
.A2(n_633),
.B(n_635),
.C(n_623),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_801),
.B(n_706),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_L g869 ( 
.A(n_815),
.B(n_702),
.C(n_697),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_836),
.A2(n_692),
.B(n_705),
.C(n_695),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_739),
.B(n_693),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_777),
.B(n_782),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_799),
.A2(n_644),
.B(n_642),
.Y(n_873)
);

AOI21xp33_ASAP7_75t_L g874 ( 
.A1(n_738),
.A2(n_694),
.B(n_685),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_793),
.A2(n_731),
.B(n_653),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_753),
.B(n_627),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_760),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_759),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_755),
.B(n_639),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_750),
.B(n_763),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_784),
.B(n_816),
.Y(n_881)
);

BUFx12f_ASAP7_75t_L g882 ( 
.A(n_742),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_784),
.B(n_640),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_803),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_745),
.B(n_640),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_786),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_826),
.B(n_813),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_805),
.Y(n_888)
);

BUFx12f_ASAP7_75t_L g889 ( 
.A(n_743),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_812),
.Y(n_890)
);

NOR3xp33_ASAP7_75t_L g891 ( 
.A(n_814),
.B(n_46),
.C(n_48),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_769),
.A2(n_652),
.B(n_103),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_829),
.B(n_49),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_785),
.A2(n_790),
.B1(n_802),
.B2(n_789),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_818),
.A2(n_51),
.B(n_52),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_820),
.A2(n_105),
.B(n_102),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_822),
.B(n_53),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_796),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_827),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_808),
.B(n_54),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_765),
.B(n_54),
.Y(n_901)
);

NOR2x1p5_ASAP7_75t_L g902 ( 
.A(n_780),
.B(n_832),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_768),
.B(n_55),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_844),
.A2(n_60),
.B1(n_56),
.B2(n_58),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_845),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_768),
.B(n_56),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_766),
.B(n_58),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_756),
.B(n_60),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_845),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_796),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_910)
);

CKINVDCx10_ASAP7_75t_R g911 ( 
.A(n_773),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_795),
.B(n_61),
.Y(n_912)
);

NAND2x1p5_ASAP7_75t_L g913 ( 
.A(n_804),
.B(n_62),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_775),
.A2(n_67),
.B1(n_64),
.B2(n_66),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_773),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_806),
.A2(n_121),
.B(n_119),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_837),
.A2(n_125),
.B(n_124),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_L g918 ( 
.A(n_804),
.B(n_126),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_778),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_762),
.B(n_71),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_771),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_781),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_807),
.B(n_72),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_809),
.B(n_73),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_811),
.B(n_75),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_850),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_877),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_905),
.B(n_747),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_868),
.B(n_748),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_859),
.A2(n_833),
.B1(n_839),
.B2(n_757),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_889),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_881),
.B(n_774),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_852),
.B(n_798),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_861),
.B(n_804),
.Y(n_934)
);

OAI21x1_ASAP7_75t_SL g935 ( 
.A1(n_895),
.A2(n_846),
.B(n_831),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_862),
.B(n_810),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_855),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_850),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_880),
.B(n_792),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_848),
.A2(n_825),
.B(n_835),
.C(n_843),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_917),
.A2(n_828),
.B(n_821),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_913),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_R g943 ( 
.A(n_911),
.B(n_743),
.Y(n_943)
);

NAND2x1p5_ASAP7_75t_L g944 ( 
.A(n_855),
.B(n_779),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_913),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_864),
.A2(n_770),
.B(n_824),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_909),
.B(n_794),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_882),
.B(n_788),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_870),
.A2(n_842),
.B(n_847),
.C(n_823),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_854),
.Y(n_950)
);

NOR2x1_ASAP7_75t_SL g951 ( 
.A(n_894),
.B(n_751),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_856),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_866),
.B(n_834),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_853),
.B(n_749),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_899),
.Y(n_955)
);

AO21x1_ASAP7_75t_L g956 ( 
.A1(n_895),
.A2(n_740),
.B(n_791),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_884),
.B(n_819),
.Y(n_957)
);

BUFx12f_ASAP7_75t_L g958 ( 
.A(n_898),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_888),
.B(n_75),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_875),
.A2(n_916),
.B(n_892),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_873),
.A2(n_867),
.B(n_858),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_890),
.Y(n_962)
);

OAI22x1_ASAP7_75t_L g963 ( 
.A1(n_910),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_857),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_851),
.A2(n_78),
.B(n_79),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_865),
.B(n_860),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_878),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_921),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_886),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_869),
.A2(n_80),
.B(n_81),
.Y(n_970)
);

OA22x2_ASAP7_75t_L g971 ( 
.A1(n_849),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_932),
.B(n_903),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_950),
.B(n_906),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_970),
.A2(n_965),
.B(n_920),
.C(n_908),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_927),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_964),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_952),
.B(n_887),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_942),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_958),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_970),
.A2(n_901),
.B(n_907),
.C(n_891),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_931),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_955),
.Y(n_982)
);

CKINVDCx11_ASAP7_75t_R g983 ( 
.A(n_948),
.Y(n_983)
);

AOI21xp33_ASAP7_75t_SL g984 ( 
.A1(n_937),
.A2(n_915),
.B(n_871),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_930),
.A2(n_872),
.B1(n_893),
.B2(n_883),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_940),
.A2(n_924),
.B(n_923),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_954),
.B(n_863),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_SL g988 ( 
.A(n_944),
.B(n_898),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_933),
.B(n_904),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_945),
.Y(n_990)
);

BUFx4f_ASAP7_75t_SL g991 ( 
.A(n_936),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_943),
.Y(n_992)
);

BUFx5_ASAP7_75t_L g993 ( 
.A(n_968),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_936),
.B(n_902),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_962),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_949),
.A2(n_939),
.B(n_947),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_947),
.B(n_897),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_969),
.B(n_900),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_929),
.B(n_885),
.Y(n_999)
);

NOR3xp33_ASAP7_75t_L g1000 ( 
.A(n_957),
.B(n_874),
.C(n_914),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_926),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_959),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_967),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_926),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_972),
.B(n_977),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_982),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_991),
.A2(n_971),
.B1(n_965),
.B2(n_934),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_995),
.B(n_967),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_980),
.A2(n_974),
.B(n_996),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_1001),
.B(n_966),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_975),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_1000),
.A2(n_935),
.B1(n_963),
.B2(n_956),
.Y(n_1012)
);

AO21x1_ASAP7_75t_SL g1013 ( 
.A1(n_1003),
.A2(n_896),
.B(n_928),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_993),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_986),
.A2(n_941),
.B(n_946),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_1001),
.A2(n_960),
.B(n_961),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_981),
.B(n_948),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_SL g1018 ( 
.A1(n_991),
.A2(n_966),
.B1(n_951),
.B2(n_938),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_976),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_987),
.B(n_953),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_993),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_993),
.Y(n_1022)
);

AO21x1_ASAP7_75t_SL g1023 ( 
.A1(n_1003),
.A2(n_990),
.B(n_978),
.Y(n_1023)
);

CKINVDCx6p67_ASAP7_75t_R g1024 ( 
.A(n_979),
.Y(n_1024)
);

BUFx8_ASAP7_75t_SL g1025 ( 
.A(n_994),
.Y(n_1025)
);

INVx6_ASAP7_75t_L g1026 ( 
.A(n_979),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_993),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_973),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_1000),
.A2(n_919),
.B1(n_922),
.B2(n_912),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1028),
.B(n_987),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1014),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_1021),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_1014),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_1022),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1022),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1006),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1011),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_1026),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1021),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1027),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_1027),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_1005),
.B(n_998),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_1008),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1019),
.Y(n_1044)
);

BUFx4f_ASAP7_75t_SL g1045 ( 
.A(n_1024),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1023),
.B(n_993),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1008),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_1023),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1016),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1015),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1009),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1036),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1031),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_1048),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_1043),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1036),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_1045),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_1049),
.A2(n_1007),
.A3(n_1020),
.B(n_985),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_1032),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1037),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_SL g1061 ( 
.A1(n_1046),
.A2(n_1026),
.B1(n_993),
.B2(n_990),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1037),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1051),
.B(n_1012),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_1032),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1047),
.B(n_1013),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1031),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_1041),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1051),
.B(n_1010),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1031),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1047),
.B(n_1013),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1055),
.B(n_1044),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_L g1072 ( 
.A(n_1063),
.B(n_1064),
.C(n_1059),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1058),
.B(n_1042),
.Y(n_1073)
);

OAI211xp5_ASAP7_75t_L g1074 ( 
.A1(n_1054),
.A2(n_983),
.B(n_1057),
.C(n_1061),
.Y(n_1074)
);

OAI221xp5_ASAP7_75t_SL g1075 ( 
.A1(n_1054),
.A2(n_1024),
.B1(n_1030),
.B2(n_1042),
.C(n_994),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_1057),
.B(n_1046),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1065),
.B(n_1039),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1056),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1070),
.A2(n_989),
.B1(n_1025),
.B2(n_1017),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_L g1080 ( 
.A(n_1067),
.B(n_1040),
.C(n_1039),
.Y(n_1080)
);

NAND4xp25_ASAP7_75t_L g1081 ( 
.A(n_1068),
.B(n_999),
.C(n_1029),
.D(n_988),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1058),
.B(n_1040),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1073),
.B(n_1058),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1078),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1071),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_1080),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1077),
.B(n_1058),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1072),
.B(n_1058),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_1076),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1082),
.B(n_1056),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1074),
.B(n_1052),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1074),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1075),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1079),
.B(n_1053),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1081),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1071),
.Y(n_1096)
);

AOI33xp33_ASAP7_75t_L g1097 ( 
.A1(n_1093),
.A2(n_992),
.A3(n_1062),
.B1(n_1060),
.B2(n_1002),
.B3(n_1018),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1092),
.B(n_1038),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1084),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1085),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1089),
.B(n_1066),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1084),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1096),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_1098),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1099),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1100),
.Y(n_1106)
);

AOI21xp33_ASAP7_75t_SL g1107 ( 
.A1(n_1103),
.A2(n_1095),
.B(n_1086),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_1104),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1106),
.B(n_1095),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_1104),
.B(n_1083),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1108),
.B(n_1107),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1109),
.B(n_1088),
.Y(n_1112)
);

OAI322xp33_ASAP7_75t_L g1113 ( 
.A1(n_1110),
.A2(n_1091),
.A3(n_1088),
.B1(n_1105),
.B2(n_1090),
.C1(n_1102),
.C2(n_1099),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1111),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1112),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1113),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_1111),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_L g1118 ( 
.A(n_1117),
.B(n_984),
.C(n_1097),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1116),
.A2(n_1101),
.B1(n_979),
.B2(n_1102),
.Y(n_1119)
);

NAND4xp25_ASAP7_75t_L g1120 ( 
.A(n_1114),
.B(n_1097),
.C(n_1025),
.D(n_1094),
.Y(n_1120)
);

AOI211xp5_ASAP7_75t_SL g1121 ( 
.A1(n_1115),
.A2(n_948),
.B(n_994),
.C(n_1026),
.Y(n_1121)
);

NAND4xp25_ASAP7_75t_L g1122 ( 
.A(n_1114),
.B(n_1094),
.C(n_997),
.D(n_1087),
.Y(n_1122)
);

NOR3x1_ASAP7_75t_L g1123 ( 
.A(n_1120),
.B(n_1122),
.C(n_1121),
.Y(n_1123)
);

NOR2x1_ASAP7_75t_L g1124 ( 
.A(n_1118),
.B(n_925),
.Y(n_1124)
);

NOR4xp25_ASAP7_75t_L g1125 ( 
.A(n_1119),
.B(n_879),
.C(n_876),
.D(n_918),
.Y(n_1125)
);

NOR3x1_ASAP7_75t_L g1126 ( 
.A(n_1119),
.B(n_1004),
.C(n_87),
.Y(n_1126)
);

AND4x1_ASAP7_75t_L g1127 ( 
.A(n_1123),
.B(n_1126),
.C(n_1124),
.D(n_1125),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1127),
.B(n_93),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_SL g1129 ( 
.A(n_1128),
.B(n_94),
.C(n_95),
.Y(n_1129)
);

AND3x1_ASAP7_75t_L g1130 ( 
.A(n_1129),
.B(n_1033),
.C(n_1069),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1130),
.A2(n_1050),
.B1(n_1034),
.B2(n_1035),
.Y(n_1131)
);

OAI322xp33_ASAP7_75t_L g1132 ( 
.A1(n_1131),
.A2(n_1050),
.A3(n_151),
.B1(n_155),
.B2(n_156),
.C1(n_157),
.C2(n_159),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1132),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_1133),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1134),
.Y(n_1135)
);

OAI331xp33_ASAP7_75t_L g1136 ( 
.A1(n_1135),
.A2(n_162),
.A3(n_163),
.B1(n_166),
.B2(n_167),
.B3(n_168),
.C1(n_169),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1136),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_1137)
);

OAI221xp5_ASAP7_75t_R g1138 ( 
.A1(n_1137),
.A2(n_180),
.B1(n_182),
.B2(n_184),
.C(n_185),
.Y(n_1138)
);

AOI211xp5_ASAP7_75t_L g1139 ( 
.A1(n_1138),
.A2(n_187),
.B(n_190),
.C(n_191),
.Y(n_1139)
);


endmodule