module fake_jpeg_1643_n_265 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_46),
.B(n_58),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_48),
.A2(n_57),
.B(n_25),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_20),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_85)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_23),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_62),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_20),
.C(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_6),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_61),
.Y(n_91)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_7),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_11),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_67),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_32),
.B(n_11),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_8),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_73),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_8),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_10),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_80),
.Y(n_114)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

CKINVDCx6p67_ASAP7_75t_R g113 ( 
.A(n_78),
.Y(n_113)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_10),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_55),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_92),
.C(n_102),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_45),
.B1(n_67),
.B2(n_54),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_87),
.A2(n_120),
.B1(n_86),
.B2(n_110),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_41),
.B1(n_26),
.B2(n_34),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_90),
.A2(n_93),
.B1(n_122),
.B2(n_97),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_34),
.B(n_29),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_99),
.A2(n_96),
.B(n_121),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_29),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_104),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_31),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_41),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_108),
.B(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_78),
.B(n_27),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_44),
.B(n_47),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_49),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_125),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_64),
.A2(n_35),
.B1(n_51),
.B2(n_60),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_124),
.B(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_56),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_118),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_130),
.Y(n_172)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_136),
.Y(n_176)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_118),
.B(n_84),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_141),
.B(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_101),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_89),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_89),
.B(n_101),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_153),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_96),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_86),
.B(n_97),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_161),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_133),
.Y(n_169)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_93),
.B(n_122),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_88),
.C(n_92),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_136),
.C(n_162),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_169),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_132),
.B(n_163),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_171),
.B(n_173),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_178),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_130),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_158),
.A2(n_159),
.B1(n_146),
.B2(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_181),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_154),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_145),
.C(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_136),
.B(n_149),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_139),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_150),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_208),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_126),
.B(n_138),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_198),
.C(n_200),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_128),
.B(n_137),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_180),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_164),
.B(n_131),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_204),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_176),
.A2(n_134),
.B(n_129),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_129),
.B1(n_175),
.B2(n_177),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_207),
.B1(n_171),
.B2(n_167),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_187),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_183),
.C(n_188),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_179),
.B1(n_169),
.B2(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_173),
.B1(n_170),
.B2(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_191),
.B1(n_193),
.B2(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_206),
.C(n_200),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_226),
.C(n_228),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_209),
.C(n_207),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_195),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_195),
.C(n_197),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_221),
.C(n_215),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_217),
.A2(n_190),
.B1(n_203),
.B2(n_184),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_213),
.Y(n_240)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_235),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_213),
.A2(n_204),
.B(n_192),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_204),
.B(n_215),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_194),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_241),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_230),
.C(n_232),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_230),
.A2(n_210),
.B1(n_212),
.B2(n_222),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_244),
.B(n_236),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_234),
.B(n_232),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_212),
.B(n_210),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_246),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_229),
.B(n_228),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_237),
.B1(n_219),
.B2(n_216),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_250),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_233),
.B(n_226),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_255),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_SL g253 ( 
.A1(n_249),
.A2(n_243),
.B(n_241),
.C(n_239),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_225),
.C(n_224),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_239),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_256),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_251),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_224),
.B1(n_208),
.B2(n_253),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_258),
.A2(n_253),
.B(n_259),
.Y(n_261)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_262),
.B(n_199),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_263),
.B(n_264),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_185),
.C(n_186),
.Y(n_264)
);


endmodule