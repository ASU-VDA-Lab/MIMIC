module fake_netlist_1_4294_n_536 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_536);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_536;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_14), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_24), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_45), .Y(n_82) );
INVxp33_ASAP7_75t_SL g83 ( .A(n_33), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_0), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_22), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_23), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_26), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_65), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_0), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_4), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_54), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_66), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_75), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_9), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_49), .Y(n_95) );
INVxp33_ASAP7_75t_L g96 ( .A(n_42), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_37), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_7), .Y(n_98) );
INVxp33_ASAP7_75t_L g99 ( .A(n_70), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_59), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_21), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_16), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_36), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_25), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_10), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_7), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_40), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_60), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_79), .Y(n_109) );
BUFx6f_ASAP7_75t_SL g110 ( .A(n_39), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_38), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_11), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_63), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_47), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_17), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_58), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_15), .Y(n_117) );
AND2x4_ASAP7_75t_L g118 ( .A(n_80), .B(n_1), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_104), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_85), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_104), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_85), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_87), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_106), .Y(n_125) );
OAI21x1_ASAP7_75t_L g126 ( .A1(n_86), .A2(n_35), .B(n_77), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_106), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
CKINVDCx9p33_ASAP7_75t_R g129 ( .A(n_86), .Y(n_129) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_114), .A2(n_34), .B(n_76), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_104), .B(n_2), .Y(n_133) );
INVx4_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_93), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_104), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_104), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_112), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_95), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_91), .B(n_3), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_134), .B(n_82), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_134), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_125), .Y(n_143) );
INVxp67_ASAP7_75t_SL g144 ( .A(n_125), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_134), .B(n_111), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_134), .B(n_118), .Y(n_146) );
INVx4_ASAP7_75t_L g147 ( .A(n_118), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_120), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_120), .Y(n_151) );
CKINVDCx8_ASAP7_75t_R g152 ( .A(n_118), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_138), .B(n_116), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_138), .Y(n_157) );
INVx5_ASAP7_75t_L g158 ( .A(n_119), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_123), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_123), .B(n_92), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_119), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_124), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_119), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_119), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_141), .B(n_140), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_141), .B(n_128), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_146), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
BUFx12f_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_161), .B(n_128), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
NOR2x1_ASAP7_75t_L g178 ( .A(n_145), .B(n_140), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_146), .Y(n_180) );
OR2x6_ASAP7_75t_SL g181 ( .A(n_154), .B(n_112), .Y(n_181) );
NAND3xp33_ASAP7_75t_SL g182 ( .A(n_152), .B(n_127), .C(n_100), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_152), .B(n_100), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_156), .B(n_131), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_156), .B(n_131), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_153), .A2(n_127), .B1(n_139), .B2(n_135), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_144), .B(n_132), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_147), .B(n_83), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_147), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_159), .A2(n_132), .B(n_135), .C(n_139), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_150), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_142), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_159), .B(n_96), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_160), .B(n_99), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_153), .B(n_95), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_160), .B(n_101), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_147), .A2(n_80), .B1(n_94), .B2(n_115), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_170), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_177), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_174), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_177), .Y(n_204) );
BUFx4_ASAP7_75t_SL g205 ( .A(n_176), .Y(n_205) );
CKINVDCx8_ASAP7_75t_R g206 ( .A(n_176), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_168), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_170), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_177), .Y(n_209) );
AO32x1_ASAP7_75t_L g210 ( .A1(n_172), .A2(n_137), .A3(n_136), .B1(n_121), .B2(n_107), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_177), .Y(n_211) );
INVx2_ASAP7_75t_SL g212 ( .A(n_170), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_168), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_173), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_173), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_172), .B(n_147), .Y(n_216) );
CKINVDCx8_ASAP7_75t_R g217 ( .A(n_198), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_171), .B(n_163), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_175), .B(n_163), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_167), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_182), .A2(n_155), .B1(n_164), .B2(n_133), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_179), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_198), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_179), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_193), .Y(n_225) );
BUFx12f_ASAP7_75t_L g226 ( .A(n_174), .Y(n_226) );
OR2x2_ASAP7_75t_L g227 ( .A(n_187), .B(n_164), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_177), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_198), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_180), .Y(n_230) );
INVx1_ASAP7_75t_SL g231 ( .A(n_174), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_180), .B(n_155), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_192), .Y(n_234) );
OR2x6_ASAP7_75t_L g235 ( .A(n_223), .B(n_169), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_207), .Y(n_236) );
CKINVDCx6p67_ASAP7_75t_R g237 ( .A(n_226), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_208), .A2(n_178), .B1(n_198), .B2(n_186), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_208), .A2(n_178), .B1(n_198), .B2(n_186), .Y(n_239) );
INVxp67_ASAP7_75t_SL g240 ( .A(n_223), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_207), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_201), .A2(n_198), .B1(n_187), .B2(n_155), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_227), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_227), .A2(n_194), .B1(n_195), .B2(n_184), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_213), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_213), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_201), .A2(n_198), .B1(n_155), .B2(n_183), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_217), .A2(n_185), .B1(n_181), .B2(n_200), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_219), .B(n_181), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_202), .A2(n_188), .B1(n_189), .B2(n_196), .Y(n_250) );
OAI22xp33_ASAP7_75t_L g251 ( .A1(n_206), .A2(n_199), .B1(n_197), .B2(n_196), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_206), .B(n_231), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_220), .Y(n_253) );
BUFx2_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_214), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_202), .B(n_189), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_226), .Y(n_257) );
BUFx2_ASAP7_75t_R g258 ( .A(n_203), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_229), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_217), .A2(n_196), .B1(n_167), .B2(n_191), .Y(n_260) );
AOI21x1_ASAP7_75t_L g261 ( .A1(n_214), .A2(n_130), .B(n_126), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_215), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_244), .A2(n_190), .B1(n_218), .B2(n_221), .C(n_215), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_253), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_249), .A2(n_202), .B1(n_212), .B2(n_232), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_248), .A2(n_202), .B1(n_212), .B2(n_232), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_251), .A2(n_224), .B1(n_222), .B2(n_225), .Y(n_267) );
OAI22xp33_ASAP7_75t_L g268 ( .A1(n_237), .A2(n_205), .B1(n_225), .B2(n_224), .Y(n_268) );
INVx4_ASAP7_75t_SL g269 ( .A(n_257), .Y(n_269) );
OAI22xp5_ASAP7_75t_SL g270 ( .A1(n_252), .A2(n_222), .B1(n_84), .B2(n_90), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_238), .A2(n_220), .B1(n_234), .B2(n_228), .Y(n_271) );
OAI22xp5_ASAP7_75t_SL g272 ( .A1(n_243), .A2(n_94), .B1(n_84), .B2(n_89), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_236), .B(n_204), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_236), .B(n_167), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_239), .A2(n_230), .B1(n_204), .B2(n_228), .Y(n_275) );
OAI211xp5_ASAP7_75t_SL g276 ( .A1(n_250), .A2(n_117), .B(n_105), .C(n_98), .Y(n_276) );
NAND3xp33_ASAP7_75t_L g277 ( .A(n_260), .B(n_211), .C(n_209), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_253), .Y(n_278) );
NOR2xp67_ASAP7_75t_SL g279 ( .A(n_259), .B(n_234), .Y(n_279) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_237), .A2(n_230), .B1(n_228), .B2(n_209), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_241), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g282 ( .A1(n_242), .A2(n_233), .B(n_216), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_241), .B(n_191), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_259), .Y(n_284) );
OAI22xp5_ASAP7_75t_SL g285 ( .A1(n_257), .A2(n_115), .B1(n_89), .B2(n_90), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_277), .A2(n_261), .B(n_130), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_264), .Y(n_287) );
AOI222xp33_ASAP7_75t_L g288 ( .A1(n_285), .A2(n_102), .B1(n_262), .B2(n_255), .C1(n_246), .C2(n_245), .Y(n_288) );
NOR3xp33_ASAP7_75t_L g289 ( .A(n_268), .B(n_108), .C(n_113), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_281), .Y(n_290) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_267), .A2(n_247), .B(n_245), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_270), .A2(n_235), .B1(n_254), .B2(n_246), .Y(n_292) );
AOI22xp5_ASAP7_75t_SL g293 ( .A1(n_284), .A2(n_254), .B1(n_240), .B2(n_259), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_281), .B(n_255), .Y(n_294) );
AOI322xp5_ASAP7_75t_L g295 ( .A1(n_266), .A2(n_262), .A3(n_108), .B1(n_113), .B2(n_107), .C1(n_109), .C2(n_103), .Y(n_295) );
OAI22xp33_ASAP7_75t_L g296 ( .A1(n_284), .A2(n_235), .B1(n_230), .B2(n_228), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_270), .A2(n_235), .B1(n_256), .B2(n_209), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_274), .B(n_235), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_272), .B(n_258), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_276), .A2(n_209), .B1(n_228), .B2(n_211), .Y(n_300) );
OAI221xp5_ASAP7_75t_L g301 ( .A1(n_285), .A2(n_204), .B1(n_230), .B2(n_81), .C(n_97), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_264), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_278), .B(n_204), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_278), .B(n_209), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_274), .B(n_209), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_283), .Y(n_306) );
NAND3xp33_ASAP7_75t_L g307 ( .A(n_263), .B(n_119), .C(n_121), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_283), .Y(n_308) );
INVx4_ASAP7_75t_L g309 ( .A(n_305), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_290), .B(n_273), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_290), .B(n_114), .Y(n_311) );
AOI22xp33_ASAP7_75t_SL g312 ( .A1(n_293), .A2(n_272), .B1(n_277), .B2(n_271), .Y(n_312) );
OAI31xp33_ASAP7_75t_L g313 ( .A1(n_301), .A2(n_265), .A3(n_280), .B(n_269), .Y(n_313) );
OR2x6_ASAP7_75t_L g314 ( .A(n_308), .B(n_279), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_302), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_305), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_302), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_293), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_302), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_287), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_289), .A2(n_110), .B1(n_282), .B2(n_275), .C(n_121), .Y(n_321) );
NOR2xp67_ASAP7_75t_L g322 ( .A(n_307), .B(n_261), .Y(n_322) );
AOI22xp33_ASAP7_75t_SL g323 ( .A1(n_299), .A2(n_269), .B1(n_110), .B2(n_279), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_287), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_308), .B(n_126), .Y(n_325) );
INVxp67_ASAP7_75t_SL g326 ( .A(n_308), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_306), .Y(n_327) );
OAI211xp5_ASAP7_75t_SL g328 ( .A1(n_288), .A2(n_137), .B(n_136), .C(n_269), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_306), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_294), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_304), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_295), .B(n_269), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_303), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_286), .Y(n_336) );
NOR3xp33_ASAP7_75t_L g337 ( .A(n_307), .B(n_136), .C(n_137), .Y(n_337) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_295), .B(n_119), .C(n_211), .Y(n_338) );
NAND2x1p5_ASAP7_75t_L g339 ( .A(n_309), .B(n_304), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_330), .B(n_298), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_327), .B(n_298), .Y(n_341) );
OAI211xp5_ASAP7_75t_SL g342 ( .A1(n_333), .A2(n_292), .B(n_297), .C(n_291), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_327), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_315), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_329), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_329), .B(n_304), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_315), .B(n_286), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_315), .B(n_126), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_338), .A2(n_300), .B1(n_296), .B2(n_228), .Y(n_349) );
NOR2xp33_ASAP7_75t_SL g350 ( .A(n_318), .B(n_211), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_330), .B(n_4), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_319), .B(n_130), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_331), .B(n_5), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_338), .B(n_119), .C(n_165), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_319), .B(n_5), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_322), .A2(n_210), .B(n_211), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_316), .B(n_309), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_331), .B(n_6), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_334), .B(n_6), .Y(n_359) );
INVxp67_ASAP7_75t_SL g360 ( .A(n_319), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_320), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_335), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_332), .B(n_8), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_323), .B(n_8), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_320), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_332), .B(n_9), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_312), .A2(n_211), .B1(n_191), .B2(n_197), .Y(n_367) );
INVx3_ASAP7_75t_SL g368 ( .A(n_314), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_324), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_309), .B(n_10), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_324), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_326), .B(n_11), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_317), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_309), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_335), .B(n_12), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_335), .B(n_12), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_334), .B(n_13), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_336), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_310), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_310), .B(n_13), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_314), .B(n_14), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_314), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_354), .A2(n_322), .B(n_321), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_380), .B(n_311), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_375), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_364), .B(n_328), .C(n_311), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_342), .A2(n_314), .B1(n_337), .B2(n_325), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_343), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_343), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_345), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g392 ( .A1(n_382), .A2(n_313), .B(n_314), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_357), .B(n_15), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_341), .B(n_16), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_357), .B(n_17), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_345), .Y(n_396) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_370), .B(n_129), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_346), .B(n_18), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_370), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_381), .B(n_18), .Y(n_400) );
CKINVDCx16_ASAP7_75t_R g401 ( .A(n_381), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_340), .B(n_19), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_354), .A2(n_210), .B(n_197), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_361), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_350), .B(n_165), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_365), .B(n_19), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_365), .B(n_20), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_369), .B(n_27), .Y(n_408) );
NAND2x1_ASAP7_75t_SL g409 ( .A(n_368), .B(n_210), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_360), .B(n_28), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_378), .B(n_29), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_376), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_350), .B(n_162), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_371), .B(n_30), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_346), .B(n_31), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_362), .B(n_32), .Y(n_416) );
XNOR2x2_ASAP7_75t_L g417 ( .A(n_382), .B(n_129), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_362), .B(n_41), .Y(n_418) );
NOR2x1_ASAP7_75t_L g419 ( .A(n_376), .B(n_210), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_344), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_378), .B(n_43), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_374), .B(n_44), .Y(n_422) );
INVxp67_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
NAND3xp33_ASAP7_75t_L g424 ( .A(n_367), .B(n_165), .C(n_162), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_374), .B(n_46), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_379), .B(n_48), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_373), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_401), .B(n_351), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_384), .B(n_368), .Y(n_429) );
AOI32xp33_ASAP7_75t_L g430 ( .A1(n_400), .A2(n_377), .A3(n_373), .B1(n_349), .B2(n_383), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_399), .B(n_355), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_427), .B(n_355), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_386), .Y(n_433) );
AOI221xp5_ASAP7_75t_SL g434 ( .A1(n_423), .A2(n_383), .B1(n_358), .B2(n_359), .C(n_353), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_389), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_387), .A2(n_368), .B1(n_363), .B2(n_366), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_390), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_393), .B(n_366), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_391), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_396), .Y(n_440) );
AND4x1_ASAP7_75t_L g441 ( .A(n_417), .B(n_363), .C(n_356), .D(n_339), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_412), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_404), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_395), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_420), .Y(n_445) );
XOR2x2_ASAP7_75t_L g446 ( .A(n_397), .B(n_339), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_397), .B(n_349), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_385), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_406), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_406), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_398), .Y(n_451) );
NOR2xp67_ASAP7_75t_SL g452 ( .A(n_418), .B(n_352), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g453 ( .A(n_394), .B(n_352), .C(n_348), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_402), .B(n_372), .Y(n_454) );
AO22x1_ASAP7_75t_L g455 ( .A1(n_416), .A2(n_347), .B1(n_348), .B2(n_210), .Y(n_455) );
NOR2x1_ASAP7_75t_L g456 ( .A(n_424), .B(n_50), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_407), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_405), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_415), .B(n_51), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_392), .B(n_52), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_392), .B(n_416), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_407), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_411), .B(n_53), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_388), .A2(n_165), .B1(n_162), .B2(n_192), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_421), .B(n_55), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_410), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_408), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_408), .Y(n_468) );
AO22x2_ASAP7_75t_L g469 ( .A1(n_384), .A2(n_56), .B1(n_57), .B2(n_61), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_414), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_419), .B(n_62), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_414), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_413), .A2(n_166), .B(n_158), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_426), .Y(n_474) );
XOR2x2_ASAP7_75t_L g475 ( .A(n_409), .B(n_64), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_426), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_422), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_422), .Y(n_478) );
XOR2xp5_ASAP7_75t_L g479 ( .A(n_425), .B(n_67), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_403), .B(n_68), .Y(n_480) );
OAI211xp5_ASAP7_75t_L g481 ( .A1(n_392), .A2(n_162), .B(n_166), .C(n_158), .Y(n_481) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_386), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_397), .A2(n_166), .B(n_158), .Y(n_483) );
XNOR2x1_ASAP7_75t_L g484 ( .A(n_417), .B(n_69), .Y(n_484) );
OAI211xp5_ASAP7_75t_L g485 ( .A1(n_392), .A2(n_166), .B(n_158), .C(n_73), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_399), .A2(n_71), .B(n_72), .C(n_74), .Y(n_486) );
AOI211xp5_ASAP7_75t_L g487 ( .A1(n_392), .A2(n_78), .B(n_192), .C(n_142), .Y(n_487) );
O2A1O1Ixp5_ASAP7_75t_L g488 ( .A1(n_400), .A2(n_158), .B(n_166), .C(n_392), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_401), .B(n_158), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_386), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_399), .B(n_427), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_389), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_401), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_493), .B(n_442), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_433), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_444), .B(n_451), .Y(n_496) );
AO22x2_ASAP7_75t_L g497 ( .A1(n_482), .A2(n_429), .B1(n_490), .B2(n_484), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_447), .A2(n_461), .B1(n_453), .B2(n_428), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_491), .Y(n_499) );
OAI211xp5_ASAP7_75t_SL g500 ( .A1(n_430), .A2(n_429), .B(n_488), .C(n_450), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_447), .A2(n_453), .B1(n_446), .B2(n_428), .Y(n_501) );
AOI211xp5_ASAP7_75t_L g502 ( .A1(n_489), .A2(n_466), .B(n_434), .C(n_483), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_438), .A2(n_449), .B1(n_472), .B2(n_436), .Y(n_503) );
XNOR2x1_ASAP7_75t_L g504 ( .A(n_475), .B(n_479), .Y(n_504) );
OAI211xp5_ASAP7_75t_L g505 ( .A1(n_436), .A2(n_487), .B(n_481), .C(n_464), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_492), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_469), .A2(n_486), .B(n_456), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_445), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_458), .A2(n_477), .B(n_485), .C(n_471), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_448), .B(n_457), .Y(n_510) );
XNOR2xp5_ASAP7_75t_L g511 ( .A(n_441), .B(n_432), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_497), .A2(n_438), .B1(n_431), .B2(n_452), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_497), .A2(n_468), .B1(n_462), .B2(n_467), .C(n_470), .Y(n_513) );
AOI211xp5_ASAP7_75t_L g514 ( .A1(n_500), .A2(n_460), .B(n_455), .C(n_463), .Y(n_514) );
NOR4xp25_ASAP7_75t_L g515 ( .A(n_501), .B(n_471), .C(n_480), .D(n_478), .Y(n_515) );
OAI211xp5_ASAP7_75t_L g516 ( .A1(n_502), .A2(n_463), .B(n_465), .C(n_458), .Y(n_516) );
AOI211xp5_ASAP7_75t_L g517 ( .A1(n_507), .A2(n_459), .B(n_480), .C(n_473), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_494), .Y(n_518) );
AOI211xp5_ASAP7_75t_L g519 ( .A1(n_505), .A2(n_454), .B(n_474), .C(n_476), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_495), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_508), .Y(n_521) );
NAND3xp33_ASAP7_75t_SL g522 ( .A(n_513), .B(n_503), .C(n_509), .Y(n_522) );
NAND3xp33_ASAP7_75t_SL g523 ( .A(n_512), .B(n_503), .C(n_498), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_516), .B(n_496), .C(n_510), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_517), .A2(n_504), .B(n_511), .Y(n_525) );
NOR3xp33_ASAP7_75t_SL g526 ( .A(n_517), .B(n_499), .C(n_506), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_524), .Y(n_527) );
OAI221xp5_ASAP7_75t_R g528 ( .A1(n_525), .A2(n_519), .B1(n_515), .B2(n_518), .C(n_520), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_522), .Y(n_529) );
AO22x2_ASAP7_75t_L g530 ( .A1(n_527), .A2(n_523), .B1(n_526), .B2(n_521), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_529), .A2(n_514), .B1(n_469), .B2(n_435), .C(n_437), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_530), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_531), .A2(n_527), .B1(n_528), .B2(n_469), .Y(n_533) );
INVxp67_ASAP7_75t_L g534 ( .A(n_532), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_534), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_535), .A2(n_533), .B1(n_443), .B2(n_439), .C(n_440), .Y(n_536) );
endmodule