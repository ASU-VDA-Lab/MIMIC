module fake_aes_6760_n_721 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_721);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_721;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_472;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_58), .Y(n_80) );
INVx1_ASAP7_75t_SL g81 ( .A(n_63), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_27), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_14), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_5), .Y(n_84) );
INVx2_ASAP7_75t_SL g85 ( .A(n_37), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_12), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_57), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_7), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_16), .Y(n_89) );
BUFx5_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_9), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_45), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_64), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_33), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_40), .Y(n_95) );
BUFx2_ASAP7_75t_L g96 ( .A(n_72), .Y(n_96) );
HB1xp67_ASAP7_75t_L g97 ( .A(n_20), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_11), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_13), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_38), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_67), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_30), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_11), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_69), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_12), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_62), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_71), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_24), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_36), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_6), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_59), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_21), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_3), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_73), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_19), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_74), .Y(n_116) );
INVxp33_ASAP7_75t_SL g117 ( .A(n_29), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_52), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_43), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_48), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_16), .Y(n_121) );
INVxp33_ASAP7_75t_L g122 ( .A(n_26), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_35), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_60), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_75), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_55), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_4), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_47), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_96), .B(n_0), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_104), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_90), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_90), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_90), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_90), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_91), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_96), .B(n_0), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_110), .B(n_1), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_114), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_110), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_80), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_80), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_82), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_87), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_112), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_87), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_116), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_92), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_123), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_88), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_113), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_92), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_108), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_85), .B(n_2), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g160 ( .A1(n_89), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_93), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_93), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_94), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_117), .Y(n_164) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_94), .A2(n_41), .B(n_78), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_100), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_102), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_109), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_98), .B(n_7), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_95), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_95), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_88), .Y(n_172) );
XOR2x2_ASAP7_75t_SL g173 ( .A(n_83), .B(n_8), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_169), .B(n_151), .Y(n_175) );
BUFx10_ASAP7_75t_L g176 ( .A(n_166), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_129), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_151), .B(n_122), .Y(n_180) );
INVxp67_ASAP7_75t_L g181 ( .A(n_169), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_153), .B(n_105), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_174), .B(n_128), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_165), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_169), .A2(n_97), .B1(n_103), .B2(n_83), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
INVxp67_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_174), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_158), .B(n_111), .Y(n_192) );
AND2x6_ASAP7_75t_L g193 ( .A(n_174), .B(n_128), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_167), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_172), .Y(n_196) );
CKINVDCx14_ASAP7_75t_R g197 ( .A(n_136), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_174), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_145), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_129), .Y(n_200) );
INVxp67_ASAP7_75t_L g201 ( .A(n_137), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_145), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_132), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_165), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_132), .Y(n_205) );
OR2x6_ASAP7_75t_L g206 ( .A(n_141), .B(n_127), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_145), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_153), .B(n_85), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_146), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_157), .B(n_127), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_146), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_132), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
AND2x6_ASAP7_75t_L g214 ( .A(n_157), .B(n_125), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_146), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_147), .Y(n_216) );
NAND2x1p5_ASAP7_75t_L g217 ( .A(n_161), .B(n_107), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_133), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_161), .B(n_101), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_162), .B(n_106), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_168), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_147), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_164), .B(n_106), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_147), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_148), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_162), .B(n_126), .Y(n_226) );
AND2x6_ASAP7_75t_L g227 ( .A(n_163), .B(n_105), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_148), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_148), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_165), .Y(n_230) );
OR2x6_ASAP7_75t_L g231 ( .A(n_141), .B(n_84), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_137), .B(n_84), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_163), .B(n_124), .Y(n_233) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_170), .B(n_121), .Y(n_234) );
AOI22x1_ASAP7_75t_L g235 ( .A1(n_185), .A2(n_149), .B1(n_171), .B2(n_172), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_178), .Y(n_236) );
NOR3xp33_ASAP7_75t_SL g237 ( .A(n_192), .B(n_160), .C(n_154), .Y(n_237) );
NOR2xp33_ASAP7_75t_R g238 ( .A(n_197), .B(n_150), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_234), .Y(n_239) );
INVxp67_ASAP7_75t_SL g240 ( .A(n_234), .Y(n_240) );
INVx4_ASAP7_75t_L g241 ( .A(n_227), .Y(n_241) );
BUFx4f_ASAP7_75t_L g242 ( .A(n_227), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_201), .B(n_170), .Y(n_243) );
NOR3xp33_ASAP7_75t_SL g244 ( .A(n_223), .B(n_160), .C(n_142), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_181), .A2(n_130), .B1(n_144), .B2(n_152), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_234), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_189), .B(n_172), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_176), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_178), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_190), .B(n_173), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_197), .Y(n_251) );
NAND2xp33_ASAP7_75t_L g252 ( .A(n_185), .B(n_171), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_175), .B(n_180), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_178), .Y(n_254) );
INVx6_ASAP7_75t_L g255 ( .A(n_194), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_175), .B(n_144), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_232), .B(n_131), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_185), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_206), .B(n_86), .Y(n_259) );
AND3x1_ASAP7_75t_L g260 ( .A(n_186), .B(n_173), .C(n_86), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_183), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_217), .B(n_173), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_183), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_232), .B(n_171), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_206), .B(n_99), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_184), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_183), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_187), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_199), .A2(n_149), .B(n_143), .C(n_140), .Y(n_269) );
NOR3xp33_ASAP7_75t_SL g270 ( .A(n_219), .B(n_121), .C(n_99), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_202), .A2(n_207), .B(n_229), .C(n_228), .Y(n_271) );
NAND2xp33_ASAP7_75t_SL g272 ( .A(n_185), .B(n_149), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_206), .B(n_118), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_176), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_206), .B(n_115), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_231), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_176), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_231), .B(n_115), .Y(n_278) );
INVx2_ASAP7_75t_SL g279 ( .A(n_231), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_217), .B(n_120), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_231), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_182), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_182), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_187), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_226), .B(n_143), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_195), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_184), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_221), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_187), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_217), .B(n_81), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_196), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_196), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_196), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_188), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_227), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_182), .B(n_140), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_184), .Y(n_297) );
AND2x6_ASAP7_75t_L g298 ( .A(n_185), .B(n_139), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_210), .B(n_119), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_191), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_220), .Y(n_301) );
BUFx10_ASAP7_75t_L g302 ( .A(n_227), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_241), .Y(n_303) );
BUFx10_ASAP7_75t_L g304 ( .A(n_248), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_266), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_288), .B(n_210), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_253), .B(n_210), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_240), .Y(n_308) );
BUFx8_ASAP7_75t_L g309 ( .A(n_276), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_248), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_266), .B(n_208), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_243), .B(n_220), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_262), .A2(n_227), .B1(n_214), .B2(n_233), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_297), .A2(n_220), .B1(n_198), .B2(n_194), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_300), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_300), .Y(n_316) );
NAND2xp33_ASAP7_75t_L g317 ( .A(n_295), .B(n_227), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_264), .B(n_216), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_241), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_287), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_287), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_239), .A2(n_213), .B1(n_194), .B2(n_224), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_246), .B(n_215), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_259), .B(n_214), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_241), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_282), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_258), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_242), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_283), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
INVx1_ASAP7_75t_SL g331 ( .A(n_277), .Y(n_331) );
CKINVDCx8_ASAP7_75t_R g332 ( .A(n_274), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_250), .A2(n_214), .B1(n_193), .B2(n_219), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_302), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_258), .Y(n_336) );
OR2x6_ASAP7_75t_SL g337 ( .A(n_274), .B(n_193), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_276), .A2(n_213), .B1(n_225), .B2(n_222), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_255), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_258), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_257), .B(n_213), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_242), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_294), .B(n_208), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_252), .A2(n_230), .B(n_204), .Y(n_344) );
INVxp67_ASAP7_75t_L g345 ( .A(n_259), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_302), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_255), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_279), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_258), .Y(n_349) );
INVx3_ASAP7_75t_SL g350 ( .A(n_286), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_252), .A2(n_230), .B(n_204), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_256), .A2(n_214), .B1(n_193), .B2(n_211), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_279), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_278), .A2(n_209), .B1(n_204), .B2(n_230), .Y(n_354) );
BUFx12f_ASAP7_75t_L g355 ( .A(n_286), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_302), .B(n_204), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_245), .B(n_214), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_247), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_256), .B(n_193), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_307), .B(n_256), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_315), .Y(n_362) );
OA21x2_ASAP7_75t_L g363 ( .A1(n_344), .A2(n_235), .B(n_271), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_318), .B(n_259), .Y(n_364) );
AO31x2_ASAP7_75t_L g365 ( .A1(n_354), .A2(n_269), .A3(n_281), .B(n_285), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_318), .B(n_265), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_308), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_306), .B(n_278), .Y(n_368) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_355), .A2(n_238), .B1(n_251), .B2(n_265), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_306), .B(n_251), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_330), .A2(n_260), .B1(n_244), .B2(n_237), .C(n_265), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_359), .B(n_275), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_316), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_355), .Y(n_374) );
INVx4_ASAP7_75t_L g375 ( .A(n_308), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_345), .A2(n_275), .B1(n_299), .B2(n_301), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_316), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_359), .A2(n_275), .B1(n_299), .B2(n_214), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_303), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_350), .A2(n_242), .B1(n_273), .B2(n_295), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_350), .B(n_301), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g382 ( .A1(n_357), .A2(n_270), .B(n_290), .C(n_280), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_327), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_358), .A2(n_272), .B(n_298), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_330), .B(n_299), .Y(n_385) );
AO31x2_ASAP7_75t_L g386 ( .A1(n_351), .A2(n_133), .A3(n_139), .B(n_138), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_303), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_358), .A2(n_255), .B1(n_293), .B2(n_268), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_310), .A2(n_193), .B1(n_230), .B2(n_204), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_303), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_312), .A2(n_193), .B1(n_254), .B2(n_292), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_326), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_350), .A2(n_292), .B1(n_254), .B2(n_236), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_321), .B(n_236), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_327), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_370), .A2(n_310), .B1(n_331), .B2(n_312), .Y(n_396) );
OAI21xp33_ASAP7_75t_L g397 ( .A1(n_382), .A2(n_343), .B(n_341), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_361), .A2(n_334), .B1(n_329), .B2(n_326), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_387), .Y(n_399) );
AOI211xp5_ASAP7_75t_L g400 ( .A1(n_371), .A2(n_334), .B(n_311), .C(n_329), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_364), .A2(n_352), .B1(n_337), .B2(n_321), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_369), .A2(n_332), .B1(n_333), .B2(n_313), .C(n_353), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_375), .A2(n_309), .B1(n_304), .B2(n_348), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_367), .A2(n_309), .B1(n_304), .B2(n_348), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_368), .A2(n_332), .B1(n_353), .B2(n_324), .C(n_338), .Y(n_405) );
OAI222xp33_ASAP7_75t_L g406 ( .A1(n_375), .A2(n_321), .B1(n_320), .B2(n_323), .C1(n_314), .C2(n_305), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_368), .B(n_323), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_366), .A2(n_337), .B1(n_320), .B2(n_305), .Y(n_408) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_375), .A2(n_309), .B1(n_304), .B2(n_311), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_375), .A2(n_311), .B1(n_272), .B2(n_230), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_372), .B(n_236), .Y(n_411) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_385), .A2(n_317), .B1(n_322), .B2(n_292), .C(n_254), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_378), .A2(n_317), .B1(n_235), .B2(n_347), .C(n_339), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_376), .A2(n_328), .B1(n_303), .B2(n_319), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_392), .B(n_249), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_360), .A2(n_339), .B1(n_347), .B2(n_249), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_360), .A2(n_377), .B1(n_373), .B2(n_362), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_362), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_373), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_374), .A2(n_328), .B1(n_303), .B2(n_319), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_374), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_392), .B(n_261), .Y(n_422) );
AOI222xp33_ASAP7_75t_L g423 ( .A1(n_372), .A2(n_134), .B1(n_135), .B2(n_138), .C1(n_268), .C2(n_263), .Y(n_423) );
INVx4_ASAP7_75t_SL g424 ( .A(n_394), .Y(n_424) );
OA21x2_ASAP7_75t_L g425 ( .A1(n_417), .A2(n_384), .B(n_336), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_424), .B(n_377), .Y(n_426) );
OAI33xp33_ASAP7_75t_L g427 ( .A1(n_419), .A2(n_393), .A3(n_381), .B1(n_134), .B2(n_135), .B3(n_388), .Y(n_427) );
NOR2x2_ASAP7_75t_L g428 ( .A(n_409), .B(n_383), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_407), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_418), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_404), .A2(n_380), .B1(n_384), .B2(n_328), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_417), .Y(n_432) );
OR2x6_ASAP7_75t_L g433 ( .A(n_408), .B(n_387), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_398), .B(n_365), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_398), .B(n_394), .Y(n_435) );
NOR2x1_ASAP7_75t_R g436 ( .A(n_403), .B(n_342), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_405), .A2(n_389), .B1(n_391), .B2(n_394), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_424), .B(n_394), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_424), .B(n_379), .Y(n_439) );
OAI22xp5_ASAP7_75t_SL g440 ( .A1(n_396), .A2(n_379), .B1(n_390), .B2(n_342), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_415), .Y(n_441) );
OR2x6_ASAP7_75t_L g442 ( .A(n_401), .B(n_387), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_400), .A2(n_293), .B1(n_263), .B2(n_267), .C(n_284), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_422), .B(n_365), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_416), .B(n_365), .Y(n_446) );
INVx3_ASAP7_75t_SL g447 ( .A(n_399), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_421), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_399), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_399), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_397), .B(n_390), .C(n_379), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_416), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_402), .A2(n_339), .B1(n_347), .B2(n_390), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_423), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_413), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_420), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_410), .B(n_365), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_412), .A2(n_387), .B1(n_395), .B2(n_383), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_410), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_446), .B(n_365), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_446), .B(n_399), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_444), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_429), .B(n_386), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_445), .B(n_386), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_444), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_457), .B(n_386), .Y(n_466) );
NAND4xp25_ASAP7_75t_L g467 ( .A(n_453), .B(n_414), .C(n_9), .D(n_10), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_457), .B(n_386), .Y(n_468) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_459), .A2(n_406), .B(n_336), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_434), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_434), .B(n_386), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_454), .B(n_432), .Y(n_472) );
INVx5_ASAP7_75t_L g473 ( .A(n_433), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_430), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_425), .Y(n_475) );
NOR2x1p5_ASAP7_75t_L g476 ( .A(n_456), .B(n_387), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_427), .A2(n_363), .B1(n_395), .B2(n_284), .Y(n_477) );
BUFx3_ASAP7_75t_L g478 ( .A(n_438), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_451), .B(n_363), .C(n_258), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_430), .B(n_8), .Y(n_480) );
INVx4_ASAP7_75t_L g481 ( .A(n_426), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_452), .B(n_10), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_455), .B(n_363), .C(n_340), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_426), .Y(n_484) );
INVx4_ASAP7_75t_L g485 ( .A(n_426), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_425), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_425), .B(n_13), .Y(n_487) );
BUFx3_ASAP7_75t_L g488 ( .A(n_438), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_441), .B(n_14), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_448), .B(n_363), .C(n_340), .Y(n_490) );
BUFx2_ASAP7_75t_L g491 ( .A(n_433), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_450), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_437), .A2(n_267), .B1(n_261), .B2(n_289), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_456), .B(n_15), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_435), .B(n_15), .Y(n_495) );
XOR2x1_ASAP7_75t_L g496 ( .A(n_428), .B(n_349), .Y(n_496) );
AOI211xp5_ASAP7_75t_SL g497 ( .A1(n_431), .A2(n_325), .B(n_349), .C(n_20), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_450), .Y(n_498) );
INVxp67_ASAP7_75t_SL g499 ( .A(n_449), .Y(n_499) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_458), .A2(n_289), .B(n_291), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_442), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_447), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_442), .B(n_65), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_442), .A2(n_319), .B1(n_325), .B2(n_291), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_449), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_438), .B(n_17), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_449), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_442), .B(n_17), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_481), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_474), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_472), .B(n_439), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_497), .A2(n_439), .B(n_443), .Y(n_512) );
OAI21xp5_ASAP7_75t_SL g513 ( .A1(n_497), .A2(n_428), .B(n_439), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_462), .B(n_447), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_474), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_462), .B(n_433), .Y(n_516) );
NOR3xp33_ASAP7_75t_SL g517 ( .A(n_467), .B(n_440), .C(n_436), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_494), .B(n_18), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_480), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_480), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_502), .B(n_18), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_478), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_478), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_465), .B(n_433), .Y(n_524) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_508), .B(n_356), .C(n_319), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_489), .B(n_21), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_468), .B(n_22), .Y(n_527) );
INVx3_ASAP7_75t_SL g528 ( .A(n_481), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_465), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_463), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_478), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_468), .B(n_466), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_482), .B(n_22), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_482), .B(n_23), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_464), .B(n_23), .Y(n_535) );
AO22x1_ASAP7_75t_L g536 ( .A1(n_481), .A2(n_485), .B1(n_473), .B2(n_508), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_492), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_488), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_492), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_498), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_498), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_468), .B(n_25), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_468), .B(n_28), .Y(n_543) );
OAI33xp33_ASAP7_75t_L g544 ( .A1(n_495), .A2(n_31), .A3(n_32), .B1(n_34), .B2(n_39), .B3(n_42), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_470), .B(n_44), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_470), .B(n_46), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_466), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_487), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_503), .B(n_319), .Y(n_549) );
OAI211xp5_ASAP7_75t_L g550 ( .A1(n_467), .A2(n_325), .B(n_346), .C(n_335), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_471), .B(n_49), .Y(n_551) );
OAI33xp33_ASAP7_75t_L g552 ( .A1(n_506), .A2(n_50), .A3(n_51), .B1(n_53), .B2(n_54), .B3(n_56), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_487), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_460), .B(n_61), .Y(n_554) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_483), .A2(n_200), .B(n_179), .Y(n_555) );
INVx4_ASAP7_75t_L g556 ( .A(n_481), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_484), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_471), .B(n_66), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_484), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_460), .B(n_68), .Y(n_560) );
NAND2xp33_ASAP7_75t_R g561 ( .A(n_503), .B(n_70), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_461), .B(n_76), .Y(n_562) );
AND4x1_ASAP7_75t_L g563 ( .A(n_493), .B(n_77), .C(n_79), .D(n_298), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_485), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_475), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_461), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_530), .B(n_485), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_547), .B(n_485), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_527), .A2(n_491), .B1(n_476), .B2(n_501), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_529), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_528), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_511), .B(n_496), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_537), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_532), .B(n_501), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_547), .B(n_488), .Y(n_575) );
AOI21xp33_ASAP7_75t_L g576 ( .A1(n_561), .A2(n_503), .B(n_488), .Y(n_576) );
AOI32xp33_ASAP7_75t_L g577 ( .A1(n_521), .A2(n_503), .A3(n_491), .B1(n_504), .B2(n_496), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_539), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_540), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_528), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_527), .B(n_496), .Y(n_581) );
INVx2_ASAP7_75t_SL g582 ( .A(n_556), .Y(n_582) );
OAI32xp33_ASAP7_75t_L g583 ( .A1(n_561), .A2(n_504), .A3(n_475), .B1(n_486), .B2(n_476), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_541), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_565), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_515), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_532), .B(n_486), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_566), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_566), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_518), .B(n_490), .C(n_500), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_510), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_510), .Y(n_592) );
OAI221xp5_ASAP7_75t_SL g593 ( .A1(n_513), .A2(n_500), .B1(n_475), .B2(n_486), .C(n_490), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_519), .B(n_499), .Y(n_594) );
AOI21xp33_ASAP7_75t_SL g595 ( .A1(n_536), .A2(n_469), .B(n_479), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_522), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_514), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_548), .B(n_553), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_520), .B(n_507), .Y(n_599) );
A2O1A1Ixp33_ASAP7_75t_L g600 ( .A1(n_517), .A2(n_473), .B(n_479), .C(n_505), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_557), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_559), .Y(n_602) );
AOI31xp33_ASAP7_75t_L g603 ( .A1(n_550), .A2(n_473), .A3(n_505), .B(n_507), .Y(n_603) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_549), .Y(n_604) );
O2A1O1Ixp5_ASAP7_75t_L g605 ( .A1(n_556), .A2(n_507), .B(n_505), .C(n_483), .Y(n_605) );
OAI21xp33_ASAP7_75t_L g606 ( .A1(n_526), .A2(n_477), .B(n_473), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_512), .A2(n_473), .B1(n_469), .B2(n_298), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_531), .B(n_473), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_565), .Y(n_609) );
OAI21xp5_ASAP7_75t_SL g610 ( .A1(n_564), .A2(n_469), .B(n_346), .Y(n_610) );
NAND2x1_ASAP7_75t_SL g611 ( .A(n_556), .B(n_469), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_546), .A2(n_346), .B1(n_335), .B2(n_255), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_516), .B(n_177), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_535), .B(n_560), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_509), .A2(n_346), .B1(n_335), .B2(n_200), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_560), .B(n_298), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_524), .B(n_298), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_551), .B(n_298), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_551), .B(n_177), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_558), .B(n_179), .Y(n_620) );
AND3x2_ASAP7_75t_L g621 ( .A(n_590), .B(n_542), .C(n_543), .Y(n_621) );
XOR2x2_ASAP7_75t_L g622 ( .A(n_571), .B(n_536), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_588), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_589), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_570), .Y(n_625) );
NOR3x1_ASAP7_75t_L g626 ( .A(n_582), .B(n_509), .C(n_534), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_587), .B(n_558), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_573), .Y(n_628) );
NOR2xp67_ASAP7_75t_SL g629 ( .A(n_582), .B(n_549), .Y(n_629) );
INVxp67_ASAP7_75t_L g630 ( .A(n_596), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_578), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_597), .B(n_533), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_579), .Y(n_633) );
OAI211xp5_ASAP7_75t_L g634 ( .A1(n_577), .A2(n_564), .B(n_538), .C(n_523), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_603), .B(n_564), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_584), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_580), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_593), .A2(n_543), .B(n_542), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_586), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_601), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_574), .B(n_562), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_602), .Y(n_642) );
NOR2xp33_ASAP7_75t_R g643 ( .A(n_569), .B(n_546), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_587), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_598), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_598), .Y(n_646) );
NAND2xp33_ASAP7_75t_SL g647 ( .A(n_569), .B(n_562), .Y(n_647) );
BUFx2_ASAP7_75t_L g648 ( .A(n_608), .Y(n_648) );
NOR2xp33_ASAP7_75t_SL g649 ( .A(n_576), .B(n_552), .Y(n_649) );
AOI22x1_ASAP7_75t_L g650 ( .A1(n_604), .A2(n_563), .B1(n_544), .B2(n_525), .Y(n_650) );
NOR3xp33_ASAP7_75t_L g651 ( .A(n_606), .B(n_554), .C(n_545), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_574), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_599), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_575), .B(n_555), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_572), .A2(n_555), .B1(n_335), .B2(n_346), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_568), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_600), .B(n_555), .Y(n_657) );
OAI211xp5_ASAP7_75t_SL g658 ( .A1(n_614), .A2(n_203), .B(n_205), .C(n_212), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_594), .B(n_203), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_625), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_628), .Y(n_661) );
OAI21x1_ASAP7_75t_SL g662 ( .A1(n_626), .A2(n_581), .B(n_622), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_644), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_631), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_648), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_653), .B(n_591), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_633), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_656), .A2(n_572), .B1(n_600), .B2(n_567), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_649), .B(n_607), .C(n_595), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_636), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_647), .A2(n_583), .B1(n_592), .B2(n_618), .C1(n_620), .C2(n_619), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g672 ( .A1(n_638), .A2(n_611), .B(n_610), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_637), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_630), .B(n_613), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_656), .Y(n_675) );
XOR2xp5_ASAP7_75t_L g676 ( .A(n_622), .B(n_616), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_643), .A2(n_634), .B1(n_650), .B2(n_632), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_639), .Y(n_678) );
XNOR2xp5_ASAP7_75t_L g679 ( .A(n_621), .B(n_618), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_640), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_652), .B(n_609), .Y(n_681) );
NAND2xp33_ASAP7_75t_SL g682 ( .A(n_643), .B(n_609), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_642), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_677), .A2(n_635), .B(n_647), .C(n_658), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_662), .A2(n_632), .B1(n_646), .B2(n_645), .C(n_623), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_681), .Y(n_686) );
INVx2_ASAP7_75t_SL g687 ( .A(n_673), .Y(n_687) );
OAI311xp33_ASAP7_75t_L g688 ( .A1(n_669), .A2(n_655), .A3(n_654), .B1(n_659), .C1(n_627), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_666), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_682), .A2(n_635), .B(n_657), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_665), .B(n_627), .Y(n_691) );
BUFx3_ASAP7_75t_L g692 ( .A(n_665), .Y(n_692) );
INVx1_ASAP7_75t_SL g693 ( .A(n_675), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_660), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g695 ( .A(n_674), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_661), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_663), .B(n_624), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g698 ( .A1(n_677), .A2(n_651), .B1(n_657), .B2(n_629), .C(n_605), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_664), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_668), .A2(n_641), .B1(n_612), .B2(n_585), .Y(n_700) );
AOI21xp33_ASAP7_75t_SL g701 ( .A1(n_671), .A2(n_612), .B(n_615), .Y(n_701) );
OAI22x1_ASAP7_75t_L g702 ( .A1(n_676), .A2(n_585), .B1(n_617), .B2(n_335), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_682), .A2(n_617), .B1(n_212), .B2(n_205), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_663), .Y(n_704) );
OAI211xp5_ASAP7_75t_SL g705 ( .A1(n_672), .A2(n_218), .B(n_674), .C(n_670), .Y(n_705) );
NAND3xp33_ASAP7_75t_SL g706 ( .A(n_667), .B(n_218), .C(n_678), .Y(n_706) );
OAI21xp33_ASAP7_75t_L g707 ( .A1(n_679), .A2(n_680), .B(n_683), .Y(n_707) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_684), .A2(n_698), .B1(n_695), .B2(n_700), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_690), .A2(n_706), .B(n_705), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_693), .B(n_687), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_692), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_689), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_708), .A2(n_685), .B1(n_707), .B2(n_695), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_710), .A2(n_687), .B1(n_702), .B2(n_692), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_709), .A2(n_688), .B(n_701), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g716 ( .A1(n_713), .A2(n_709), .B1(n_711), .B2(n_712), .Y(n_716) );
AOI22xp33_ASAP7_75t_R g717 ( .A1(n_715), .A2(n_689), .B1(n_696), .B2(n_699), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_717), .A2(n_714), .B1(n_716), .B2(n_703), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_717), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g720 ( .A1(n_719), .A2(n_694), .B1(n_686), .B2(n_704), .C1(n_697), .C2(n_691), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_720), .A2(n_718), .B(n_686), .Y(n_721) );
endmodule