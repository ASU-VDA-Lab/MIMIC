module fake_netlist_1_5166_n_486 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_486);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_486;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_141;
wire n_119;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g67 ( .A(n_55), .Y(n_67) );
INVxp33_ASAP7_75t_SL g68 ( .A(n_39), .Y(n_68) );
CKINVDCx20_ASAP7_75t_R g69 ( .A(n_1), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_45), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_32), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_17), .Y(n_72) );
BUFx2_ASAP7_75t_L g73 ( .A(n_36), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_19), .Y(n_74) );
INVxp33_ASAP7_75t_L g75 ( .A(n_8), .Y(n_75) );
INVxp67_ASAP7_75t_SL g76 ( .A(n_4), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_26), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_57), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_37), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_41), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_17), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_8), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_64), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_53), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_56), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_27), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_4), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_58), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_11), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_66), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_52), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_5), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_28), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_48), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_62), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_18), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_21), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_46), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_63), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_59), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_18), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_73), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_73), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_103), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_103), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_82), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_103), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_68), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_67), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_72), .B(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_70), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_75), .B(n_0), .Y(n_115) );
AND2x2_ASAP7_75t_L g116 ( .A(n_72), .B(n_74), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_79), .Y(n_117) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_71), .A2(n_1), .B(n_2), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_80), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_74), .Y(n_120) );
INVx4_ASAP7_75t_L g121 ( .A(n_83), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_84), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_71), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_81), .B(n_2), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_104), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_104), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_121), .B(n_77), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_104), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_104), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_120), .B(n_116), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_115), .A2(n_98), .B1(n_76), .B2(n_81), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_116), .B(n_87), .Y(n_132) );
OR2x2_ASAP7_75t_SL g133 ( .A(n_118), .B(n_87), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_104), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_116), .B(n_90), .Y(n_135) );
BUFx3_ASAP7_75t_L g136 ( .A(n_104), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_121), .B(n_91), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_121), .B(n_102), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_104), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_109), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_104), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_123), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_121), .B(n_102), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_123), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_123), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_123), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_130), .B(n_106), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_132), .B(n_121), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_130), .B(n_106), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_138), .B(n_114), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
NOR2xp33_ASAP7_75t_R g152 ( .A(n_140), .B(n_109), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_144), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_145), .Y(n_154) );
OR2x2_ASAP7_75t_L g155 ( .A(n_131), .B(n_115), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_142), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_132), .B(n_115), .Y(n_158) );
BUFx2_ASAP7_75t_L g159 ( .A(n_132), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_135), .A2(n_114), .B1(n_120), .B2(n_124), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_142), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
BUFx4f_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_145), .B(n_120), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_145), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_131), .B(n_108), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_143), .B(n_108), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_142), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
BUFx8_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_150), .A2(n_137), .B(n_127), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_157), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_151), .B(n_105), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
AOI222xp33_ASAP7_75t_L g181 ( .A1(n_171), .A2(n_69), .B1(n_99), .B2(n_113), .C1(n_124), .C2(n_111), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_168), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
AOI22xp5_ASAP7_75t_SL g186 ( .A1(n_151), .A2(n_118), .B1(n_111), .B2(n_113), .Y(n_186) );
CKINVDCx11_ASAP7_75t_R g187 ( .A(n_171), .Y(n_187) );
BUFx2_ASAP7_75t_SL g188 ( .A(n_163), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_168), .B(n_118), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_157), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_172), .B(n_112), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_150), .A2(n_128), .B(n_141), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_153), .A2(n_128), .B(n_141), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_168), .Y(n_195) );
INVx5_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
INVx2_ASAP7_75t_SL g197 ( .A(n_168), .Y(n_197) );
NOR2xp33_ASAP7_75t_SL g198 ( .A(n_168), .B(n_121), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_175), .A2(n_114), .B1(n_118), .B2(n_146), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_166), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_175), .A2(n_118), .B1(n_146), .B2(n_107), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_176), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_166), .Y(n_203) );
INVx1_ASAP7_75t_SL g204 ( .A(n_152), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_147), .B(n_112), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_163), .B(n_119), .Y(n_206) );
OAI21x1_ASAP7_75t_L g207 ( .A1(n_194), .A2(n_167), .B(n_162), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_186), .A2(n_161), .B(n_148), .C(n_165), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g209 ( .A1(n_200), .A2(n_161), .B1(n_160), .B2(n_159), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_193), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_181), .A2(n_163), .B1(n_158), .B2(n_159), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_184), .B(n_158), .Y(n_212) );
AO22x1_ASAP7_75t_L g213 ( .A1(n_204), .A2(n_176), .B1(n_171), .B2(n_147), .Y(n_213) );
NAND2xp33_ASAP7_75t_SL g214 ( .A(n_200), .B(n_163), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_202), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_202), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_187), .Y(n_217) );
OR2x6_ASAP7_75t_L g218 ( .A(n_188), .B(n_159), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_199), .A2(n_148), .B(n_170), .Y(n_219) );
AOI221xp5_ASAP7_75t_L g220 ( .A1(n_191), .A2(n_149), .B1(n_171), .B2(n_158), .C(n_155), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_203), .A2(n_160), .B1(n_164), .B2(n_165), .Y(n_221) );
OAI221xp5_ASAP7_75t_L g222 ( .A1(n_205), .A2(n_149), .B1(n_155), .B2(n_160), .C(n_164), .Y(n_222) );
AOI222xp33_ASAP7_75t_L g223 ( .A1(n_179), .A2(n_171), .B1(n_172), .B2(n_169), .C1(n_94), .C2(n_90), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_205), .A2(n_155), .B(n_169), .C(n_172), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_185), .A2(n_165), .B1(n_154), .B2(n_156), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_179), .A2(n_119), .B1(n_122), .B2(n_117), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_184), .A2(n_122), .B1(n_154), .B2(n_156), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_195), .B(n_154), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_185), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_188), .A2(n_154), .B1(n_156), .B2(n_176), .Y(n_230) );
INVxp67_ASAP7_75t_L g231 ( .A(n_195), .Y(n_231) );
BUFx8_ASAP7_75t_SL g232 ( .A(n_217), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_218), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_211), .A2(n_182), .B1(n_197), .B2(n_206), .Y(n_234) );
OAI211xp5_ASAP7_75t_SL g235 ( .A1(n_226), .A2(n_94), .B(n_110), .C(n_107), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_224), .A2(n_186), .B(n_199), .Y(n_236) );
OAI21xp5_ASAP7_75t_SL g237 ( .A1(n_211), .A2(n_197), .B(n_182), .Y(n_237) );
AOI221xp5_ASAP7_75t_L g238 ( .A1(n_222), .A2(n_177), .B1(n_203), .B2(n_107), .C(n_110), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_220), .A2(n_196), .B1(n_198), .B2(n_156), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_210), .B(n_196), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_223), .A2(n_196), .B1(n_198), .B2(n_156), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_208), .A2(n_201), .B1(n_196), .B2(n_189), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_209), .B(n_201), .Y(n_243) );
OAI211xp5_ASAP7_75t_L g244 ( .A1(n_208), .A2(n_110), .B(n_196), .C(n_86), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_219), .A2(n_189), .B(n_192), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_229), .Y(n_246) );
OAI221xp5_ASAP7_75t_L g247 ( .A1(n_212), .A2(n_189), .B1(n_196), .B2(n_154), .C(n_170), .Y(n_247) );
OAI221xp5_ASAP7_75t_L g248 ( .A1(n_225), .A2(n_77), .B1(n_78), .B2(n_85), .C(n_88), .Y(n_248) );
OAI211xp5_ASAP7_75t_SL g249 ( .A1(n_227), .A2(n_78), .B(n_85), .C(n_88), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_218), .A2(n_183), .B1(n_180), .B2(n_178), .Y(n_250) );
OAI21xp33_ASAP7_75t_L g251 ( .A1(n_230), .A2(n_146), .B(n_92), .Y(n_251) );
OAI221xp5_ASAP7_75t_SL g252 ( .A1(n_237), .A2(n_218), .B1(n_231), .B2(n_225), .C(n_215), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_236), .A2(n_207), .B(n_221), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_233), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_246), .B(n_213), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_235), .A2(n_214), .B1(n_216), .B2(n_215), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_246), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_243), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_233), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_233), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_243), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_250), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_249), .A2(n_214), .B1(n_216), .B2(n_217), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_237), .B(n_118), .Y(n_264) );
NOR2xp33_ASAP7_75t_SL g265 ( .A(n_242), .B(n_176), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_245), .B(n_146), .Y(n_266) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_244), .A2(n_89), .B(n_92), .Y(n_267) );
AOI31xp33_ASAP7_75t_SL g268 ( .A1(n_234), .A2(n_3), .A3(n_5), .B(n_6), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_247), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_251), .Y(n_270) );
OAI33xp33_ASAP7_75t_L g271 ( .A1(n_251), .A2(n_101), .A3(n_93), .B1(n_95), .B2(n_96), .B3(n_97), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_261), .B(n_248), .Y(n_272) );
INVxp67_ASAP7_75t_SL g273 ( .A(n_262), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_261), .B(n_238), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_258), .B(n_239), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_258), .B(n_89), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_257), .Y(n_277) );
AOI211xp5_ASAP7_75t_L g278 ( .A1(n_268), .A2(n_240), .B(n_95), .C(n_96), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_257), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_257), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_258), .B(n_241), .Y(n_281) );
OAI222xp33_ASAP7_75t_L g282 ( .A1(n_252), .A2(n_101), .B1(n_100), .B2(n_97), .C1(n_93), .C2(n_228), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_259), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_259), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_266), .B(n_146), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_264), .B(n_100), .Y(n_286) );
OAI33xp33_ASAP7_75t_L g287 ( .A1(n_255), .A2(n_3), .A3(n_6), .B1(n_7), .B2(n_9), .B3(n_10), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_255), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_259), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_254), .Y(n_290) );
OAI31xp33_ASAP7_75t_SL g291 ( .A1(n_264), .A2(n_232), .A3(n_9), .B(n_10), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_264), .A2(n_176), .B1(n_232), .B2(n_146), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_262), .Y(n_293) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_253), .A2(n_173), .B(n_174), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_254), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_260), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_260), .Y(n_298) );
OAI31xp33_ASAP7_75t_L g299 ( .A1(n_252), .A2(n_7), .A3(n_11), .B(n_12), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_277), .B(n_266), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_288), .B(n_262), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_277), .B(n_266), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_277), .B(n_280), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_280), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_283), .Y(n_305) );
BUFx2_ASAP7_75t_SL g306 ( .A(n_289), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_288), .B(n_262), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_280), .B(n_253), .Y(n_308) );
NOR3xp33_ASAP7_75t_L g309 ( .A(n_287), .B(n_271), .C(n_268), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_279), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_293), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_279), .B(n_270), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_296), .B(n_270), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_286), .B(n_269), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_286), .B(n_269), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_289), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_296), .B(n_265), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_290), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_290), .Y(n_319) );
OAI33xp33_ASAP7_75t_L g320 ( .A1(n_295), .A2(n_269), .A3(n_13), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_293), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_297), .B(n_265), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_293), .B(n_269), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_273), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_283), .Y(n_325) );
AND2x2_ASAP7_75t_SL g326 ( .A(n_284), .B(n_263), .Y(n_326) );
NOR2xp67_ASAP7_75t_L g327 ( .A(n_289), .B(n_12), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_276), .B(n_295), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_276), .B(n_267), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_297), .B(n_267), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_298), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_276), .B(n_267), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_298), .B(n_267), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_275), .B(n_267), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_284), .B(n_285), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_285), .B(n_13), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_275), .B(n_281), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_281), .B(n_263), .Y(n_339) );
OR2x4_ASAP7_75t_L g340 ( .A(n_291), .B(n_271), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_299), .A2(n_256), .B1(n_190), .B2(n_183), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_339), .A2(n_278), .B1(n_287), .B2(n_292), .Y(n_342) );
OAI221xp5_ASAP7_75t_L g343 ( .A1(n_341), .A2(n_291), .B1(n_299), .B2(n_278), .C(n_339), .Y(n_343) );
NAND2xp33_ASAP7_75t_L g344 ( .A(n_309), .B(n_272), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_318), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_318), .Y(n_346) );
NAND2x1_ASAP7_75t_L g347 ( .A(n_316), .B(n_285), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_319), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_338), .B(n_272), .Y(n_349) );
NAND2xp33_ASAP7_75t_L g350 ( .A(n_305), .B(n_282), .Y(n_350) );
AND2x4_ASAP7_75t_SL g351 ( .A(n_337), .B(n_335), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_338), .B(n_274), .Y(n_352) );
NOR3xp33_ASAP7_75t_L g353 ( .A(n_320), .B(n_282), .C(n_274), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_337), .B(n_273), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_328), .B(n_294), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_328), .B(n_294), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_319), .A2(n_256), .B1(n_294), .B2(n_139), .C(n_134), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_310), .Y(n_358) );
OAI21xp33_ASAP7_75t_L g359 ( .A1(n_316), .A2(n_125), .B(n_126), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_310), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_336), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
AOI21xp33_ASAP7_75t_SL g363 ( .A1(n_326), .A2(n_14), .B(n_15), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_331), .B(n_333), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_340), .A2(n_294), .B(n_190), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_335), .B(n_16), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_304), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_340), .A2(n_190), .B1(n_183), .B2(n_180), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_311), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_304), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_303), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_340), .A2(n_125), .B1(n_126), .B2(n_129), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_300), .B(n_19), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_312), .Y(n_374) );
AOI31xp33_ASAP7_75t_L g375 ( .A1(n_336), .A2(n_20), .A3(n_21), .B(n_22), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_312), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_313), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_326), .A2(n_157), .B1(n_183), .B2(n_180), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_313), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_326), .A2(n_157), .B1(n_183), .B2(n_180), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_330), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_330), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_300), .B(n_20), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_333), .B(n_22), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_302), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_302), .Y(n_386) );
OAI32xp33_ASAP7_75t_L g387 ( .A1(n_325), .A2(n_23), .A3(n_25), .B1(n_29), .B2(n_30), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_301), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_301), .Y(n_389) );
OAI21xp5_ASAP7_75t_SL g390 ( .A1(n_329), .A2(n_23), .B(n_190), .Y(n_390) );
NOR3xp33_ASAP7_75t_L g391 ( .A(n_375), .B(n_327), .C(n_334), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_351), .B(n_361), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_349), .B(n_325), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_352), .B(n_334), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_374), .Y(n_395) );
INVx5_ASAP7_75t_SL g396 ( .A(n_354), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_376), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_345), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_346), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_348), .Y(n_400) );
INVxp67_ASAP7_75t_L g401 ( .A(n_344), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_377), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_379), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_388), .B(n_308), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_389), .B(n_308), .Y(n_405) );
NAND3xp33_ASAP7_75t_L g406 ( .A(n_344), .B(n_332), .C(n_329), .Y(n_406) );
OAI21xp5_ASAP7_75t_SL g407 ( .A1(n_390), .A2(n_337), .B(n_317), .Y(n_407) );
NOR4xp25_ASAP7_75t_SL g408 ( .A(n_363), .B(n_306), .C(n_317), .D(n_322), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_383), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_364), .B(n_308), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_362), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_381), .B(n_308), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_347), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_382), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_385), .B(n_307), .Y(n_415) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_350), .B(n_306), .Y(n_416) );
NAND2xp33_ASAP7_75t_SL g417 ( .A(n_383), .B(n_322), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_354), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_386), .B(n_307), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_371), .B(n_323), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_368), .B(n_324), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_358), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_360), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_366), .B(n_323), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_350), .A2(n_314), .B(n_315), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_367), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_354), .B(n_323), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_370), .Y(n_428) );
XNOR2xp5_ASAP7_75t_L g429 ( .A(n_373), .B(n_315), .Y(n_429) );
NAND2x1_ASAP7_75t_L g430 ( .A(n_369), .B(n_324), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_394), .B(n_356), .Y(n_431) );
AOI221x1_ASAP7_75t_L g432 ( .A1(n_391), .A2(n_353), .B1(n_365), .B2(n_384), .C(n_359), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_394), .B(n_355), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_414), .B(n_369), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_414), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_425), .B(n_342), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_430), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_401), .A2(n_343), .B1(n_353), .B2(n_372), .C(n_387), .Y(n_438) );
AOI322xp5_ASAP7_75t_L g439 ( .A1(n_401), .A2(n_380), .A3(n_378), .B1(n_314), .B2(n_357), .C1(n_324), .C2(n_321), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_426), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_406), .A2(n_380), .B1(n_321), .B2(n_311), .C(n_129), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_393), .B(n_321), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_407), .A2(n_311), .B(n_190), .Y(n_443) );
XOR2x2_ASAP7_75t_L g444 ( .A(n_391), .B(n_31), .Y(n_444) );
AOI21xp33_ASAP7_75t_L g445 ( .A1(n_416), .A2(n_33), .B(n_34), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_395), .B(n_38), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_392), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_410), .B(n_40), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_404), .B(n_42), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_409), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_413), .Y(n_451) );
NOR3xp33_ASAP7_75t_L g452 ( .A(n_417), .B(n_174), .C(n_173), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_428), .Y(n_453) );
OAI31xp33_ASAP7_75t_L g454 ( .A1(n_413), .A2(n_136), .A3(n_44), .B(n_47), .Y(n_454) );
AOI211xp5_ASAP7_75t_L g455 ( .A1(n_438), .A2(n_429), .B(n_418), .C(n_421), .Y(n_455) );
NOR2xp33_ASAP7_75t_R g456 ( .A(n_436), .B(n_418), .Y(n_456) );
OAI211xp5_ASAP7_75t_SL g457 ( .A1(n_439), .A2(n_421), .B(n_402), .C(n_403), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_451), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_431), .A2(n_397), .B1(n_399), .B2(n_400), .C(n_423), .Y(n_459) );
NOR2xp33_ASAP7_75t_R g460 ( .A(n_450), .B(n_447), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g461 ( .A1(n_432), .A2(n_408), .B(n_412), .C(n_405), .Y(n_461) );
NOR2xp67_ASAP7_75t_SL g462 ( .A(n_448), .B(n_396), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_434), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_452), .B(n_396), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_431), .B(n_420), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g466 ( .A1(n_433), .A2(n_419), .B1(n_415), .B2(n_422), .C(n_398), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_445), .A2(n_427), .B(n_424), .C(n_411), .Y(n_467) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_444), .A2(n_162), .B1(n_178), .B2(n_136), .C(n_51), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_445), .A2(n_136), .B(n_49), .C(n_50), .Y(n_469) );
OR3x2_ASAP7_75t_L g470 ( .A(n_435), .B(n_43), .C(n_54), .Y(n_470) );
OAI211xp5_ASAP7_75t_L g471 ( .A1(n_454), .A2(n_178), .B(n_60), .C(n_61), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_440), .A2(n_65), .B1(n_453), .B2(n_442), .C(n_434), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_443), .A2(n_441), .B1(n_437), .B2(n_449), .Y(n_473) );
OAI321xp33_ASAP7_75t_L g474 ( .A1(n_446), .A2(n_401), .A3(n_436), .B1(n_438), .B2(n_406), .C(n_451), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_458), .B(n_474), .Y(n_475) );
NOR4xp25_ASAP7_75t_L g476 ( .A(n_457), .B(n_461), .C(n_466), .D(n_471), .Y(n_476) );
OAI211xp5_ASAP7_75t_SL g477 ( .A1(n_455), .A2(n_472), .B(n_468), .C(n_467), .Y(n_477) );
INVx1_ASAP7_75t_SL g478 ( .A(n_460), .Y(n_478) );
INVx5_ASAP7_75t_L g479 ( .A(n_478), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_476), .B(n_475), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_477), .A2(n_457), .B1(n_473), .B2(n_456), .C(n_459), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_479), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_480), .Y(n_483) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_482), .A2(n_481), .B1(n_464), .B2(n_462), .C(n_469), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_484), .A2(n_482), .B1(n_483), .B2(n_470), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_485), .A2(n_463), .B(n_465), .Y(n_486) );
endmodule