module real_jpeg_28103_n_11 (n_5, n_4, n_8, n_0, n_251, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_251;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_244;
wire n_213;
wire n_179;
wire n_128;
wire n_216;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_50),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_0),
.A2(n_36),
.B1(n_37),
.B2(n_50),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_0),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_213)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_1),
.Y(n_100)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_1),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_5),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_5),
.A2(n_19),
.B1(n_28),
.B2(n_29),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_19),
.B1(n_43),
.B2(n_44),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_5),
.A2(n_19),
.B1(n_36),
.B2(n_37),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_SL g111 ( 
.A1(n_5),
.A2(n_25),
.B(n_29),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_72),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g134 ( 
.A1(n_5),
.A2(n_6),
.B(n_37),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_5),
.B(n_65),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_5),
.A2(n_8),
.B(n_28),
.C(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_35)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_46),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_194)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_80),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_78),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_66),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_14),
.B(n_66),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_17),
.C(n_61),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_15),
.A2(n_16),
.B1(n_17),
.B2(n_60),
.Y(n_243)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_60),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_58),
.C(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_17),
.B(n_47),
.C(n_58),
.Y(n_77)
);

AOI211xp5_ASAP7_75t_L g88 ( 
.A1(n_17),
.A2(n_89),
.B(n_91),
.C(n_95),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_17),
.A2(n_60),
.B1(n_92),
.B2(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_17),
.A2(n_60),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_17),
.A2(n_60),
.B1(n_208),
.B2(n_209),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_17),
.A2(n_60),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_17),
.A2(n_208),
.B(n_228),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_22),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_18),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_19),
.A2(n_20),
.B(n_26),
.C(n_111),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_19),
.A2(n_39),
.B(n_44),
.C(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_19),
.B(n_35),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_19),
.B(n_147),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_19),
.A2(n_43),
.B(n_55),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_20),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_28),
.A2(n_29),
.B1(n_53),
.B2(n_55),
.Y(n_56)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_32),
.A2(n_58),
.B1(n_62),
.B2(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_45),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_34),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_35),
.A2(n_40),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_35),
.A2(n_40),
.B1(n_45),
.B2(n_213),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_36),
.B(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_37),
.B(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_44),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_56),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_92),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_60),
.B(n_92),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_61),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_62),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_76),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_77),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_235),
.A3(n_244),
.B1(n_247),
.B2(n_248),
.C(n_251),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_219),
.B(n_234),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_200),
.B(n_218),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_126),
.B(n_182),
.C(n_199),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_116),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_85),
.B(n_116),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_105),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_96),
.B2(n_97),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_87),
.B(n_97),
.C(n_105),
.Y(n_183)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_94),
.B1(n_98),
.B2(n_104),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_89),
.A2(n_94),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_89),
.A2(n_94),
.B1(n_133),
.B2(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_112),
.C(n_137),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_89),
.A2(n_94),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_89),
.B(n_165),
.C(n_171),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_89),
.B(n_98),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_89),
.A2(n_94),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_89),
.B(n_191),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_90),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_92),
.A2(n_94),
.B(n_159),
.C(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_92),
.A2(n_93),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_112),
.C(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_93),
.A2(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_93),
.B(n_225),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_95),
.A2(n_115),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_95),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_100),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_99),
.A2(n_103),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_115),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_106),
.A2(n_107),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_106),
.A2(n_107),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_113),
.B1(n_136),
.B2(n_139),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_112),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_113),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_112),
.A2(n_113),
.B1(n_124),
.B2(n_125),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_112),
.B(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_149),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_123),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_117),
.A2(n_118),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_119),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_120),
.B1(n_155),
.B2(n_159),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_123),
.Y(n_178)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_181),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_174),
.B(n_180),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_161),
.B(n_173),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_152),
.B(n_160),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_140),
.B(n_151),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_135),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_133),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_164),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_170),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_176),
.Y(n_180)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_184),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_197),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_189),
.B1(n_195),
.B2(n_196),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_189),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_195),
.C(n_197),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_198),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_202),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_215),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_207),
.C(n_215),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_205),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_216),
.B(n_217),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_214),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_211),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_211),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_221),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_232),
.B2(n_233),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_227),
.C(n_233),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_237),
.C(n_241),
.Y(n_236)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_226),
.B(n_237),
.CI(n_241),
.CON(n_246),
.SN(n_246)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_230),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_242),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_242),
.Y(n_248)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_246),
.Y(n_250)
);


endmodule