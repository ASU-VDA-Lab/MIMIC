module fake_jpeg_21142_n_252 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_R g43 ( 
.A(n_34),
.B(n_1),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_46),
.Y(n_71)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_32),
.Y(n_52)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_30),
.B1(n_23),
.B2(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_20),
.Y(n_66)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_49),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_3),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_62),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_67),
.B(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_55),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_30),
.B1(n_23),
.B2(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_47),
.B1(n_44),
.B2(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_70),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_30),
.B1(n_23),
.B2(n_17),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_68),
.B1(n_21),
.B2(n_33),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_66),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_18),
.B1(n_33),
.B2(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_22),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_31),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_31),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_26),
.C(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_51),
.Y(n_104)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_82),
.Y(n_120)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2x1_ASAP7_75t_R g116 ( 
.A(n_83),
.B(n_88),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_93),
.Y(n_122)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_19),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_72),
.B1(n_78),
.B2(n_25),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_18),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_106),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_100),
.Y(n_119)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_104),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_35),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_64),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_41),
.B1(n_40),
.B2(n_29),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_67),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_25),
.B1(n_21),
.B2(n_19),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_123),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_126),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_53),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_135),
.B(n_110),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_71),
.B1(n_75),
.B2(n_72),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_118),
.B1(n_133),
.B2(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_58),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_58),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_86),
.B(n_35),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_19),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_92),
.A2(n_24),
.B1(n_26),
.B2(n_6),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_107),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_90),
.C(n_108),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_157),
.C(n_115),
.Y(n_181)
);

OAI22x1_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_91),
.B1(n_109),
.B2(n_60),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_152),
.B1(n_133),
.B2(n_126),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_122),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_143),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_149),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_135),
.A2(n_100),
.B1(n_79),
.B2(n_80),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_89),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_81),
.B1(n_99),
.B2(n_24),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_150),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_26),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_12),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_96),
.B(n_81),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_4),
.B(n_5),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_12),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_161),
.B(n_16),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_156),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_162),
.B(n_166),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_174),
.B1(n_144),
.B2(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_118),
.B1(n_125),
.B2(n_128),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_179),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_115),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_158),
.B1(n_148),
.B2(n_161),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_172),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_134),
.C(n_121),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_136),
.C(n_147),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_146),
.B(n_139),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_187),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_141),
.B1(n_152),
.B2(n_137),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_188),
.A2(n_195),
.B1(n_196),
.B2(n_201),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_137),
.Y(n_189)
);

OAI322xp33_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_163),
.A3(n_174),
.B1(n_166),
.B2(n_162),
.C1(n_176),
.C2(n_168),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_153),
.B(n_141),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_165),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_194),
.C(n_200),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_144),
.B1(n_121),
.B2(n_111),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_164),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_111),
.B1(n_132),
.B2(n_157),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_179),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_204),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_177),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_171),
.B1(n_173),
.B2(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_151),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_211),
.A2(n_192),
.B(n_185),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_165),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_215),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_107),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_192),
.C(n_185),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_189),
.B1(n_198),
.B2(n_191),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_221),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_205),
.A2(n_198),
.B(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_223),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_190),
.Y(n_223)
);

NOR3xp33_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_15),
.C(n_11),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_14),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_212),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_229),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_206),
.C(n_204),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_203),
.B1(n_214),
.B2(n_202),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_231),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_216),
.B(n_206),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_221),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_220),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_236),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_217),
.B(n_216),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_239),
.B(n_14),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_224),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_229),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_244),
.B(n_243),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_247),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_235),
.C(n_7),
.Y(n_247)
);

NOR4xp25_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_6),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_248),
.C(n_7),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_9),
.Y(n_252)
);


endmodule