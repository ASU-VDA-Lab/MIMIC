module fake_netlist_5_57_n_7687 (n_924, n_1263, n_977, n_1378, n_611, n_1126, n_1423, n_1729, n_1166, n_1751, n_469, n_1508, n_82, n_785, n_549, n_532, n_1161, n_1859, n_1677, n_1150, n_226, n_1780, n_1488, n_667, n_790, n_1055, n_1501, n_111, n_880, n_544, n_1007, n_155, n_552, n_1528, n_1370, n_1292, n_1198, n_1360, n_1099, n_956, n_564, n_423, n_1738, n_21, n_105, n_1021, n_4, n_551, n_1323, n_1466, n_688, n_1695, n_1353, n_800, n_1347, n_1535, n_1789, n_1666, n_671, n_819, n_1451, n_1022, n_915, n_1545, n_864, n_173, n_859, n_951, n_1264, n_447, n_247, n_1494, n_292, n_625, n_854, n_1462, n_1799, n_1580, n_674, n_417, n_1806, n_516, n_933, n_1152, n_497, n_1869, n_1607, n_1563, n_606, n_275, n_26, n_877, n_2, n_1696, n_755, n_1118, n_6, n_1686, n_947, n_1285, n_373, n_307, n_1860, n_1359, n_530, n_87, n_150, n_1107, n_1728, n_556, n_1230, n_668, n_375, n_301, n_1896, n_929, n_1124, n_1818, n_902, n_1576, n_191, n_1104, n_1294, n_659, n_51, n_1705, n_1257, n_171, n_1182, n_579, n_1698, n_1261, n_938, n_1098, n_320, n_1154, n_1242, n_1135, n_24, n_406, n_519, n_1016, n_1243, n_546, n_101, n_1280, n_1845, n_281, n_240, n_291, n_231, n_257, n_731, n_371, n_1483, n_1314, n_1512, n_709, n_1490, n_317, n_1236, n_1633, n_569, n_1778, n_227, n_920, n_1289, n_1517, n_94, n_335, n_1669, n_370, n_976, n_343, n_1449, n_308, n_1566, n_297, n_156, n_1078, n_1670, n_775, n_219, n_157, n_600, n_1484, n_1374, n_1328, n_223, n_264, n_1877, n_1831, n_1598, n_1723, n_955, n_1850, n_163, n_339, n_1146, n_882, n_183, n_243, n_1036, n_1097, n_1749, n_347, n_59, n_550, n_696, n_897, n_215, n_350, n_196, n_798, n_646, n_1428, n_436, n_1394, n_1414, n_1216, n_290, n_580, n_1040, n_1872, n_1852, n_578, n_926, n_344, n_1218, n_422, n_475, n_777, n_1070, n_1547, n_1030, n_72, n_1755, n_415, n_1071, n_485, n_1165, n_1267, n_1561, n_496, n_1801, n_1391, n_958, n_1034, n_670, n_1513, n_1600, n_48, n_521, n_663, n_845, n_1862, n_673, n_837, n_1239, n_528, n_1796, n_680, n_1473, n_1587, n_395, n_164, n_553, n_901, n_813, n_1521, n_1284, n_1590, n_214, n_1748, n_1672, n_675, n_888, n_1880, n_1167, n_1626, n_637, n_1384, n_1556, n_184, n_446, n_1863, n_1064, n_144, n_858, n_114, n_96, n_923, n_691, n_1151, n_881, n_1405, n_1706, n_468, n_213, n_129, n_342, n_464, n_363, n_1582, n_197, n_1069, n_1784, n_1075, n_1836, n_1450, n_1322, n_1471, n_1750, n_1459, n_460, n_889, n_973, n_1700, n_477, n_571, n_1585, n_461, n_1599, n_1211, n_1197, n_1523, n_907, n_1447, n_1377, n_190, n_989, n_1039, n_34, n_228, n_283, n_1403, n_488, n_736, n_892, n_1000, n_1202, n_1278, n_1002, n_1463, n_1581, n_49, n_310, n_54, n_593, n_12, n_748, n_586, n_1058, n_1667, n_838, n_332, n_1053, n_1224, n_349, n_1248, n_230, n_1331, n_953, n_279, n_1014, n_1241, n_70, n_289, n_963, n_1052, n_954, n_627, n_1385, n_440, n_793, n_478, n_1819, n_476, n_1527, n_534, n_1882, n_884, n_345, n_944, n_1754, n_1623, n_1854, n_91, n_1565, n_1809, n_1856, n_182, n_143, n_647, n_237, n_407, n_1072, n_832, n_857, n_207, n_561, n_1319, n_1825, n_1883, n_1906, n_1712, n_1387, n_1532, n_18, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_686, n_847, n_1393, n_596, n_1775, n_1368, n_558, n_702, n_1276, n_822, n_1412, n_1709, n_728, n_266, n_1162, n_272, n_1538, n_1838, n_1199, n_1847, n_1779, n_352, n_1884, n_53, n_1038, n_520, n_1369, n_409, n_1841, n_1660, n_887, n_1905, n_154, n_71, n_300, n_809, n_870, n_931, n_599, n_1711, n_1662, n_1891, n_1481, n_434, n_1544, n_868, n_639, n_914, n_411, n_414, n_1629, n_1293, n_965, n_1876, n_1743, n_935, n_121, n_1175, n_817, n_360, n_36, n_1479, n_1810, n_64, n_1888, n_759, n_1892, n_28, n_806, n_1766, n_1477, n_324, n_1635, n_1571, n_187, n_1189, n_103, n_97, n_11, n_7, n_1259, n_1690, n_706, n_746, n_1649, n_747, n_52, n_784, n_110, n_1733, n_1244, n_431, n_1194, n_1815, n_615, n_851, n_1759, n_843, n_1788, n_523, n_913, n_1537, n_705, n_865, n_61, n_678, n_697, n_127, n_1222, n_75, n_1679, n_776, n_1798, n_1790, n_1415, n_367, n_452, n_525, n_1260, n_1746, n_1647, n_1829, n_1464, n_649, n_547, n_43, n_1444, n_1191, n_1674, n_1833, n_116, n_1830, n_1710, n_284, n_1128, n_139, n_1734, n_744, n_590, n_629, n_1308, n_1767, n_254, n_1680, n_1233, n_23, n_1615, n_1529, n_526, n_1916, n_293, n_372, n_677, n_244, n_47, n_1333, n_1121, n_314, n_368, n_433, n_604, n_8, n_949, n_100, n_1443, n_1008, n_946, n_1539, n_1001, n_1503, n_498, n_1468, n_1559, n_1765, n_1866, n_689, n_738, n_1624, n_640, n_1510, n_252, n_624, n_1380, n_1744, n_1617, n_295, n_133, n_1010, n_1231, n_739, n_1279, n_1406, n_1195, n_1837, n_1839, n_610, n_1760, n_936, n_568, n_1500, n_39, n_1090, n_757, n_633, n_439, n_106, n_1832, n_259, n_448, n_1851, n_758, n_999, n_93, n_1656, n_1158, n_1509, n_1874, n_563, n_1145, n_878, n_524, n_204, n_394, n_1678, n_1049, n_1153, n_741, n_1639, n_1306, n_1068, n_1871, n_122, n_331, n_10, n_906, n_1163, n_1207, n_919, n_908, n_90, n_724, n_1781, n_658, n_1740, n_1362, n_1586, n_456, n_959, n_535, n_152, n_940, n_1445, n_9, n_1492, n_1923, n_1773, n_592, n_1169, n_45, n_1596, n_1692, n_1017, n_123, n_978, n_1434, n_1054, n_1474, n_1665, n_1269, n_1095, n_1828, n_1614, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_603, n_1431, n_484, n_1593, n_1033, n_442, n_131, n_636, n_660, n_1640, n_1732, n_1009, n_1148, n_109, n_742, n_750, n_995, n_454, n_1609, n_374, n_185, n_396, n_1887, n_1383, n_1073, n_255, n_662, n_459, n_218, n_962, n_1215, n_1171, n_1578, n_723, n_1920, n_1065, n_1592, n_1336, n_1721, n_1758, n_1574, n_473, n_1921, n_1309, n_1878, n_1426, n_1043, n_355, n_486, n_1800, n_1548, n_614, n_337, n_1421, n_88, n_1286, n_1177, n_1355, n_168, n_974, n_727, n_1159, n_957, n_773, n_208, n_142, n_743, n_299, n_303, n_296, n_613, n_1119, n_1240, n_1820, n_65, n_829, n_1612, n_1416, n_1724, n_361, n_700, n_1237, n_573, n_69, n_1420, n_1132, n_388, n_1366, n_1300, n_1127, n_761, n_1785, n_1568, n_1006, n_329, n_274, n_1270, n_1664, n_1486, n_582, n_1332, n_1390, n_73, n_19, n_1870, n_309, n_30, n_512, n_1591, n_84, n_130, n_322, n_1682, n_1249, n_652, n_1111, n_1365, n_25, n_1349, n_1093, n_288, n_1031, n_263, n_609, n_1041, n_1265, n_1909, n_44, n_224, n_1562, n_383, n_834, n_112, n_765, n_893, n_1015, n_1140, n_891, n_1651, n_239, n_630, n_1902, n_55, n_1913, n_504, n_1823, n_511, n_874, n_358, n_1101, n_77, n_102, n_1106, n_1456, n_1875, n_1304, n_1324, n_987, n_1846, n_261, n_174, n_1885, n_1455, n_767, n_993, n_1903, n_1407, n_1551, n_545, n_441, n_860, n_450, n_1805, n_1816, n_429, n_948, n_1217, n_628, n_365, n_1849, n_729, n_1131, n_1084, n_970, n_911, n_1430, n_83, n_513, n_1094, n_1354, n_560, n_1534, n_340, n_1351, n_1044, n_1205, n_346, n_1209, n_1552, n_495, n_602, n_574, n_1435, n_879, n_16, n_58, n_623, n_405, n_824, n_359, n_1645, n_490, n_1327, n_996, n_921, n_1684, n_233, n_1717, n_572, n_366, n_815, n_1795, n_128, n_1821, n_120, n_327, n_135, n_1381, n_1611, n_1037, n_1080, n_1274, n_1316, n_1708, n_426, n_1438, n_1082, n_1840, n_589, n_716, n_1630, n_562, n_1436, n_62, n_1691, n_952, n_1229, n_391, n_701, n_1437, n_1023, n_645, n_539, n_803, n_1092, n_238, n_1776, n_531, n_1757, n_890, n_1897, n_764, n_1919, n_1056, n_1424, n_162, n_960, n_1893, n_222, n_1290, n_1123, n_1467, n_1047, n_634, n_199, n_32, n_1252, n_348, n_1382, n_1029, n_925, n_1206, n_424, n_1311, n_1519, n_256, n_950, n_1553, n_1811, n_380, n_419, n_1346, n_444, n_1299, n_1808, n_1060, n_1141, n_316, n_389, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_451, n_619, n_408, n_1386, n_1699, n_376, n_967, n_1442, n_74, n_1139, n_515, n_57, n_351, n_885, n_397, n_1432, n_1357, n_483, n_683, n_1632, n_1057, n_1051, n_1085, n_1066, n_721, n_1157, n_841, n_1050, n_22, n_802, n_46, n_1608, n_983, n_1844, n_38, n_280, n_1305, n_873, n_1826, n_378, n_1112, n_762, n_1283, n_1644, n_17, n_690, n_33, n_583, n_302, n_1343, n_1203, n_1631, n_821, n_1763, n_1768, n_321, n_1179, n_621, n_753, n_455, n_1048, n_1719, n_1288, n_212, n_385, n_507, n_1560, n_1605, n_330, n_1228, n_972, n_692, n_820, n_1200, n_1911, n_1301, n_1363, n_1668, n_1185, n_991, n_828, n_779, n_576, n_1143, n_1579, n_1329, n_1312, n_1439, n_804, n_537, n_1688, n_945, n_492, n_153, n_1504, n_943, n_341, n_250, n_992, n_543, n_260, n_842, n_650, n_984, n_694, n_286, n_1643, n_883, n_470, n_325, n_449, n_1594, n_132, n_1214, n_1342, n_1400, n_900, n_856, n_1793, n_918, n_942, n_1804, n_189, n_1147, n_1557, n_1610, n_13, n_1077, n_1422, n_540, n_618, n_896, n_323, n_195, n_356, n_894, n_1636, n_1730, n_831, n_964, n_1373, n_1350, n_1511, n_1865, n_1470, n_1096, n_234, n_1575, n_1697, n_1735, n_833, n_5, n_1646, n_225, n_1307, n_1881, n_988, n_814, n_192, n_1549, n_1201, n_1114, n_655, n_1616, n_1446, n_669, n_472, n_1458, n_1176, n_1472, n_1807, n_387, n_1149, n_398, n_1671, n_635, n_763, n_1020, n_1062, n_211, n_1824, n_1917, n_1219, n_3, n_1204, n_178, n_1814, n_1035, n_287, n_555, n_783, n_1848, n_1188, n_1722, n_661, n_41, n_1802, n_849, n_15, n_336, n_584, n_681, n_1638, n_1786, n_50, n_430, n_510, n_216, n_311, n_830, n_1296, n_1413, n_801, n_241, n_875, n_357, n_1110, n_1655, n_445, n_749, n_1895, n_1134, n_1358, n_717, n_165, n_939, n_482, n_1088, n_588, n_1173, n_789, n_1232, n_1603, n_734, n_638, n_866, n_107, n_969, n_1401, n_1019, n_1105, n_249, n_304, n_1338, n_577, n_1522, n_1687, n_1637, n_1419, n_338, n_149, n_1653, n_693, n_1506, n_14, n_836, n_990, n_1886, n_1389, n_1894, n_975, n_1908, n_1256, n_1702, n_567, n_1465, n_778, n_1122, n_151, n_306, n_458, n_770, n_1375, n_1102, n_1843, n_711, n_1499, n_85, n_1187, n_1441, n_1392, n_1597, n_1164, n_1659, n_1834, n_489, n_1174, n_1371, n_617, n_1303, n_1572, n_876, n_1516, n_1190, n_1736, n_1685, n_118, n_601, n_917, n_1714, n_966, n_253, n_1116, n_1661, n_1212, n_1541, n_172, n_206, n_217, n_726, n_982, n_1573, n_1453, n_1731, n_818, n_861, n_1713, n_1183, n_1658, n_899, n_1253, n_210, n_1737, n_1904, n_774, n_1628, n_1335, n_1514, n_1777, n_1059, n_1345, n_176, n_1133, n_1771, n_1912, n_1899, n_557, n_1410, n_1005, n_607, n_1003, n_679, n_710, n_527, n_1168, n_707, n_937, n_1427, n_393, n_108, n_487, n_1584, n_665, n_1726, n_1835, n_66, n_1440, n_177, n_421, n_1853, n_1356, n_1787, n_910, n_1657, n_768, n_1475, n_1302, n_1774, n_1725, n_205, n_1136, n_1313, n_1491, n_754, n_1496, n_179, n_1125, n_125, n_410, n_708, n_529, n_1812, n_735, n_232, n_1915, n_1109, n_126, n_895, n_1310, n_1803, n_202, n_427, n_1399, n_1543, n_791, n_732, n_1533, n_193, n_808, n_797, n_1025, n_500, n_1067, n_1720, n_148, n_435, n_159, n_766, n_1457, n_541, n_538, n_1117, n_799, n_687, n_715, n_1742, n_1480, n_1482, n_1213, n_1266, n_536, n_872, n_594, n_200, n_1291, n_1297, n_1753, n_1782, n_1155, n_1418, n_89, n_1524, n_1689, n_1485, n_115, n_1011, n_1184, n_985, n_1855, n_869, n_810, n_416, n_827, n_401, n_1703, n_1352, n_626, n_1650, n_1144, n_1137, n_1570, n_1170, n_305, n_137, n_676, n_294, n_318, n_653, n_642, n_1602, n_194, n_855, n_1178, n_1461, n_850, n_684, n_124, n_268, n_664, n_503, n_235, n_1372, n_605, n_1273, n_1822, n_353, n_620, n_643, n_916, n_1081, n_493, n_1235, n_703, n_698, n_980, n_1115, n_1282, n_1318, n_1783, n_780, n_998, n_1454, n_467, n_1227, n_1531, n_840, n_1334, n_1907, n_501, n_823, n_245, n_725, n_1388, n_1417, n_1295, n_672, n_1898, n_581, n_382, n_554, n_1625, n_898, n_1762, n_1013, n_1452, n_718, n_265, n_1120, n_719, n_443, n_1791, n_198, n_1890, n_1747, n_714, n_1683, n_1817, n_909, n_1497, n_1530, n_997, n_932, n_612, n_1409, n_788, n_1326, n_119, n_1268, n_559, n_825, n_508, n_506, n_1320, n_1663, n_737, n_1718, n_986, n_509, n_1317, n_147, n_1518, n_1715, n_1281, n_67, n_1192, n_1024, n_1063, n_1889, n_209, n_1792, n_1564, n_1868, n_1613, n_733, n_1489, n_1922, n_1376, n_941, n_981, n_1569, n_68, n_867, n_186, n_134, n_587, n_63, n_792, n_756, n_1429, n_399, n_1238, n_548, n_812, n_298, n_518, n_505, n_1772, n_282, n_752, n_905, n_1476, n_1108, n_782, n_1100, n_1861, n_1395, n_862, n_1425, n_760, n_1901, n_1900, n_1620, n_381, n_220, n_390, n_1330, n_1867, n_31, n_481, n_1675, n_1727, n_1554, n_1745, n_769, n_42, n_1046, n_271, n_934, n_1618, n_826, n_1813, n_886, n_1221, n_654, n_1172, n_167, n_379, n_428, n_1341, n_570, n_1641, n_1361, n_1707, n_853, n_377, n_751, n_786, n_1083, n_1142, n_1129, n_392, n_158, n_704, n_787, n_1770, n_138, n_961, n_1756, n_771, n_276, n_95, n_1716, n_1225, n_1520, n_169, n_522, n_1287, n_1262, n_400, n_930, n_181, n_1873, n_1411, n_221, n_622, n_1577, n_1087, n_386, n_994, n_1701, n_848, n_1550, n_1498, n_1223, n_1272, n_104, n_682, n_1567, n_56, n_141, n_1247, n_922, n_816, n_1648, n_591, n_145, n_1536, n_1857, n_1344, n_313, n_631, n_479, n_1246, n_1339, n_1478, n_1797, n_432, n_1769, n_839, n_1210, n_1364, n_328, n_140, n_1250, n_369, n_1842, n_871, n_598, n_685, n_928, n_608, n_1367, n_78, n_1460, n_772, n_1555, n_499, n_1589, n_517, n_98, n_402, n_413, n_1086, n_796, n_1858, n_1619, n_236, n_1502, n_1469, n_1012, n_1, n_1396, n_1348, n_903, n_1525, n_1752, n_740, n_203, n_384, n_1404, n_80, n_1794, n_35, n_1315, n_277, n_1061, n_92, n_1910, n_333, n_1298, n_1652, n_462, n_1193, n_1676, n_1255, n_258, n_1113, n_29, n_79, n_1226, n_722, n_1277, n_188, n_844, n_201, n_471, n_852, n_1487, n_40, n_1864, n_1028, n_1601, n_781, n_474, n_542, n_463, n_1546, n_595, n_502, n_466, n_420, n_1337, n_1495, n_632, n_699, n_979, n_1515, n_1627, n_1245, n_846, n_1673, n_465, n_76, n_362, n_1321, n_170, n_27, n_161, n_273, n_585, n_1739, n_270, n_616, n_81, n_1914, n_745, n_1654, n_1103, n_648, n_1379, n_312, n_1076, n_1091, n_1408, n_494, n_1761, n_641, n_730, n_1325, n_1595, n_354, n_575, n_480, n_425, n_795, n_695, n_180, n_656, n_1606, n_1220, n_37, n_1694, n_1540, n_229, n_437, n_1642, n_60, n_403, n_453, n_1130, n_720, n_0, n_1918, n_1526, n_863, n_805, n_1604, n_1275, n_1764, n_113, n_712, n_246, n_1583, n_1042, n_1402, n_269, n_285, n_412, n_1493, n_657, n_644, n_1741, n_1160, n_1397, n_491, n_1258, n_1074, n_1621, n_251, n_160, n_566, n_565, n_1448, n_1507, n_1398, n_1879, n_597, n_1181, n_1505, n_1634, n_1196, n_651, n_1340, n_334, n_811, n_1558, n_807, n_835, n_175, n_666, n_262, n_1433, n_1704, n_99, n_1254, n_1026, n_1234, n_319, n_364, n_1138, n_927, n_20, n_1089, n_1004, n_1186, n_1032, n_242, n_1681, n_1018, n_1693, n_438, n_713, n_904, n_1588, n_1622, n_166, n_1180, n_1827, n_1271, n_533, n_1542, n_1251, n_278, n_7687);

input n_924;
input n_1263;
input n_977;
input n_1378;
input n_611;
input n_1126;
input n_1423;
input n_1729;
input n_1166;
input n_1751;
input n_469;
input n_1508;
input n_82;
input n_785;
input n_549;
input n_532;
input n_1161;
input n_1859;
input n_1677;
input n_1150;
input n_226;
input n_1780;
input n_1488;
input n_667;
input n_790;
input n_1055;
input n_1501;
input n_111;
input n_880;
input n_544;
input n_1007;
input n_155;
input n_552;
input n_1528;
input n_1370;
input n_1292;
input n_1198;
input n_1360;
input n_1099;
input n_956;
input n_564;
input n_423;
input n_1738;
input n_21;
input n_105;
input n_1021;
input n_4;
input n_551;
input n_1323;
input n_1466;
input n_688;
input n_1695;
input n_1353;
input n_800;
input n_1347;
input n_1535;
input n_1789;
input n_1666;
input n_671;
input n_819;
input n_1451;
input n_1022;
input n_915;
input n_1545;
input n_864;
input n_173;
input n_859;
input n_951;
input n_1264;
input n_447;
input n_247;
input n_1494;
input n_292;
input n_625;
input n_854;
input n_1462;
input n_1799;
input n_1580;
input n_674;
input n_417;
input n_1806;
input n_516;
input n_933;
input n_1152;
input n_497;
input n_1869;
input n_1607;
input n_1563;
input n_606;
input n_275;
input n_26;
input n_877;
input n_2;
input n_1696;
input n_755;
input n_1118;
input n_6;
input n_1686;
input n_947;
input n_1285;
input n_373;
input n_307;
input n_1860;
input n_1359;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_1728;
input n_556;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_1896;
input n_929;
input n_1124;
input n_1818;
input n_902;
input n_1576;
input n_191;
input n_1104;
input n_1294;
input n_659;
input n_51;
input n_1705;
input n_1257;
input n_171;
input n_1182;
input n_579;
input n_1698;
input n_1261;
input n_938;
input n_1098;
input n_320;
input n_1154;
input n_1242;
input n_1135;
input n_24;
input n_406;
input n_519;
input n_1016;
input n_1243;
input n_546;
input n_101;
input n_1280;
input n_1845;
input n_281;
input n_240;
input n_291;
input n_231;
input n_257;
input n_731;
input n_371;
input n_1483;
input n_1314;
input n_1512;
input n_709;
input n_1490;
input n_317;
input n_1236;
input n_1633;
input n_569;
input n_1778;
input n_227;
input n_920;
input n_1289;
input n_1517;
input n_94;
input n_335;
input n_1669;
input n_370;
input n_976;
input n_343;
input n_1449;
input n_308;
input n_1566;
input n_297;
input n_156;
input n_1078;
input n_1670;
input n_775;
input n_219;
input n_157;
input n_600;
input n_1484;
input n_1374;
input n_1328;
input n_223;
input n_264;
input n_1877;
input n_1831;
input n_1598;
input n_1723;
input n_955;
input n_1850;
input n_163;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_1036;
input n_1097;
input n_1749;
input n_347;
input n_59;
input n_550;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_646;
input n_1428;
input n_436;
input n_1394;
input n_1414;
input n_1216;
input n_290;
input n_580;
input n_1040;
input n_1872;
input n_1852;
input n_578;
input n_926;
input n_344;
input n_1218;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1547;
input n_1030;
input n_72;
input n_1755;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_1267;
input n_1561;
input n_496;
input n_1801;
input n_1391;
input n_958;
input n_1034;
input n_670;
input n_1513;
input n_1600;
input n_48;
input n_521;
input n_663;
input n_845;
input n_1862;
input n_673;
input n_837;
input n_1239;
input n_528;
input n_1796;
input n_680;
input n_1473;
input n_1587;
input n_395;
input n_164;
input n_553;
input n_901;
input n_813;
input n_1521;
input n_1284;
input n_1590;
input n_214;
input n_1748;
input n_1672;
input n_675;
input n_888;
input n_1880;
input n_1167;
input n_1626;
input n_637;
input n_1384;
input n_1556;
input n_184;
input n_446;
input n_1863;
input n_1064;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_691;
input n_1151;
input n_881;
input n_1405;
input n_1706;
input n_468;
input n_213;
input n_129;
input n_342;
input n_464;
input n_363;
input n_1582;
input n_197;
input n_1069;
input n_1784;
input n_1075;
input n_1836;
input n_1450;
input n_1322;
input n_1471;
input n_1750;
input n_1459;
input n_460;
input n_889;
input n_973;
input n_1700;
input n_477;
input n_571;
input n_1585;
input n_461;
input n_1599;
input n_1211;
input n_1197;
input n_1523;
input n_907;
input n_1447;
input n_1377;
input n_190;
input n_989;
input n_1039;
input n_34;
input n_228;
input n_283;
input n_1403;
input n_488;
input n_736;
input n_892;
input n_1000;
input n_1202;
input n_1278;
input n_1002;
input n_1463;
input n_1581;
input n_49;
input n_310;
input n_54;
input n_593;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_1667;
input n_838;
input n_332;
input n_1053;
input n_1224;
input n_349;
input n_1248;
input n_230;
input n_1331;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_1385;
input n_440;
input n_793;
input n_478;
input n_1819;
input n_476;
input n_1527;
input n_534;
input n_1882;
input n_884;
input n_345;
input n_944;
input n_1754;
input n_1623;
input n_1854;
input n_91;
input n_1565;
input n_1809;
input n_1856;
input n_182;
input n_143;
input n_647;
input n_237;
input n_407;
input n_1072;
input n_832;
input n_857;
input n_207;
input n_561;
input n_1319;
input n_1825;
input n_1883;
input n_1906;
input n_1712;
input n_1387;
input n_1532;
input n_18;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_686;
input n_847;
input n_1393;
input n_596;
input n_1775;
input n_1368;
input n_558;
input n_702;
input n_1276;
input n_822;
input n_1412;
input n_1709;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1538;
input n_1838;
input n_1199;
input n_1847;
input n_1779;
input n_352;
input n_1884;
input n_53;
input n_1038;
input n_520;
input n_1369;
input n_409;
input n_1841;
input n_1660;
input n_887;
input n_1905;
input n_154;
input n_71;
input n_300;
input n_809;
input n_870;
input n_931;
input n_599;
input n_1711;
input n_1662;
input n_1891;
input n_1481;
input n_434;
input n_1544;
input n_868;
input n_639;
input n_914;
input n_411;
input n_414;
input n_1629;
input n_1293;
input n_965;
input n_1876;
input n_1743;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_360;
input n_36;
input n_1479;
input n_1810;
input n_64;
input n_1888;
input n_759;
input n_1892;
input n_28;
input n_806;
input n_1766;
input n_1477;
input n_324;
input n_1635;
input n_1571;
input n_187;
input n_1189;
input n_103;
input n_97;
input n_11;
input n_7;
input n_1259;
input n_1690;
input n_706;
input n_746;
input n_1649;
input n_747;
input n_52;
input n_784;
input n_110;
input n_1733;
input n_1244;
input n_431;
input n_1194;
input n_1815;
input n_615;
input n_851;
input n_1759;
input n_843;
input n_1788;
input n_523;
input n_913;
input n_1537;
input n_705;
input n_865;
input n_61;
input n_678;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_1679;
input n_776;
input n_1798;
input n_1790;
input n_1415;
input n_367;
input n_452;
input n_525;
input n_1260;
input n_1746;
input n_1647;
input n_1829;
input n_1464;
input n_649;
input n_547;
input n_43;
input n_1444;
input n_1191;
input n_1674;
input n_1833;
input n_116;
input n_1830;
input n_1710;
input n_284;
input n_1128;
input n_139;
input n_1734;
input n_744;
input n_590;
input n_629;
input n_1308;
input n_1767;
input n_254;
input n_1680;
input n_1233;
input n_23;
input n_1615;
input n_1529;
input n_526;
input n_1916;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1333;
input n_1121;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_949;
input n_100;
input n_1443;
input n_1008;
input n_946;
input n_1539;
input n_1001;
input n_1503;
input n_498;
input n_1468;
input n_1559;
input n_1765;
input n_1866;
input n_689;
input n_738;
input n_1624;
input n_640;
input n_1510;
input n_252;
input n_624;
input n_1380;
input n_1744;
input n_1617;
input n_295;
input n_133;
input n_1010;
input n_1231;
input n_739;
input n_1279;
input n_1406;
input n_1195;
input n_1837;
input n_1839;
input n_610;
input n_1760;
input n_936;
input n_568;
input n_1500;
input n_39;
input n_1090;
input n_757;
input n_633;
input n_439;
input n_106;
input n_1832;
input n_259;
input n_448;
input n_1851;
input n_758;
input n_999;
input n_93;
input n_1656;
input n_1158;
input n_1509;
input n_1874;
input n_563;
input n_1145;
input n_878;
input n_524;
input n_204;
input n_394;
input n_1678;
input n_1049;
input n_1153;
input n_741;
input n_1639;
input n_1306;
input n_1068;
input n_1871;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_1207;
input n_919;
input n_908;
input n_90;
input n_724;
input n_1781;
input n_658;
input n_1740;
input n_1362;
input n_1586;
input n_456;
input n_959;
input n_535;
input n_152;
input n_940;
input n_1445;
input n_9;
input n_1492;
input n_1923;
input n_1773;
input n_592;
input n_1169;
input n_45;
input n_1596;
input n_1692;
input n_1017;
input n_123;
input n_978;
input n_1434;
input n_1054;
input n_1474;
input n_1665;
input n_1269;
input n_1095;
input n_1828;
input n_1614;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_603;
input n_1431;
input n_484;
input n_1593;
input n_1033;
input n_442;
input n_131;
input n_636;
input n_660;
input n_1640;
input n_1732;
input n_1009;
input n_1148;
input n_109;
input n_742;
input n_750;
input n_995;
input n_454;
input n_1609;
input n_374;
input n_185;
input n_396;
input n_1887;
input n_1383;
input n_1073;
input n_255;
input n_662;
input n_459;
input n_218;
input n_962;
input n_1215;
input n_1171;
input n_1578;
input n_723;
input n_1920;
input n_1065;
input n_1592;
input n_1336;
input n_1721;
input n_1758;
input n_1574;
input n_473;
input n_1921;
input n_1309;
input n_1878;
input n_1426;
input n_1043;
input n_355;
input n_486;
input n_1800;
input n_1548;
input n_614;
input n_337;
input n_1421;
input n_88;
input n_1286;
input n_1177;
input n_1355;
input n_168;
input n_974;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_743;
input n_299;
input n_303;
input n_296;
input n_613;
input n_1119;
input n_1240;
input n_1820;
input n_65;
input n_829;
input n_1612;
input n_1416;
input n_1724;
input n_361;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1420;
input n_1132;
input n_388;
input n_1366;
input n_1300;
input n_1127;
input n_761;
input n_1785;
input n_1568;
input n_1006;
input n_329;
input n_274;
input n_1270;
input n_1664;
input n_1486;
input n_582;
input n_1332;
input n_1390;
input n_73;
input n_19;
input n_1870;
input n_309;
input n_30;
input n_512;
input n_1591;
input n_84;
input n_130;
input n_322;
input n_1682;
input n_1249;
input n_652;
input n_1111;
input n_1365;
input n_25;
input n_1349;
input n_1093;
input n_288;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_1265;
input n_1909;
input n_44;
input n_224;
input n_1562;
input n_383;
input n_834;
input n_112;
input n_765;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_1651;
input n_239;
input n_630;
input n_1902;
input n_55;
input n_1913;
input n_504;
input n_1823;
input n_511;
input n_874;
input n_358;
input n_1101;
input n_77;
input n_102;
input n_1106;
input n_1456;
input n_1875;
input n_1304;
input n_1324;
input n_987;
input n_1846;
input n_261;
input n_174;
input n_1885;
input n_1455;
input n_767;
input n_993;
input n_1903;
input n_1407;
input n_1551;
input n_545;
input n_441;
input n_860;
input n_450;
input n_1805;
input n_1816;
input n_429;
input n_948;
input n_1217;
input n_628;
input n_365;
input n_1849;
input n_729;
input n_1131;
input n_1084;
input n_970;
input n_911;
input n_1430;
input n_83;
input n_513;
input n_1094;
input n_1354;
input n_560;
input n_1534;
input n_340;
input n_1351;
input n_1044;
input n_1205;
input n_346;
input n_1209;
input n_1552;
input n_495;
input n_602;
input n_574;
input n_1435;
input n_879;
input n_16;
input n_58;
input n_623;
input n_405;
input n_824;
input n_359;
input n_1645;
input n_490;
input n_1327;
input n_996;
input n_921;
input n_1684;
input n_233;
input n_1717;
input n_572;
input n_366;
input n_815;
input n_1795;
input n_128;
input n_1821;
input n_120;
input n_327;
input n_135;
input n_1381;
input n_1611;
input n_1037;
input n_1080;
input n_1274;
input n_1316;
input n_1708;
input n_426;
input n_1438;
input n_1082;
input n_1840;
input n_589;
input n_716;
input n_1630;
input n_562;
input n_1436;
input n_62;
input n_1691;
input n_952;
input n_1229;
input n_391;
input n_701;
input n_1437;
input n_1023;
input n_645;
input n_539;
input n_803;
input n_1092;
input n_238;
input n_1776;
input n_531;
input n_1757;
input n_890;
input n_1897;
input n_764;
input n_1919;
input n_1056;
input n_1424;
input n_162;
input n_960;
input n_1893;
input n_222;
input n_1290;
input n_1123;
input n_1467;
input n_1047;
input n_634;
input n_199;
input n_32;
input n_1252;
input n_348;
input n_1382;
input n_1029;
input n_925;
input n_1206;
input n_424;
input n_1311;
input n_1519;
input n_256;
input n_950;
input n_1553;
input n_1811;
input n_380;
input n_419;
input n_1346;
input n_444;
input n_1299;
input n_1808;
input n_1060;
input n_1141;
input n_316;
input n_389;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_451;
input n_619;
input n_408;
input n_1386;
input n_1699;
input n_376;
input n_967;
input n_1442;
input n_74;
input n_1139;
input n_515;
input n_57;
input n_351;
input n_885;
input n_397;
input n_1432;
input n_1357;
input n_483;
input n_683;
input n_1632;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_1157;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_46;
input n_1608;
input n_983;
input n_1844;
input n_38;
input n_280;
input n_1305;
input n_873;
input n_1826;
input n_378;
input n_1112;
input n_762;
input n_1283;
input n_1644;
input n_17;
input n_690;
input n_33;
input n_583;
input n_302;
input n_1343;
input n_1203;
input n_1631;
input n_821;
input n_1763;
input n_1768;
input n_321;
input n_1179;
input n_621;
input n_753;
input n_455;
input n_1048;
input n_1719;
input n_1288;
input n_212;
input n_385;
input n_507;
input n_1560;
input n_1605;
input n_330;
input n_1228;
input n_972;
input n_692;
input n_820;
input n_1200;
input n_1911;
input n_1301;
input n_1363;
input n_1668;
input n_1185;
input n_991;
input n_828;
input n_779;
input n_576;
input n_1143;
input n_1579;
input n_1329;
input n_1312;
input n_1439;
input n_804;
input n_537;
input n_1688;
input n_945;
input n_492;
input n_153;
input n_1504;
input n_943;
input n_341;
input n_250;
input n_992;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_286;
input n_1643;
input n_883;
input n_470;
input n_325;
input n_449;
input n_1594;
input n_132;
input n_1214;
input n_1342;
input n_1400;
input n_900;
input n_856;
input n_1793;
input n_918;
input n_942;
input n_1804;
input n_189;
input n_1147;
input n_1557;
input n_1610;
input n_13;
input n_1077;
input n_1422;
input n_540;
input n_618;
input n_896;
input n_323;
input n_195;
input n_356;
input n_894;
input n_1636;
input n_1730;
input n_831;
input n_964;
input n_1373;
input n_1350;
input n_1511;
input n_1865;
input n_1470;
input n_1096;
input n_234;
input n_1575;
input n_1697;
input n_1735;
input n_833;
input n_5;
input n_1646;
input n_225;
input n_1307;
input n_1881;
input n_988;
input n_814;
input n_192;
input n_1549;
input n_1201;
input n_1114;
input n_655;
input n_1616;
input n_1446;
input n_669;
input n_472;
input n_1458;
input n_1176;
input n_1472;
input n_1807;
input n_387;
input n_1149;
input n_398;
input n_1671;
input n_635;
input n_763;
input n_1020;
input n_1062;
input n_211;
input n_1824;
input n_1917;
input n_1219;
input n_3;
input n_1204;
input n_178;
input n_1814;
input n_1035;
input n_287;
input n_555;
input n_783;
input n_1848;
input n_1188;
input n_1722;
input n_661;
input n_41;
input n_1802;
input n_849;
input n_15;
input n_336;
input n_584;
input n_681;
input n_1638;
input n_1786;
input n_50;
input n_430;
input n_510;
input n_216;
input n_311;
input n_830;
input n_1296;
input n_1413;
input n_801;
input n_241;
input n_875;
input n_357;
input n_1110;
input n_1655;
input n_445;
input n_749;
input n_1895;
input n_1134;
input n_1358;
input n_717;
input n_165;
input n_939;
input n_482;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_1232;
input n_1603;
input n_734;
input n_638;
input n_866;
input n_107;
input n_969;
input n_1401;
input n_1019;
input n_1105;
input n_249;
input n_304;
input n_1338;
input n_577;
input n_1522;
input n_1687;
input n_1637;
input n_1419;
input n_338;
input n_149;
input n_1653;
input n_693;
input n_1506;
input n_14;
input n_836;
input n_990;
input n_1886;
input n_1389;
input n_1894;
input n_975;
input n_1908;
input n_1256;
input n_1702;
input n_567;
input n_1465;
input n_778;
input n_1122;
input n_151;
input n_306;
input n_458;
input n_770;
input n_1375;
input n_1102;
input n_1843;
input n_711;
input n_1499;
input n_85;
input n_1187;
input n_1441;
input n_1392;
input n_1597;
input n_1164;
input n_1659;
input n_1834;
input n_489;
input n_1174;
input n_1371;
input n_617;
input n_1303;
input n_1572;
input n_876;
input n_1516;
input n_1190;
input n_1736;
input n_1685;
input n_118;
input n_601;
input n_917;
input n_1714;
input n_966;
input n_253;
input n_1116;
input n_1661;
input n_1212;
input n_1541;
input n_172;
input n_206;
input n_217;
input n_726;
input n_982;
input n_1573;
input n_1453;
input n_1731;
input n_818;
input n_861;
input n_1713;
input n_1183;
input n_1658;
input n_899;
input n_1253;
input n_210;
input n_1737;
input n_1904;
input n_774;
input n_1628;
input n_1335;
input n_1514;
input n_1777;
input n_1059;
input n_1345;
input n_176;
input n_1133;
input n_1771;
input n_1912;
input n_1899;
input n_557;
input n_1410;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_527;
input n_1168;
input n_707;
input n_937;
input n_1427;
input n_393;
input n_108;
input n_487;
input n_1584;
input n_665;
input n_1726;
input n_1835;
input n_66;
input n_1440;
input n_177;
input n_421;
input n_1853;
input n_1356;
input n_1787;
input n_910;
input n_1657;
input n_768;
input n_1475;
input n_1302;
input n_1774;
input n_1725;
input n_205;
input n_1136;
input n_1313;
input n_1491;
input n_754;
input n_1496;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_708;
input n_529;
input n_1812;
input n_735;
input n_232;
input n_1915;
input n_1109;
input n_126;
input n_895;
input n_1310;
input n_1803;
input n_202;
input n_427;
input n_1399;
input n_1543;
input n_791;
input n_732;
input n_1533;
input n_193;
input n_808;
input n_797;
input n_1025;
input n_500;
input n_1067;
input n_1720;
input n_148;
input n_435;
input n_159;
input n_766;
input n_1457;
input n_541;
input n_538;
input n_1117;
input n_799;
input n_687;
input n_715;
input n_1742;
input n_1480;
input n_1482;
input n_1213;
input n_1266;
input n_536;
input n_872;
input n_594;
input n_200;
input n_1291;
input n_1297;
input n_1753;
input n_1782;
input n_1155;
input n_1418;
input n_89;
input n_1524;
input n_1689;
input n_1485;
input n_115;
input n_1011;
input n_1184;
input n_985;
input n_1855;
input n_869;
input n_810;
input n_416;
input n_827;
input n_401;
input n_1703;
input n_1352;
input n_626;
input n_1650;
input n_1144;
input n_1137;
input n_1570;
input n_1170;
input n_305;
input n_137;
input n_676;
input n_294;
input n_318;
input n_653;
input n_642;
input n_1602;
input n_194;
input n_855;
input n_1178;
input n_1461;
input n_850;
input n_684;
input n_124;
input n_268;
input n_664;
input n_503;
input n_235;
input n_1372;
input n_605;
input n_1273;
input n_1822;
input n_353;
input n_620;
input n_643;
input n_916;
input n_1081;
input n_493;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_1282;
input n_1318;
input n_1783;
input n_780;
input n_998;
input n_1454;
input n_467;
input n_1227;
input n_1531;
input n_840;
input n_1334;
input n_1907;
input n_501;
input n_823;
input n_245;
input n_725;
input n_1388;
input n_1417;
input n_1295;
input n_672;
input n_1898;
input n_581;
input n_382;
input n_554;
input n_1625;
input n_898;
input n_1762;
input n_1013;
input n_1452;
input n_718;
input n_265;
input n_1120;
input n_719;
input n_443;
input n_1791;
input n_198;
input n_1890;
input n_1747;
input n_714;
input n_1683;
input n_1817;
input n_909;
input n_1497;
input n_1530;
input n_997;
input n_932;
input n_612;
input n_1409;
input n_788;
input n_1326;
input n_119;
input n_1268;
input n_559;
input n_825;
input n_508;
input n_506;
input n_1320;
input n_1663;
input n_737;
input n_1718;
input n_986;
input n_509;
input n_1317;
input n_147;
input n_1518;
input n_1715;
input n_1281;
input n_67;
input n_1192;
input n_1024;
input n_1063;
input n_1889;
input n_209;
input n_1792;
input n_1564;
input n_1868;
input n_1613;
input n_733;
input n_1489;
input n_1922;
input n_1376;
input n_941;
input n_981;
input n_1569;
input n_68;
input n_867;
input n_186;
input n_134;
input n_587;
input n_63;
input n_792;
input n_756;
input n_1429;
input n_399;
input n_1238;
input n_548;
input n_812;
input n_298;
input n_518;
input n_505;
input n_1772;
input n_282;
input n_752;
input n_905;
input n_1476;
input n_1108;
input n_782;
input n_1100;
input n_1861;
input n_1395;
input n_862;
input n_1425;
input n_760;
input n_1901;
input n_1900;
input n_1620;
input n_381;
input n_220;
input n_390;
input n_1330;
input n_1867;
input n_31;
input n_481;
input n_1675;
input n_1727;
input n_1554;
input n_1745;
input n_769;
input n_42;
input n_1046;
input n_271;
input n_934;
input n_1618;
input n_826;
input n_1813;
input n_886;
input n_1221;
input n_654;
input n_1172;
input n_167;
input n_379;
input n_428;
input n_1341;
input n_570;
input n_1641;
input n_1361;
input n_1707;
input n_853;
input n_377;
input n_751;
input n_786;
input n_1083;
input n_1142;
input n_1129;
input n_392;
input n_158;
input n_704;
input n_787;
input n_1770;
input n_138;
input n_961;
input n_1756;
input n_771;
input n_276;
input n_95;
input n_1716;
input n_1225;
input n_1520;
input n_169;
input n_522;
input n_1287;
input n_1262;
input n_400;
input n_930;
input n_181;
input n_1873;
input n_1411;
input n_221;
input n_622;
input n_1577;
input n_1087;
input n_386;
input n_994;
input n_1701;
input n_848;
input n_1550;
input n_1498;
input n_1223;
input n_1272;
input n_104;
input n_682;
input n_1567;
input n_56;
input n_141;
input n_1247;
input n_922;
input n_816;
input n_1648;
input n_591;
input n_145;
input n_1536;
input n_1857;
input n_1344;
input n_313;
input n_631;
input n_479;
input n_1246;
input n_1339;
input n_1478;
input n_1797;
input n_432;
input n_1769;
input n_839;
input n_1210;
input n_1364;
input n_328;
input n_140;
input n_1250;
input n_369;
input n_1842;
input n_871;
input n_598;
input n_685;
input n_928;
input n_608;
input n_1367;
input n_78;
input n_1460;
input n_772;
input n_1555;
input n_499;
input n_1589;
input n_517;
input n_98;
input n_402;
input n_413;
input n_1086;
input n_796;
input n_1858;
input n_1619;
input n_236;
input n_1502;
input n_1469;
input n_1012;
input n_1;
input n_1396;
input n_1348;
input n_903;
input n_1525;
input n_1752;
input n_740;
input n_203;
input n_384;
input n_1404;
input n_80;
input n_1794;
input n_35;
input n_1315;
input n_277;
input n_1061;
input n_92;
input n_1910;
input n_333;
input n_1298;
input n_1652;
input n_462;
input n_1193;
input n_1676;
input n_1255;
input n_258;
input n_1113;
input n_29;
input n_79;
input n_1226;
input n_722;
input n_1277;
input n_188;
input n_844;
input n_201;
input n_471;
input n_852;
input n_1487;
input n_40;
input n_1864;
input n_1028;
input n_1601;
input n_781;
input n_474;
input n_542;
input n_463;
input n_1546;
input n_595;
input n_502;
input n_466;
input n_420;
input n_1337;
input n_1495;
input n_632;
input n_699;
input n_979;
input n_1515;
input n_1627;
input n_1245;
input n_846;
input n_1673;
input n_465;
input n_76;
input n_362;
input n_1321;
input n_170;
input n_27;
input n_161;
input n_273;
input n_585;
input n_1739;
input n_270;
input n_616;
input n_81;
input n_1914;
input n_745;
input n_1654;
input n_1103;
input n_648;
input n_1379;
input n_312;
input n_1076;
input n_1091;
input n_1408;
input n_494;
input n_1761;
input n_641;
input n_730;
input n_1325;
input n_1595;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_695;
input n_180;
input n_656;
input n_1606;
input n_1220;
input n_37;
input n_1694;
input n_1540;
input n_229;
input n_437;
input n_1642;
input n_60;
input n_403;
input n_453;
input n_1130;
input n_720;
input n_0;
input n_1918;
input n_1526;
input n_863;
input n_805;
input n_1604;
input n_1275;
input n_1764;
input n_113;
input n_712;
input n_246;
input n_1583;
input n_1042;
input n_1402;
input n_269;
input n_285;
input n_412;
input n_1493;
input n_657;
input n_644;
input n_1741;
input n_1160;
input n_1397;
input n_491;
input n_1258;
input n_1074;
input n_1621;
input n_251;
input n_160;
input n_566;
input n_565;
input n_1448;
input n_1507;
input n_1398;
input n_1879;
input n_597;
input n_1181;
input n_1505;
input n_1634;
input n_1196;
input n_651;
input n_1340;
input n_334;
input n_811;
input n_1558;
input n_807;
input n_835;
input n_175;
input n_666;
input n_262;
input n_1433;
input n_1704;
input n_99;
input n_1254;
input n_1026;
input n_1234;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_1681;
input n_1018;
input n_1693;
input n_438;
input n_713;
input n_904;
input n_1588;
input n_1622;
input n_166;
input n_1180;
input n_1827;
input n_1271;
input n_533;
input n_1542;
input n_1251;
input n_278;

output n_7687;

wire n_6643;
wire n_6122;
wire n_2417;
wire n_2253;
wire n_2756;
wire n_4706;
wire n_5567;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_6579;
wire n_7164;
wire n_5287;
wire n_6546;
wire n_2327;
wire n_2899;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_5978;
wire n_2395;
wire n_5161;
wire n_5776;
wire n_6551;
wire n_5512;
wire n_5207;
wire n_2347;
wire n_6786;
wire n_7206;
wire n_7303;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_7461;
wire n_2487;
wire n_6649;
wire n_7154;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_6810;
wire n_7660;
wire n_6276;
wire n_6072;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_7686;
wire n_4211;
wire n_7024;
wire n_3448;
wire n_7205;
wire n_6742;
wire n_3019;
wire n_2096;
wire n_6694;
wire n_3776;
wire n_7616;
wire n_2530;
wire n_4517;
wire n_2483;
wire n_7486;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_4615;
wire n_2076;
wire n_6090;
wire n_6580;
wire n_7010;
wire n_5480;
wire n_6549;
wire n_6913;
wire n_2147;
wire n_3010;
wire n_7315;
wire n_7004;
wire n_2770;
wire n_4131;
wire n_5402;
wire n_2584;
wire n_5851;
wire n_3188;
wire n_5509;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_7641;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_3283;
wire n_7468;
wire n_5469;
wire n_2323;
wire n_6431;
wire n_5744;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_5202;
wire n_5648;
wire n_7667;
wire n_6931;
wire n_6618;
wire n_6408;
wire n_3214;
wire n_7523;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_5922;
wire n_6698;
wire n_4678;
wire n_2032;
wire n_2587;
wire n_5848;
wire n_5406;
wire n_6085;
wire n_3947;
wire n_3490;
wire n_7421;
wire n_7306;
wire n_6214;
wire n_7493;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_6939;
wire n_2384;
wire n_7528;
wire n_3156;
wire n_3376;
wire n_7562;
wire n_5037;
wire n_4468;
wire n_5661;
wire n_6991;
wire n_3653;
wire n_5562;
wire n_3702;
wire n_4976;
wire n_6586;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_6096;
wire n_2276;
wire n_6707;
wire n_5852;
wire n_2089;
wire n_3420;
wire n_6920;
wire n_6868;
wire n_5144;
wire n_3361;
wire n_4758;
wire n_7402;
wire n_4255;
wire n_5577;
wire n_4484;
wire n_7592;
wire n_3668;
wire n_7152;
wire n_6512;
wire n_4237;
wire n_2934;
wire n_3550;
wire n_5689;
wire n_5894;
wire n_2079;
wire n_2238;
wire n_7463;
wire n_3418;
wire n_4901;
wire n_6725;
wire n_7613;
wire n_2859;
wire n_3395;
wire n_7083;
wire n_4917;
wire n_7086;
wire n_7349;
wire n_6464;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_7647;
wire n_5825;
wire n_2968;
wire n_7316;
wire n_6820;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_4421;
wire n_6098;
wire n_7019;
wire n_6686;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_4469;
wire n_4414;
wire n_6561;
wire n_6584;
wire n_7452;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3735;
wire n_3349;
wire n_7323;
wire n_2248;
wire n_7195;
wire n_6701;
wire n_7478;
wire n_3007;
wire n_6769;
wire n_7683;
wire n_6592;
wire n_5686;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_6062;
wire n_6191;
wire n_2258;
wire n_3983;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_4195;
wire n_4969;
wire n_4504;
wire n_5909;
wire n_7575;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_4531;
wire n_6043;
wire n_2987;
wire n_6271;
wire n_7171;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_6793;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_7127;
wire n_5397;
wire n_4471;
wire n_6550;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_5709;
wire n_7568;
wire n_3208;
wire n_6021;
wire n_3331;
wire n_4983;
wire n_2379;
wire n_5695;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_5860;
wire n_6926;
wire n_3649;
wire n_4302;
wire n_7589;
wire n_6928;
wire n_2514;
wire n_5862;
wire n_6304;
wire n_5189;
wire n_6956;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_7026;
wire n_4160;
wire n_6782;
wire n_2293;
wire n_5854;
wire n_5516;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_7002;
wire n_3981;
wire n_7141;
wire n_5936;
wire n_6126;
wire n_6027;
wire n_6598;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_6342;
wire n_6638;
wire n_7308;
wire n_5254;
wire n_3526;
wire n_6900;
wire n_2546;
wire n_3790;
wire n_7264;
wire n_3491;
wire n_7457;
wire n_4613;
wire n_4649;
wire n_7617;
wire n_6269;
wire n_5615;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_5902;
wire n_4028;
wire n_5479;
wire n_3819;
wire n_6013;
wire n_7357;
wire n_2449;
wire n_5083;
wire n_6927;
wire n_6503;
wire n_5888;
wire n_2297;
wire n_4186;
wire n_7310;
wire n_4731;
wire n_2177;
wire n_3747;
wire n_5698;
wire n_5592;
wire n_7521;
wire n_2227;
wire n_4618;
wire n_3346;
wire n_2190;
wire n_4742;
wire n_7593;
wire n_6256;
wire n_2876;
wire n_4099;
wire n_7406;
wire n_7600;
wire n_3484;
wire n_3620;
wire n_2479;
wire n_5870;
wire n_4295;
wire n_5303;
wire n_7076;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_6982;
wire n_4697;
wire n_7286;
wire n_7137;
wire n_4190;
wire n_3994;
wire n_2607;
wire n_4810;
wire n_6727;
wire n_3317;
wire n_7539;
wire n_7229;
wire n_4391;
wire n_5954;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_4638;
wire n_3455;
wire n_6097;
wire n_5047;
wire n_3452;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_7125;
wire n_6677;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_6624;
wire n_7121;
wire n_2796;
wire n_6466;
wire n_2342;
wire n_4156;
wire n_4848;
wire n_2937;
wire n_6008;
wire n_3095;
wire n_2805;
wire n_5624;
wire n_4918;
wire n_5714;
wire n_5806;
wire n_3856;
wire n_7624;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_6221;
wire n_7160;
wire n_4002;
wire n_6805;
wire n_6185;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_6568;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_6004;
wire n_6351;
wire n_7552;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_6901;
wire n_2947;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_4801;
wire n_7183;
wire n_6411;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_3287;
wire n_3378;
wire n_5435;
wire n_6873;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_5745;
wire n_7139;
wire n_4294;
wire n_5279;
wire n_4232;
wire n_4125;
wire n_4949;
wire n_2941;
wire n_6594;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_2536;
wire n_6387;
wire n_7223;
wire n_2952;
wire n_4847;
wire n_6179;
wire n_7338;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_6019;
wire n_6222;
wire n_7165;
wire n_3505;
wire n_6223;
wire n_4610;
wire n_6435;
wire n_3730;
wire n_4489;
wire n_7235;
wire n_5210;
wire n_6976;
wire n_4967;
wire n_6486;
wire n_5657;
wire n_6889;
wire n_6083;
wire n_4992;
wire n_6844;
wire n_3001;
wire n_7404;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_6295;
wire n_3597;
wire n_4198;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_5857;
wire n_4534;
wire n_4500;
wire n_7437;
wire n_5014;
wire n_6241;
wire n_3185;
wire n_6087;
wire n_3523;
wire n_2829;
wire n_4597;
wire n_6846;
wire n_4329;
wire n_4087;
wire n_3811;
wire n_3200;
wire n_5756;
wire n_2231;
wire n_6041;
wire n_2017;
wire n_2604;
wire n_6994;
wire n_4257;
wire n_3453;
wire n_7449;
wire n_7329;
wire n_2390;
wire n_5708;
wire n_3213;
wire n_6790;
wire n_3077;
wire n_7194;
wire n_6273;
wire n_3474;
wire n_3984;
wire n_6807;
wire n_5927;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_5638;
wire n_7115;
wire n_4189;
wire n_5670;
wire n_2803;
wire n_3707;
wire n_5584;
wire n_3429;
wire n_3849;
wire n_3946;
wire n_5965;
wire n_3229;
wire n_4463;
wire n_4687;
wire n_5751;
wire n_5664;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_5641;
wire n_4037;
wire n_6218;
wire n_7281;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_6824;
wire n_6189;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_6993;
wire n_3683;
wire n_6037;
wire n_7245;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_5963;
wire n_5980;
wire n_4763;
wire n_3590;
wire n_5310;
wire n_4594;
wire n_6153;
wire n_3424;
wire n_5970;
wire n_6418;
wire n_6564;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_7192;
wire n_3171;
wire n_6671;
wire n_6591;
wire n_6266;
wire n_7161;
wire n_7580;
wire n_7153;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_6517;
wire n_3468;
wire n_2910;
wire n_7350;
wire n_5690;
wire n_2163;
wire n_6967;
wire n_5885;
wire n_2254;
wire n_6433;
wire n_3546;
wire n_7535;
wire n_6893;
wire n_2647;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_7178;
wire n_7480;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_7632;
wire n_3244;
wire n_6501;
wire n_6028;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_5362;
wire n_6709;
wire n_4355;
wire n_3494;
wire n_6798;
wire n_5702;
wire n_5050;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_3110;
wire n_3073;
wire n_4572;
wire n_5527;
wire n_6986;
wire n_5609;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_5266;
wire n_7471;
wire n_3178;
wire n_5355;
wire n_2334;
wire n_6745;
wire n_4521;
wire n_4488;
wire n_5977;
wire n_6811;
wire n_2289;
wire n_3051;
wire n_2783;
wire n_6209;
wire n_2263;
wire n_6875;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_6853;
wire n_4519;
wire n_5551;
wire n_7594;
wire n_3715;
wire n_7340;
wire n_6699;
wire n_6073;
wire n_5767;
wire n_6324;
wire n_3040;
wire n_1938;
wire n_5640;
wire n_2499;
wire n_3568;
wire n_5655;
wire n_5475;
wire n_3737;
wire n_6138;
wire n_7603;
wire n_1967;
wire n_3255;
wire n_5692;
wire n_4856;
wire n_7494;
wire n_2997;
wire n_5921;
wire n_4400;
wire n_5168;
wire n_3326;
wire n_6477;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_6159;
wire n_6283;
wire n_7396;
wire n_5322;
wire n_7116;
wire n_4352;
wire n_7519;
wire n_4441;
wire n_6943;
wire n_4761;
wire n_6827;
wire n_6173;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_6312;
wire n_2533;
wire n_2364;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_3601;
wire n_6997;
wire n_5418;
wire n_2973;
wire n_2094;
wire n_2393;
wire n_7664;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_6300;
wire n_2043;
wire n_2751;
wire n_6131;
wire n_4893;
wire n_5032;
wire n_1934;
wire n_6537;
wire n_5933;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_4406;
wire n_2758;
wire n_7023;
wire n_2618;
wire n_7428;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_6783;
wire n_4748;
wire n_7465;
wire n_2295;
wire n_3931;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_2441;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_7149;
wire n_2795;
wire n_6459;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_5644;
wire n_2098;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_6869;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_3198;
wire n_2641;
wire n_4728;
wire n_7117;
wire n_4247;
wire n_4933;
wire n_6977;
wire n_4018;
wire n_3900;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_6313;
wire n_3872;
wire n_4336;
wire n_6569;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_2496;
wire n_2259;
wire n_6555;
wire n_3877;
wire n_6639;
wire n_7516;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_7596;
wire n_4052;
wire n_5864;
wire n_6536;
wire n_3459;
wire n_4398;
wire n_3155;
wire n_6490;
wire n_2633;
wire n_6961;
wire n_4954;
wire n_2435;
wire n_2097;
wire n_5460;
wire n_7628;
wire n_4304;
wire n_6761;
wire n_3911;
wire n_5333;
wire n_6294;
wire n_6767;
wire n_4431;
wire n_7427;
wire n_4192;
wire n_6802;
wire n_7527;
wire n_5570;
wire n_3736;
wire n_6326;
wire n_4805;
wire n_4885;
wire n_5983;
wire n_5804;
wire n_6376;
wire n_3565;
wire n_6167;
wire n_4701;
wire n_2575;
wire n_5910;
wire n_7411;
wire n_7101;
wire n_5040;
wire n_6730;
wire n_6948;
wire n_6582;
wire n_6996;
wire n_6974;
wire n_6765;
wire n_7577;
wire n_6921;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_6898;
wire n_6710;
wire n_5717;
wire n_7162;
wire n_5464;
wire n_6565;
wire n_5886;
wire n_7080;
wire n_3639;
wire n_7302;
wire n_6533;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_6960;
wire n_6426;
wire n_6634;
wire n_7180;
wire n_5610;
wire n_6836;
wire n_5239;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1979;
wire n_6972;
wire n_2924;
wire n_7111;
wire n_7549;
wire n_4111;
wire n_2484;
wire n_5785;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_6344;
wire n_5305;
wire n_5994;
wire n_4538;
wire n_6093;
wire n_6010;
wire n_7247;
wire n_6833;
wire n_2754;
wire n_5376;
wire n_2489;
wire n_7481;
wire n_5204;
wire n_7292;
wire n_2012;
wire n_4094;
wire n_3503;
wire n_7150;
wire n_2866;
wire n_3561;
wire n_2917;
wire n_2425;
wire n_3661;
wire n_3536;
wire n_4150;
wire n_4878;
wire n_6265;
wire n_6821;
wire n_3934;
wire n_4985;
wire n_6373;
wire n_6988;
wire n_5788;
wire n_3922;
wire n_3846;
wire n_5897;
wire n_6887;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_3074;
wire n_1999;
wire n_6676;
wire n_2372;
wire n_3673;
wire n_6347;
wire n_6492;
wire n_7016;
wire n_3768;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_5795;
wire n_7072;
wire n_5508;
wire n_5582;
wire n_4022;
wire n_7374;
wire n_7440;
wire n_4852;
wire n_7547;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_7201;
wire n_4035;
wire n_2316;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_5746;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_6648;
wire n_4601;
wire n_2687;
wire n_4220;
wire n_1944;
wire n_5630;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_7513;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_7413;
wire n_4403;
wire n_1981;
wire n_7540;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_5504;
wire n_7622;
wire n_7005;
wire n_4223;
wire n_7353;
wire n_6219;
wire n_6965;
wire n_5025;
wire n_2966;
wire n_2326;
wire n_6720;
wire n_2188;
wire n_6032;
wire n_7174;
wire n_6205;
wire n_6362;
wire n_6402;
wire n_4644;
wire n_7166;
wire n_4456;
wire n_5060;
wire n_7607;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_7591;
wire n_5775;
wire n_3311;
wire n_2748;
wire n_3272;
wire n_7282;
wire n_6491;
wire n_2898;
wire n_2717;
wire n_7151;
wire n_6229;
wire n_5731;
wire n_5581;
wire n_3691;
wire n_3628;
wire n_6668;
wire n_7446;
wire n_4235;
wire n_1945;
wire n_3018;
wire n_7053;
wire n_5831;
wire n_2573;
wire n_7473;
wire n_4435;
wire n_2939;
wire n_6835;
wire n_6419;
wire n_6039;
wire n_3807;
wire n_5884;
wire n_2447;
wire n_4764;
wire n_5653;
wire n_6258;
wire n_7070;
wire n_5394;
wire n_6755;
wire n_2774;
wire n_7276;
wire n_7351;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_6084;
wire n_4827;
wire n_7412;
wire n_7157;
wire n_6436;
wire n_2488;
wire n_7666;
wire n_6472;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_7211;
wire n_4399;
wire n_6531;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_4782;
wire n_4363;
wire n_2887;
wire n_4864;
wire n_2691;
wire n_7368;
wire n_3054;
wire n_4335;
wire n_6567;
wire n_5889;
wire n_6771;
wire n_2526;
wire n_6389;
wire n_2703;
wire n_2167;
wire n_5764;
wire n_5428;
wire n_6910;
wire n_6442;
wire n_3391;
wire n_6102;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_6441;
wire n_5543;
wire n_5678;
wire n_5935;
wire n_4865;
wire n_4056;
wire n_4564;
wire n_3840;
wire n_7677;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_5950;
wire n_2173;
wire n_3738;
wire n_5995;
wire n_6162;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_6331;
wire n_6006;
wire n_3245;
wire n_4417;
wire n_6109;
wire n_6278;
wire n_6787;
wire n_6872;
wire n_4899;
wire n_6208;
wire n_2119;
wire n_2157;
wire n_2552;
wire n_6632;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_7027;
wire n_3509;
wire n_3352;
wire n_5671;
wire n_3076;
wire n_6990;
wire n_3535;
wire n_2182;
wire n_6349;
wire n_3251;
wire n_2931;
wire n_7631;
wire n_6830;
wire n_5185;
wire n_6359;
wire n_3118;
wire n_3511;
wire n_3443;
wire n_2146;
wire n_7498;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_7377;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_6301;
wire n_3232;
wire n_2918;
wire n_5945;
wire n_2112;
wire n_2958;
wire n_6744;
wire n_4981;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_6439;
wire n_7381;
wire n_5565;
wire n_4081;
wire n_3132;
wire n_4407;
wire n_7291;
wire n_3951;
wire n_4894;
wire n_5780;
wire n_5643;
wire n_3238;
wire n_3210;
wire n_5846;
wire n_2036;
wire n_7430;
wire n_3267;
wire n_4995;
wire n_5524;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_6104;
wire n_3884;
wire n_6475;
wire n_6465;
wire n_3726;
wire n_6496;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_6998;
wire n_6145;
wire n_3577;
wire n_2820;
wire n_7305;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_4057;
wire n_4332;
wire n_4314;
wire n_3347;
wire n_3216;
wire n_3809;
wire n_2113;
wire n_7075;
wire n_7545;
wire n_4288;
wire n_6076;
wire n_3567;
wire n_6194;
wire n_5066;
wire n_3939;
wire n_6092;
wire n_7275;
wire n_5401;
wire n_6357;
wire n_5843;
wire n_4241;
wire n_3321;
wire n_7537;
wire n_3212;
wire n_3152;
wire n_2256;
wire n_7489;
wire n_5106;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_6335;
wire n_5883;
wire n_6985;
wire n_5319;
wire n_2247;
wire n_7451;
wire n_6238;
wire n_3705;
wire n_6548;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_2268;
wire n_3778;
wire n_5706;
wire n_5337;
wire n_6366;
wire n_3304;
wire n_3912;
wire n_7236;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_7269;
wire n_5223;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_6602;
wire n_4419;
wire n_4477;
wire n_6620;
wire n_3179;
wire n_6502;
wire n_3256;
wire n_7560;
wire n_7326;
wire n_7060;
wire n_2386;
wire n_7572;
wire n_3086;
wire n_6885;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_2568;
wire n_5364;
wire n_6529;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_5895;
wire n_4639;
wire n_6951;
wire n_3713;
wire n_3663;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_7169;
wire n_6423;
wire n_3246;
wire n_2495;
wire n_7140;
wire n_7233;
wire n_5088;
wire n_2302;
wire n_6558;
wire n_5457;
wire n_7352;
wire n_7134;
wire n_5532;
wire n_2069;
wire n_6950;
wire n_7246;
wire n_6525;
wire n_7650;
wire n_3434;
wire n_6631;
wire n_6892;
wire n_7663;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_7056;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_6683;
wire n_2482;
wire n_2677;
wire n_6292;
wire n_5544;
wire n_3832;
wire n_3987;
wire n_7339;
wire n_5987;
wire n_6180;
wire n_5352;
wire n_5824;
wire n_4991;
wire n_5538;
wire n_6658;
wire n_6264;
wire n_6925;
wire n_5919;
wire n_2329;
wire n_2142;
wire n_6176;
wire n_5410;
wire n_3332;
wire n_7146;
wire n_3048;
wire n_3937;
wire n_6124;
wire n_7672;
wire n_2203;
wire n_4525;
wire n_3782;
wire n_7482;
wire n_6864;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_7090;
wire n_3786;
wire n_7158;
wire n_2888;
wire n_7156;
wire n_5742;
wire n_3638;
wire n_5992;
wire n_6494;
wire n_5503;
wire n_4177;
wire n_6199;
wire n_3763;
wire n_2669;
wire n_2306;
wire n_5958;
wire n_6614;
wire n_3022;
wire n_4264;
wire n_7504;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_7360;
wire n_7681;
wire n_7301;
wire n_5129;
wire n_2149;
wire n_7375;
wire n_7102;
wire n_5500;
wire n_3060;
wire n_4276;
wire n_7366;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_5654;
wire n_2408;
wire n_7025;
wire n_5320;
wire n_3049;
wire n_6947;
wire n_5107;
wire n_5999;
wire n_4485;
wire n_7309;
wire n_4626;
wire n_6863;
wire n_6637;
wire n_6100;
wire n_6735;
wire n_2659;
wire n_4975;
wire n_6358;
wire n_5602;
wire n_3089;
wire n_6050;
wire n_2470;
wire n_7244;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_7610;
wire n_2551;
wire n_5903;
wire n_2682;
wire n_6371;
wire n_7043;
wire n_3440;
wire n_6171;
wire n_6510;
wire n_4569;
wire n_6468;
wire n_2699;
wire n_4897;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_2615;
wire n_3940;
wire n_5842;
wire n_6352;
wire n_2985;
wire n_5722;
wire n_7534;
wire n_5636;
wire n_5065;
wire n_2753;
wire n_7287;
wire n_7032;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_2868;
wire n_5492;
wire n_3141;
wire n_5084;
wire n_6850;
wire n_5667;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_7119;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_6354;
wire n_5918;
wire n_7634;
wire n_4503;
wire n_3507;
wire n_6959;
wire n_3821;
wire n_6909;
wire n_2700;
wire n_6332;
wire n_3367;
wire n_4464;
wire n_7006;
wire n_5877;
wire n_3096;
wire n_6306;
wire n_7682;
wire n_3496;
wire n_4114;
wire n_2544;
wire n_6434;
wire n_2356;
wire n_6751;
wire n_7068;
wire n_4556;
wire n_6322;
wire n_5454;
wire n_2620;
wire n_6667;
wire n_7526;
wire n_6530;
wire n_4089;
wire n_7376;
wire n_6156;
wire n_5913;
wire n_7268;
wire n_7044;
wire n_5621;
wire n_2919;
wire n_4327;
wire n_4218;
wire n_6429;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_7239;
wire n_2757;
wire n_5573;
wire n_6405;
wire n_6613;
wire n_4353;
wire n_2042;
wire n_6248;
wire n_2921;
wire n_2720;
wire n_4990;
wire n_6088;
wire n_5529;
wire n_6894;
wire n_7267;
wire n_4959;
wire n_4161;
wire n_5800;
wire n_3992;
wire n_2616;
wire n_4103;
wire n_4466;
wire n_2262;
wire n_6204;
wire n_2462;
wire n_3625;
wire n_7387;
wire n_7431;
wire n_7654;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_4844;
wire n_6296;
wire n_2979;
wire n_5257;
wire n_6290;
wire n_6288;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2548;
wire n_5645;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_5779;
wire n_4388;
wire n_4206;
wire n_6140;
wire n_7441;
wire n_4738;
wire n_6211;
wire n_3909;
wire n_6307;
wire n_6164;
wire n_3207;
wire n_3944;
wire n_7394;
wire n_4434;
wire n_4837;
wire n_7022;
wire n_3042;
wire n_1942;
wire n_6860;
wire n_2510;
wire n_4219;
wire n_3659;
wire n_2804;
wire n_2120;
wire n_5012;
wire n_4620;
wire n_5697;
wire n_7188;
wire n_7573;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_7087;
wire n_2222;
wire n_3510;
wire n_6147;
wire n_3218;
wire n_2667;
wire n_6515;
wire n_6011;
wire n_6645;
wire n_3150;
wire n_6984;
wire n_4325;
wire n_2413;
wire n_7193;
wire n_3775;
wire n_4133;
wire n_6897;
wire n_7256;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_6460;
wire n_4379;
wire n_7128;
wire n_7595;
wire n_2181;
wire n_6183;
wire n_7522;
wire n_5882;
wire n_4030;
wire n_7436;
wire n_4490;
wire n_3138;
wire n_7380;
wire n_7012;
wire n_4397;
wire n_7502;
wire n_2928;
wire n_7335;
wire n_7103;
wire n_4820;
wire n_6246;
wire n_3770;
wire n_5094;
wire n_6383;
wire n_4938;
wire n_7020;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_2723;
wire n_5672;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_5548;
wire n_5601;
wire n_7248;
wire n_7662;
wire n_3855;
wire n_2054;
wire n_5339;
wire n_4931;
wire n_6099;
wire n_3158;
wire n_5693;
wire n_2623;
wire n_3113;
wire n_6904;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_2856;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_7533;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_6626;
wire n_6563;
wire n_5486;
wire n_6611;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_5599;
wire n_6116;
wire n_7186;
wire n_4356;
wire n_6819;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_6473;
wire n_4291;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_6310;
wire n_2982;
wire n_2481;
wire n_7429;
wire n_3545;
wire n_6688;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_2339;
wire n_7148;
wire n_5782;
wire n_6714;
wire n_4637;
wire n_7017;
wire n_7250;
wire n_7462;
wire n_7658;
wire n_4935;
wire n_6365;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_5608;
wire n_3741;
wire n_3410;
wire n_7401;
wire n_6828;
wire n_2029;
wire n_5298;
wire n_6355;
wire n_5596;
wire n_4413;
wire n_6777;
wire n_5728;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_6420;
wire n_6945;
wire n_2882;
wire n_7356;
wire n_2338;
wire n_5726;
wire n_7288;
wire n_7637;
wire n_7124;
wire n_3672;
wire n_7294;
wire n_5290;
wire n_3197;
wire n_7018;
wire n_3109;
wire n_2721;
wire n_7321;
wire n_5095;
wire n_3002;
wire n_6754;
wire n_6583;
wire n_6622;
wire n_6936;
wire n_5324;
wire n_3897;
wire n_5928;
wire n_3845;
wire n_7108;
wire n_6882;
wire n_2081;
wire n_7585;
wire n_4570;
wire n_7386;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_5019;
wire n_5911;
wire n_7362;
wire n_7417;
wire n_2418;
wire n_7187;
wire n_5589;
wire n_5841;
wire n_2179;
wire n_2521;
wire n_7544;
wire n_3458;
wire n_5712;
wire n_3330;
wire n_4606;
wire n_6166;
wire n_4774;
wire n_2477;
wire n_6966;
wire n_3887;
wire n_7542;
wire n_6781;
wire n_7255;
wire n_4093;
wire n_7120;
wire n_7218;
wire n_4672;
wire n_7147;
wire n_3519;
wire n_7221;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_2367;
wire n_4766;
wire n_5633;
wire n_2896;
wire n_4074;
wire n_4600;
wire n_6980;
wire n_1927;
wire n_5583;
wire n_4460;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_6064;
wire n_6110;
wire n_6237;
wire n_7196;
wire n_2255;
wire n_2272;
wire n_6341;
wire n_1965;
wire n_6590;
wire n_1941;
wire n_5501;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_6697;
wire n_5652;
wire n_6453;
wire n_6135;
wire n_7559;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_7081;
wire n_3189;
wire n_2066;
wire n_6449;
wire n_3154;
wire n_6141;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_2220;
wire n_4349;
wire n_7584;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_6983;
wire n_1935;
wire n_6036;
wire n_3366;
wire n_2696;
wire n_4863;
wire n_7222;
wire n_3242;
wire n_6071;
wire n_3525;
wire n_3486;
wire n_6808;
wire n_2405;
wire n_6724;
wire n_3995;
wire n_2953;
wire n_2088;
wire n_4036;
wire n_6571;
wire n_5100;
wire n_7470;
wire n_5849;
wire n_6251;
wire n_7400;
wire n_2578;
wire n_3483;
wire n_6635;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_7623;
wire n_3524;
wire n_5616;
wire n_7597;
wire n_5034;
wire n_6733;
wire n_7071;
wire n_5988;
wire n_6467;
wire n_6035;
wire n_3549;
wire n_6522;
wire n_7109;
wire n_2092;
wire n_5959;
wire n_2075;
wire n_7645;
wire n_3658;
wire n_6732;
wire n_4807;
wire n_6562;
wire n_6150;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_4230;
wire n_3419;
wire n_2053;
wire n_1958;
wire n_5917;
wire n_5754;
wire n_6016;
wire n_3784;
wire n_3941;
wire n_2969;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_7212;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_5628;
wire n_6726;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_7009;
wire n_6554;
wire n_6689;
wire n_2731;
wire n_6143;
wire n_5614;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_7355;
wire n_3979;
wire n_7365;
wire n_4582;
wire n_2998;
wire n_6277;
wire n_4684;
wire n_7395;
wire n_5981;
wire n_6095;
wire n_7671;
wire n_6247;
wire n_4840;
wire n_3162;
wire n_2760;
wire n_6880;
wire n_3377;
wire n_3749;
wire n_5720;
wire n_3962;
wire n_2304;
wire n_5325;
wire n_5696;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_6499;
wire n_6837;
wire n_4423;
wire n_4096;
wire n_7393;
wire n_2881;
wire n_6616;
wire n_3282;
wire n_3231;
wire n_1966;
wire n_6946;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_5759;
wire n_4478;
wire n_5753;
wire n_2646;
wire n_5536;
wire n_7484;
wire n_5173;
wire n_6305;
wire n_6317;
wire n_3920;
wire n_4890;
wire n_5691;
wire n_5794;
wire n_5027;
wire n_5647;
wire n_7231;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_7272;
wire n_4106;
wire n_3717;
wire n_5738;
wire n_2743;
wire n_2675;
wire n_7649;
wire n_3052;
wire n_5215;
wire n_7324;
wire n_6693;
wire n_3743;
wire n_6734;
wire n_7135;
wire n_7014;
wire n_1932;
wire n_4721;
wire n_5597;
wire n_5635;
wire n_6382;
wire n_7328;
wire n_1983;
wire n_7635;
wire n_6404;
wire n_5975;
wire n_4029;
wire n_3870;
wire n_6379;
wire n_7066;
wire n_4496;
wire n_3529;
wire n_7358;
wire n_1977;
wire n_2153;
wire n_6235;
wire n_4338;
wire n_7277;
wire n_6504;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_7265;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_6789;
wire n_7184;
wire n_6440;
wire n_6417;
wire n_2318;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_7491;
wire n_5942;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_7219;
wire n_7479;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_7270;
wire n_5940;
wire n_7390;
wire n_5121;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_5555;
wire n_6914;
wire n_2446;
wire n_3488;
wire n_7182;
wire n_4547;
wire n_2893;
wire n_4004;
wire n_2588;
wire n_2962;
wire n_5784;
wire n_6272;
wire n_6484;
wire n_7674;
wire n_6236;
wire n_5576;
wire n_4668;
wire n_4953;
wire n_5466;
wire n_6958;
wire n_6840;
wire n_3898;
wire n_6871;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_6768;
wire n_4759;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_7506;
wire n_2340;
wire n_3552;
wire n_6717;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_7048;
wire n_5578;
wire n_2361;
wire n_4113;
wire n_1998;
wire n_4686;
wire n_5530;
wire n_3759;
wire n_6196;
wire n_7416;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_5741;
wire n_5991;
wire n_3933;
wire n_7330;
wire n_3206;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_5221;
wire n_6992;
wire n_4183;
wire n_4068;
wire n_4872;
wire n_6000;
wire n_4233;
wire n_7283;
wire n_3192;
wire n_7099;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_6448;
wire n_2649;
wire n_6655;
wire n_7304;
wire n_5792;
wire n_6657;
wire n_1929;
wire n_5575;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_7626;
wire n_3742;
wire n_7474;
wire n_2252;
wire n_7612;
wire n_6113;
wire n_4819;
wire n_6242;
wire n_7088;
wire n_6519;
wire n_4900;
wire n_2576;
wire n_6842;
wire n_7588;
wire n_3390;
wire n_6206;
wire n_6414;
wire n_3746;
wire n_2373;
wire n_3817;
wire n_2745;
wire n_6801;
wire n_2493;
wire n_4930;
wire n_7680;
wire n_5276;
wire n_6308;
wire n_7398;
wire n_6906;
wire n_5078;
wire n_4537;
wire n_7230;
wire n_2885;
wire n_6629;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_6968;
wire n_4282;
wire n_6615;
wire n_3485;
wire n_4180;
wire n_7378;
wire n_3839;
wire n_5205;
wire n_3333;
wire n_5651;
wire n_2845;
wire n_6144;
wire n_4143;
wire n_4659;
wire n_6188;
wire n_2602;
wire n_5819;
wire n_4579;
wire n_4616;
wire n_3014;
wire n_2547;
wire n_5998;
wire n_6398;
wire n_5023;
wire n_4105;
wire n_5721;
wire n_5673;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_3329;
wire n_2765;
wire n_6415;
wire n_2994;
wire n_6857;
wire n_3135;
wire n_2401;
wire n_5476;
wire n_2003;
wire n_5856;
wire n_5446;
wire n_4895;
wire n_6722;
wire n_3573;
wire n_3148;
wire n_6428;
wire n_5944;
wire n_7618;
wire n_2264;
wire n_3534;
wire n_6413;
wire n_7679;
wire n_4275;
wire n_3970;
wire n_6361;
wire n_3438;
wire n_6231;
wire n_4098;
wire n_5684;
wire n_5861;
wire n_5976;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_2184;
wire n_5312;
wire n_5850;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_5111;
wire n_5890;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_7167;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_7643;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_6712;
wire n_5687;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_5839;
wire n_3397;
wire n_3740;
wire n_6953;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_2977;
wire n_6303;
wire n_6474;
wire n_6182;
wire n_3723;
wire n_5674;
wire n_3600;
wire n_6573;
wire n_4134;
wire n_6053;
wire n_7234;
wire n_2836;
wire n_5682;
wire n_6392;
wire n_2130;
wire n_5167;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_5612;
wire n_6125;
wire n_6599;
wire n_6685;
wire n_2850;
wire n_4251;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_6560;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_6253;
wire n_4740;
wire n_7382;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_7615;
wire n_5898;
wire n_2221;
wire n_3576;
wire n_7298;
wire n_7581;
wire n_4049;
wire n_6641;
wire n_5214;
wire n_3862;
wire n_5487;
wire n_5563;
wire n_6593;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_6673;
wire n_7172;
wire n_7074;
wire n_5497;
wire n_4724;
wire n_5832;
wire n_7190;
wire n_7112;
wire n_7678;
wire n_5526;
wire n_2818;
wire n_3646;
wire n_6367;
wire n_2129;
wire n_3345;
wire n_4546;
wire n_6195;
wire n_6356;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_7001;
wire n_5593;
wire n_5021;
wire n_6514;
wire n_2772;
wire n_7369;
wire n_5444;
wire n_1924;
wire n_4382;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_6559;
wire n_7359;
wire n_2260;
wire n_5389;
wire n_7144;
wire n_4833;
wire n_6841;
wire n_3056;
wire n_2345;
wire n_5110;
wire n_6653;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_7450;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_5737;
wire n_2579;
wire n_6825;
wire n_6923;
wire n_4228;
wire n_4401;
wire n_6112;
wire n_2788;
wire n_6547;
wire n_2984;
wire n_6198;
wire n_7439;
wire n_3364;
wire n_5560;
wire n_6399;
wire n_3201;
wire n_6275;
wire n_5666;
wire n_6575;
wire n_3472;
wire n_6151;
wire n_2874;
wire n_5179;
wire n_7227;
wire n_7040;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_7325;
wire n_4968;
wire n_6469;
wire n_6756;
wire n_5030;
wire n_3949;
wire n_5961;
wire n_3543;
wire n_7191;
wire n_7459;
wire n_7096;
wire n_3050;
wire n_3903;
wire n_4834;
wire n_5272;
wire n_2742;
wire n_2183;
wire n_3314;
wire n_4158;
wire n_6826;
wire n_2360;
wire n_6015;
wire n_3254;
wire n_5361;
wire n_5683;
wire n_4171;
wire n_5847;
wire n_7551;
wire n_4045;
wire n_6678;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_5740;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_5729;
wire n_7485;
wire n_6748;
wire n_2030;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_6752;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_6553;
wire n_2209;
wire n_7652;
wire n_6500;
wire n_4270;
wire n_2797;
wire n_7051;
wire n_5152;
wire n_2321;
wire n_3680;
wire n_6628;
wire n_6297;
wire n_5905;
wire n_3497;
wire n_6975;
wire n_5409;
wire n_6329;
wire n_2940;
wire n_7536;
wire n_5688;
wire n_2612;
wire n_5128;
wire n_4566;
wire n_2841;
wire n_6293;
wire n_3322;
wire n_4576;
wire n_2427;
wire n_2505;
wire n_7676;
wire n_4061;
wire n_3250;
wire n_2070;
wire n_7553;
wire n_6905;
wire n_7425;
wire n_2594;
wire n_5798;
wire n_6381;
wire n_6521;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_5986;
wire n_3112;
wire n_2349;
wire n_6581;
wire n_3874;
wire n_6215;
wire n_7095;
wire n_5415;
wire n_4676;
wire n_5770;
wire n_7064;
wire n_5892;
wire n_4544;
wire n_2170;
wire n_6577;
wire n_6899;
wire n_5676;
wire n_7307;
wire n_6545;
wire n_5802;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_6370;
wire n_3266;
wire n_7210;
wire n_4646;
wire n_5769;
wire n_6065;
wire n_7039;
wire n_6987;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_6190;
wire n_6859;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_6309;
wire n_6623;
wire n_2426;
wire n_6527;
wire n_7443;
wire n_5341;
wire n_4320;
wire n_5930;
wire n_5814;
wire n_4881;
wire n_5979;
wire n_5271;
wire n_5089;
wire n_7015;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_6929;
wire n_4012;
wire n_5518;
wire n_4636;
wire n_5637;
wire n_4584;
wire n_5622;
wire n_3910;
wire n_4711;
wire n_3319;
wire n_7348;
wire n_5240;
wire n_3335;
wire n_5813;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_5546;
wire n_2689;
wire n_3259;
wire n_7143;
wire n_5482;
wire n_7312;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_7155;
wire n_3688;
wire n_6865;
wire n_3016;
wire n_5393;
wire n_2599;
wire n_6535;
wire n_3338;
wire n_7213;
wire n_3414;
wire n_4671;
wire n_4209;
wire n_5966;
wire n_7456;
wire n_5041;
wire n_7420;
wire n_5431;
wire n_3261;
wire n_2200;
wire n_6482;
wire n_5026;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_5059;
wire n_5505;
wire n_3127;
wire n_3732;
wire n_6605;
wire n_4250;
wire n_5329;
wire n_3596;
wire n_4699;
wire n_7007;
wire n_3906;
wire n_4127;
wire n_3297;
wire n_2683;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_5908;
wire n_6018;
wire n_4202;
wire n_7168;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_5939;
wire n_7177;
wire n_3766;
wire n_2880;
wire n_7379;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_7444;
wire n_5931;
wire n_7435;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_7030;
wire n_5420;
wire n_6311;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_6424;
wire n_6654;
wire n_6816;
wire n_6220;
wire n_3621;
wire n_5234;
wire n_6740;
wire n_7122;
wire n_5835;
wire n_7049;
wire n_7567;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_6029;
wire n_6879;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_5679;
wire n_3710;
wire n_5938;
wire n_6702;
wire n_4155;
wire n_2031;
wire n_3891;
wire n_5891;
wire n_4144;
wire n_5724;
wire n_5774;
wire n_2165;
wire n_6452;
wire n_3379;
wire n_4374;
wire n_6791;
wire n_3532;
wire n_5131;
wire n_7280;
wire n_2127;
wire n_6915;
wire n_7110;
wire n_7511;
wire n_6856;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_7232;
wire n_4548;
wire n_7345;
wire n_5923;
wire n_5790;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_6364;
wire n_6451;
wire n_6552;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_6328;
wire n_4816;
wire n_6363;
wire n_2983;
wire n_7159;
wire n_3810;
wire n_2715;
wire n_6132;
wire n_6578;
wire n_6406;
wire n_5598;
wire n_2085;
wire n_5306;
wire n_6978;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_2672;
wire n_2651;
wire n_4358;
wire n_7477;
wire n_5147;
wire n_3656;
wire n_6918;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_4793;
wire n_7363;
wire n_6612;
wire n_5677;
wire n_4168;
wire n_3446;
wire n_5997;
wire n_5511;
wire n_5680;
wire n_3028;
wire n_4806;
wire n_4350;
wire n_7295;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_5280;
wire n_6375;
wire n_6479;
wire n_6866;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_3389;
wire n_6170;
wire n_1931;
wire n_4187;
wire n_4166;
wire n_6447;
wire n_6263;
wire n_7093;
wire n_5206;
wire n_3222;
wire n_7466;
wire n_5419;
wire n_6130;
wire n_2970;
wire n_7651;
wire n_2235;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_3755;
wire n_5803;
wire n_4258;
wire n_6014;
wire n_4498;
wire n_6935;
wire n_7530;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_5985;
wire n_2944;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_6907;
wire n_6158;
wire n_7661;
wire n_6541;
wire n_3262;
wire n_6119;
wire n_5018;
wire n_4006;
wire n_5896;
wire n_4861;
wire n_3690;
wire n_2358;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_2833;
wire n_4712;
wire n_6226;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_7145;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_6338;
wire n_1950;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_7467;
wire n_5097;
wire n_2750;
wire n_5730;
wire n_3899;
wire n_7550;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_5816;
wire n_4069;
wire n_2784;
wire n_7541;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_7241;
wire n_2557;
wire n_5300;
wire n_4850;
wire n_6625;
wire n_3781;
wire n_4912;
wire n_4813;
wire n_7464;
wire n_2590;
wire n_6302;
wire n_2330;
wire n_5748;
wire n_2942;
wire n_6759;
wire n_5525;
wire n_3106;
wire n_3328;
wire n_6706;
wire n_3889;
wire n_6139;
wire n_4256;
wire n_7434;
wire n_7636;
wire n_7054;
wire n_6999;
wire n_4224;
wire n_6403;
wire n_3508;
wire n_6483;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_6228;
wire n_5650;
wire n_2636;
wire n_1951;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_7299;
wire n_4702;
wire n_6888;
wire n_4252;
wire n_4457;
wire n_6063;
wire n_6800;
wire n_5139;
wire n_2319;
wire n_6922;
wire n_3481;
wire n_5481;
wire n_6890;
wire n_7503;
wire n_2808;
wire n_6070;
wire n_2676;
wire n_2679;
wire n_6651;
wire n_5821;
wire n_7091;
wire n_4491;
wire n_7296;
wire n_6647;
wire n_7273;
wire n_2930;
wire n_5733;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_5871;
wire n_7543;
wire n_2611;
wire n_4261;
wire n_6184;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_7507;
wire n_2698;
wire n_5043;
wire n_7555;
wire n_5707;
wire n_4001;
wire n_3047;
wire n_2454;
wire n_4371;
wire n_5836;
wire n_5281;
wire n_6716;
wire n_6422;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_4268;
wire n_5048;
wire n_5521;
wire n_7578;
wire n_5028;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_7475;
wire n_4194;
wire n_5585;
wire n_6397;
wire n_4824;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_2990;
wire n_7033;
wire n_6121;
wire n_3119;
wire n_7531;
wire n_4142;
wire n_4082;
wire n_5561;
wire n_3479;
wire n_4085;
wire n_4260;
wire n_4073;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_6981;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_6954;
wire n_3279;
wire n_2621;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_5875;
wire n_4262;
wire n_2671;
wire n_6646;
wire n_4720;
wire n_7131;
wire n_6903;
wire n_4685;
wire n_6101;
wire n_5968;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_6941;
wire n_2073;
wire n_4511;
wire n_5812;
wire n_6148;
wire n_5515;
wire n_6106;
wire n_6604;
wire n_4014;
wire n_7418;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_5607;
wire n_4175;
wire n_2005;
wire n_4648;
wire n_5006;
wire n_6566;
wire n_5734;
wire n_6081;
wire n_4892;
wire n_7204;
wire n_3823;
wire n_4173;
wire n_4970;
wire n_3816;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_6047;
wire n_2960;
wire n_5438;
wire n_4627;
wire n_7448;
wire n_7354;
wire n_6244;
wire n_2290;
wire n_6861;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_2145;
wire n_5725;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_7571;
wire n_5163;
wire n_2039;
wire n_5768;
wire n_4961;
wire n_7556;
wire n_3753;
wire n_7640;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_7422;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_6588;
wire n_3396;
wire n_7050;
wire n_4023;
wire n_4420;
wire n_5685;
wire n_5773;
wire n_7136;
wire n_7318;
wire n_6055;
wire n_5138;
wire n_5374;
wire n_6108;
wire n_2116;
wire n_6165;
wire n_6621;
wire n_2320;
wire n_7175;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_6323;
wire n_4396;
wire n_5127;
wire n_6587;
wire n_4367;
wire n_6480;
wire n_2087;
wire n_6731;
wire n_5485;
wire n_5766;
wire n_5216;
wire n_6597;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_6933;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_6881;
wire n_7289;
wire n_5805;
wire n_7665;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_6216;
wire n_3830;
wire n_2585;
wire n_6817;
wire n_7170;
wire n_7314;
wire n_2725;
wire n_6949;
wire n_6509;
wire n_5175;
wire n_3883;
wire n_7260;
wire n_4152;
wire n_2565;
wire n_7263;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_6911;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_5900;
wire n_3466;
wire n_4962;
wire n_6327;
wire n_2595;
wire n_6607;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_7509;
wire n_7209;
wire n_5171;
wire n_3586;
wire n_6401;
wire n_5554;
wire n_6227;
wire n_7240;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_5427;
wire n_5639;
wire n_3065;
wire n_4361;
wire n_5417;
wire n_4614;
wire n_2681;
wire n_3103;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_7609;
wire n_7278;
wire n_7630;
wire n_2775;
wire n_6416;
wire n_4693;
wire n_5488;
wire n_4326;
wire n_6695;
wire n_3557;
wire n_2230;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_6127;
wire n_7565;
wire n_2851;
wire n_4305;
wire n_5781;
wire n_6600;
wire n_2490;
wire n_7410;
wire n_4213;
wire n_2849;
wire n_7097;
wire n_3692;
wire n_2204;
wire n_6421;
wire n_5747;
wire n_7414;
wire n_7495;
wire n_5969;
wire n_4929;
wire n_1961;
wire n_4964;
wire n_6079;
wire n_4802;
wire n_6192;
wire n_6458;
wire n_4139;
wire n_3029;
wire n_6746;
wire n_2508;
wire n_4031;
wire n_7586;
wire n_6719;
wire n_2416;
wire n_5437;
wire n_5826;
wire n_7659;
wire n_3881;
wire n_2461;
wire n_6506;
wire n_2243;
wire n_4583;
wire n_6287;
wire n_6662;
wire n_4210;
wire n_5245;
wire n_7189;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_2368;
wire n_6851;
wire n_6687;
wire n_2890;
wire n_6884;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_4540;
wire n_3961;
wire n_6780;
wire n_6513;
wire n_4891;
wire n_6619;
wire n_5603;
wire n_6804;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_5716;
wire n_3993;
wire n_4940;
wire n_6516;
wire n_5208;
wire n_7490;
wire n_3588;
wire n_6924;
wire n_2308;
wire n_4590;
wire n_7492;
wire n_5606;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_5456;
wire n_3160;
wire n_7073;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_6040;
wire n_3847;
wire n_4946;
wire n_4906;
wire n_5727;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_7114;
wire n_5347;
wire n_3298;
wire n_3033;
wire n_2824;
wire n_6788;
wire n_2440;
wire n_4883;
wire n_2923;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_6393;
wire n_2333;
wire n_2916;
wire n_6249;
wire n_4297;
wire n_5833;
wire n_6849;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_7271;
wire n_3991;
wire n_3134;
wire n_6572;
wire n_4172;
wire n_4791;
wire n_6739;
wire n_4536;
wire n_5149;
wire n_5967;
wire n_2463;
wire n_5151;
wire n_7569;
wire n_7003;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_6666;
wire n_2472;
wire n_4611;
wire n_6812;
wire n_4755;
wire n_5982;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_7419;
wire n_5827;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_6200;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_6123;
wire n_6934;
wire n_2589;
wire n_7094;
wire n_7500;
wire n_3482;
wire n_6082;
wire n_2233;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_7129;
wire n_3956;
wire n_5758;
wire n_5323;
wire n_3572;
wire n_4215;
wire n_6952;
wire n_4280;
wire n_7062;
wire n_3375;
wire n_4047;
wire n_5471;
wire n_7642;
wire n_5434;
wire n_2082;
wire n_5941;
wire n_7045;
wire n_5879;
wire n_3167;
wire n_5558;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_7238;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_7126;
wire n_5669;
wire n_3854;
wire n_2468;
wire n_3078;
wire n_6979;
wire n_6203;
wire n_7405;
wire n_3253;
wire n_7207;
wire n_4027;
wire n_2280;
wire n_7454;
wire n_4599;
wire n_5830;
wire n_6796;
wire n_3363;
wire n_4812;
wire n_5760;
wire n_6368;
wire n_3689;
wire n_6556;
wire n_2020;
wire n_4628;
wire n_5668;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_5878;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_5765;
wire n_3950;
wire n_4458;
wire n_6596;
wire n_4121;
wire n_5090;
wire n_6870;
wire n_7639;
wire n_4476;
wire n_5613;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_7251;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_6080;
wire n_7059;
wire n_7035;
wire n_5571;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_6713;
wire n_5513;
wire n_6747;
wire n_6281;
wire n_4803;
wire n_5972;
wire n_4079;
wire n_4091;
wire n_5916;
wire n_5984;
wire n_7029;
wire n_7317;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_6094;
wire n_2935;
wire n_6444;
wire n_5132;
wire n_5191;
wire n_6333;
wire n_6262;
wire n_3085;
wire n_5869;
wire n_5925;
wire n_6240;
wire n_5359;
wire n_6412;
wire n_2574;
wire n_5293;
wire n_7220;
wire n_4316;
wire n_3697;
wire n_7438;
wire n_2638;
wire n_7515;
wire n_7574;
wire n_4044;
wire n_4062;
wire n_6684;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_7065;
wire n_5510;
wire n_6046;
wire n_2016;
wire n_6973;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_7285;
wire n_5200;
wire n_5659;
wire n_5618;
wire n_6325;
wire n_2867;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_6737;
wire n_6454;
wire n_4253;
wire n_5356;
wire n_6721;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_7008;
wire n_3517;
wire n_3100;
wire n_2522;
wire n_6111;
wire n_7505;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_6260;
wire n_7501;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_6665;
wire n_7566;
wire n_7055;
wire n_3506;
wire n_3605;
wire n_2409;
wire n_5858;
wire n_5817;
wire n_6690;
wire n_3402;
wire n_5723;
wire n_5295;
wire n_6137;
wire n_4679;
wire n_4115;
wire n_6201;
wire n_7113;
wire n_4998;
wire n_2988;
wire n_1970;
wire n_2766;
wire n_5627;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_7242;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_6461;
wire n_2205;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_6212;
wire n_3401;
wire n_6908;
wire n_3226;
wire n_6570;
wire n_6498;
wire n_3902;
wire n_4730;
wire n_7228;
wire n_6692;
wire n_6074;
wire n_2779;
wire n_7561;
wire n_6380;
wire n_3654;
wire n_2164;
wire n_5996;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_6045;
wire n_4713;
wire n_5137;
wire n_6505;
wire n_2811;
wire n_3348;
wire n_7415;
wire n_5796;
wire n_7598;
wire n_6320;
wire n_6489;
wire n_6068;
wire n_3358;
wire n_5791;
wire n_2121;
wire n_4204;
wire n_5098;
wire n_6772;
wire n_1991;
wire n_2224;
wire n_6877;
wire n_6823;
wire n_6806;
wire n_7426;
wire n_5906;
wire n_4743;
wire n_3805;
wire n_3825;
wire n_6831;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_7217;
wire n_2692;
wire n_2008;
wire n_6284;
wire n_7058;
wire n_4654;
wire n_6157;
wire n_5423;
wire n_7497;
wire n_6785;
wire n_6374;
wire n_6930;
wire n_4733;
wire n_3792;
wire n_6017;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_2283;
wire n_3278;
wire n_4269;
wire n_4695;
wire n_6838;
wire n_5736;
wire n_6937;
wire n_6443;
wire n_3312;
wire n_6105;
wire n_2197;
wire n_7558;
wire n_2199;
wire n_5069;
wire n_7442;
wire n_5700;
wire n_6543;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_6091;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_6674;
wire n_2480;
wire n_6034;
wire n_7499;
wire n_2363;
wire n_4072;
wire n_5579;
wire n_7085;
wire n_4781;
wire n_3606;
wire n_6652;
wire n_7098;
wire n_5004;
wire n_2550;
wire n_6762;
wire n_7341;
wire n_4424;
wire n_7611;
wire n_7391;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_5837;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_6895;
wire n_3878;
wire n_7646;
wire n_4450;
wire n_5642;
wire n_3553;
wire n_7224;
wire n_5880;
wire n_6169;
wire n_4746;
wire n_7524;
wire n_5713;
wire n_6005;
wire n_7627;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_3850;
wire n_4459;
wire n_2996;
wire n_5793;
wire n_5591;
wire n_4050;
wire n_7496;
wire n_2315;
wire n_3228;
wire n_2102;
wire n_5623;
wire n_5681;
wire n_4853;
wire n_7399;
wire n_2422;
wire n_6213;
wire n_2239;
wire n_6118;
wire n_5256;
wire n_2950;
wire n_7605;
wire n_5220;
wire n_5732;
wire n_3852;
wire n_5178;
wire n_4520;
wire n_6814;
wire n_7342;
wire n_2057;
wire n_4008;
wire n_5507;
wire n_7214;
wire n_7472;
wire n_5077;
wire n_5872;
wire n_3858;
wire n_7408;
wire n_6115;
wire n_4502;
wire n_6858;
wire n_3032;
wire n_4851;
wire n_5735;
wire n_7254;
wire n_6944;
wire n_7384;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_3924;
wire n_4571;
wire n_2006;
wire n_6430;
wire n_6193;
wire n_5314;
wire n_6462;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_6757;
wire n_6822;
wire n_2535;
wire n_4205;
wire n_5953;
wire n_2726;
wire n_7599;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_6779;
wire n_6518;
wire n_6797;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_5952;
wire n_4739;
wire n_5820;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_5718;
wire n_6916;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_3926;
wire n_6152;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_2854;
wire n_4181;
wire n_5777;
wire n_2764;
wire n_7046;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_4153;
wire n_5156;
wire n_5926;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_4783;
wire n_2964;
wire n_3769;
wire n_6589;
wire n_7579;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_7173;
wire n_5951;
wire n_7092;
wire n_2442;
wire n_6197;
wire n_6971;
wire n_1943;
wire n_7460;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_6154;
wire n_7344;
wire n_6020;
wire n_2883;
wire n_4182;
wire n_2912;
wire n_4825;
wire n_5701;
wire n_4440;
wire n_4549;
wire n_3955;
wire n_7079;
wire n_5120;
wire n_5470;
wire n_4565;
wire n_7675;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_5797;
wire n_6696;
wire n_4839;
wire n_5222;
wire n_5743;
wire n_4016;
wire n_6210;
wire n_5772;
wire n_3435;
wire n_3575;
wire n_6964;
wire n_5801;
wire n_6117;
wire n_4231;
wire n_6202;
wire n_7279;
wire n_3165;
wire n_7670;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_6681;
wire n_4083;
wire n_1937;
wire n_5971;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_2381;
wire n_6661;
wire n_3303;
wire n_6640;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_7371;
wire n_6962;
wire n_4101;
wire n_6455;
wire n_3591;
wire n_2196;
wire n_4273;
wire n_3024;
wire n_7606;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_6963;
wire n_6644;
wire n_4389;
wire n_6896;
wire n_3930;
wire n_4448;
wire n_6832;
wire n_2161;
wire n_6160;
wire n_7564;
wire n_2404;
wire n_2083;
wire n_6718;
wire n_2503;
wire n_6542;
wire n_1936;
wire n_6031;
wire n_5502;
wire n_2027;
wire n_5568;
wire n_2642;
wire n_2500;
wire n_7653;
wire n_5656;
wire n_6763;
wire n_4831;
wire n_2513;
wire n_5974;
wire n_3480;
wire n_2695;
wire n_3057;
wire n_3194;
wire n_6280;
wire n_2414;
wire n_6438;
wire n_3662;
wire n_6316;
wire n_7383;
wire n_4319;
wire n_5474;
wire n_2229;
wire n_4596;
wire n_5413;
wire n_6758;
wire n_2004;
wire n_5412;
wire n_3694;
wire n_2586;
wire n_6069;
wire n_5752;
wire n_6874;
wire n_4726;
wire n_4751;
wire n_4222;
wire n_2274;
wire n_3225;
wire n_2972;
wire n_6030;
wire n_6077;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_6299;
wire n_4474;
wire n_6386;
wire n_5217;
wire n_5957;
wire n_2511;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_7655;
wire n_5490;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_6708;
wire n_7433;
wire n_4366;
wire n_4009;
wire n_7347;
wire n_4580;
wire n_6792;
wire n_7633;
wire n_6177;
wire n_5912;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_6033;
wire n_5557;
wire n_7397;
wire n_7389;
wire n_5472;
wire n_7602;
wire n_2955;
wire n_4112;
wire n_6002;
wire n_4337;
wire n_5711;
wire n_4138;
wire n_7554;
wire n_5396;
wire n_5335;
wire n_2520;
wire n_6557;
wire n_7300;
wire n_2134;
wire n_5960;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_7532;
wire n_5143;
wire n_4238;
wire n_6142;
wire n_6917;
wire n_7510;
wire n_2374;
wire n_5859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_2396;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_6163;
wire n_4635;
wire n_3501;
wire n_7118;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_6285;
wire n_6778;
wire n_6025;
wire n_7257;
wire n_4242;
wire n_6862;
wire n_6319;
wire n_7067;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_3180;
wire n_5283;
wire n_7669;
wire n_5268;
wire n_6318;
wire n_4561;
wire n_2639;
wire n_6089;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_6315;
wire n_3186;
wire n_4955;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_3650;
wire n_5840;
wire n_2761;
wire n_6343;
wire n_3157;
wire n_2537;
wire n_2144;
wire n_6049;
wire n_6919;
wire n_7423;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_6052;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_7069;
wire n_6886;
wire n_1949;
wire n_2936;
wire n_1946;
wire n_6912;
wire n_5914;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_6061;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_7252;
wire n_5542;
wire n_4394;
wire n_7133;
wire n_6883;
wire n_5519;
wire n_3101;
wire n_3669;
wire n_6009;
wire n_7061;
wire n_5278;
wire n_2663;
wire n_7518;
wire n_5586;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_6378;
wire n_5187;
wire n_4944;
wire n_5675;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_2632;
wire n_6601;
wire n_5771;
wire n_7216;
wire n_6407;
wire n_6749;
wire n_6839;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_6051;
wire n_4716;
wire n_4942;
wire n_6217;
wire n_6680;
wire n_5844;
wire n_2432;
wire n_6532;
wire n_3405;
wire n_4745;
wire n_6155;
wire n_6446;
wire n_6738;
wire n_6250;
wire n_7458;
wire n_7614;
wire n_2337;
wire n_3907;
wire n_6736;
wire n_5344;
wire n_6526;
wire n_4629;
wire n_6339;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_6350;
wire n_7013;
wire n_3306;
wire n_5662;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_3986;
wire n_4376;
wire n_5705;
wire n_4753;
wire n_4552;
wire n_7656;
wire n_3885;
wire n_6845;
wire n_7105;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_6829;
wire n_5574;
wire n_5126;
wire n_6508;
wire n_2214;
wire n_3427;
wire n_2055;
wire n_4067;
wire n_5553;
wire n_4042;
wire n_4176;
wire n_7570;
wire n_4385;
wire n_3320;
wire n_7052;
wire n_5009;
wire n_7262;
wire n_2688;
wire n_5368;
wire n_5626;
wire n_6603;
wire n_6114;
wire n_6576;
wire n_3651;
wire n_4333;
wire n_7364;
wire n_3359;
wire n_7208;
wire n_6245;
wire n_2865;
wire n_2706;
wire n_5499;
wire n_6703;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_7202;
wire n_4246;
wire n_3580;
wire n_7011;
wire n_2139;
wire n_4609;
wire n_7621;
wire n_5291;
wire n_5876;
wire n_6970;
wire n_5114;
wire n_2674;
wire n_6409;
wire n_6704;
wire n_6876;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_7028;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_7313;
wire n_6255;
wire n_7320;
wire n_7343;
wire n_5288;
wire n_2305;
wire n_5540;
wire n_5699;
wire n_7525;
wire n_2450;
wire n_3447;
wire n_5810;
wire n_3305;
wire n_4151;
wire n_4148;
wire n_3528;
wire n_6938;
wire n_4373;
wire n_5762;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_7337;
wire n_6989;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_6427;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_3296;
wire n_2762;
wire n_7038;
wire n_4683;
wire n_5366;
wire n_2767;
wire n_6360;
wire n_2603;
wire n_3116;
wire n_3602;
wire n_2967;
wire n_6146;
wire n_6270;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_5451;
wire n_3923;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_5086;
wire n_2801;
wire n_5901;
wire n_6353;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_3643;
wire n_2825;
wire n_4876;
wire n_6345;
wire n_1997;
wire n_6691;
wire n_3748;
wire n_3142;
wire n_4278;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_7392;
wire n_2215;
wire n_5053;
wire n_6239;
wire n_4553;
wire n_6803;
wire n_3978;
wire n_6340;
wire n_7583;
wire n_4809;
wire n_5226;
wire n_7657;
wire n_1925;
wire n_3660;
wire n_6048;
wire n_5867;
wire n_2491;
wire n_5079;
wire n_5590;
wire n_6773;
wire n_3833;
wire n_5632;
wire n_4841;
wire n_2022;
wire n_6336;
wire n_3814;
wire n_7041;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_7370;
wire n_3513;
wire n_3133;
wire n_5660;
wire n_4645;
wire n_7557;
wire n_2992;
wire n_6174;
wire n_3725;
wire n_4920;
wire n_4972;
wire n_6023;
wire n_2517;
wire n_6776;
wire n_3128;
wire n_5426;
wire n_6463;
wire n_2631;
wire n_2178;
wire n_6372;
wire n_7176;
wire n_2469;
wire n_5625;
wire n_5778;
wire n_6396;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_6669;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_5531;
wire n_3000;
wire n_5429;
wire n_3108;
wire n_3111;
wire n_5818;
wire n_5646;
wire n_6940;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_6394;
wire n_2875;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_7590;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_6995;
wire n_7185;
wire n_3564;
wire n_3988;
wire n_6254;
wire n_6161;
wire n_3457;
wire n_4324;
wire n_4821;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_7332;
wire n_6660;
wire n_4771;
wire n_5719;
wire n_7225;
wire n_6128;
wire n_4086;
wire n_2412;
wire n_7037;
wire n_4814;
wire n_2084;
wire n_3648;
wire n_5749;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_7409;
wire n_4692;
wire n_3031;
wire n_7258;
wire n_7432;
wire n_3701;
wire n_3243;
wire n_6334;
wire n_2666;
wire n_3385;
wire n_6848;
wire n_2171;
wire n_4708;
wire n_6321;
wire n_2768;
wire n_2314;
wire n_6794;
wire n_4826;
wire n_3343;
wire n_2420;
wire n_7197;
wire n_5489;
wire n_6400;
wire n_3767;
wire n_2299;
wire n_2540;
wire n_4589;
wire n_2873;
wire n_5057;
wire n_4578;
wire n_6705;
wire n_2162;
wire n_7619;
wire n_2847;
wire n_2051;
wire n_3221;
wire n_5436;
wire n_5907;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_6044;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_6495;
wire n_5013;
wire n_2312;
wire n_7403;
wire n_6902;
wire n_6470;
wire n_3015;
wire n_5569;
wire n_5439;
wire n_5619;
wire n_4147;
wire n_2048;
wire n_6481;
wire n_3607;
wire n_4925;
wire n_7548;
wire n_6534;
wire n_4974;
wire n_4932;
wire n_4510;
wire n_2571;
wire n_6181;
wire n_3276;
wire n_6728;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_5715;
wire n_6133;
wire n_6528;
wire n_7604;
wire n_7407;
wire n_3827;
wire n_3354;
wire n_2519;
wire n_2724;
wire n_4447;
wire n_6670;
wire n_6774;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_6741;
wire n_7424;
wire n_6038;
wire n_4818;
wire n_4514;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_6282;
wire n_2110;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_6700;
wire n_7334;
wire n_2033;
wire n_7684;
wire n_4341;
wire n_4312;
wire n_3399;
wire n_2628;
wire n_5932;
wire n_6178;
wire n_2132;
wire n_6234;
wire n_6012;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_3387;
wire n_5186;
wire n_7367;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_6715;
wire n_5828;
wire n_2831;
wire n_7200;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_7582;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_3037;
wire n_6337;
wire n_4868;
wire n_2452;
wire n_6770;
wire n_6743;
wire n_3925;
wire n_2176;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_6682;
wire n_5054;
wire n_7673;
wire n_5631;
wire n_2467;
wire n_6539;
wire n_7243;
wire n_7179;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_6314;
wire n_6617;
wire n_3592;
wire n_5694;
wire n_4650;
wire n_4888;
wire n_7274;
wire n_5326;
wire n_3394;
wire n_4874;
wire n_7608;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_6595;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_4060;
wire n_2658;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_6385;
wire n_6289;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_4796;
wire n_7373;
wire n_3589;
wire n_2534;
wire n_6186;
wire n_4799;
wire n_5153;
wire n_6257;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_6852;
wire n_2789;
wire n_6346;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_5809;
wire n_5365;
wire n_2933;
wire n_7587;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_6274;
wire n_7372;
wire n_2328;
wire n_4248;
wire n_5915;
wire n_6818;
wire n_5452;
wire n_7226;
wire n_4754;
wire n_7057;
wire n_7685;
wire n_4554;
wire n_5595;
wire n_6609;
wire n_4845;
wire n_6753;
wire n_6815;
wire n_3053;
wire n_3893;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_6764;
wire n_5535;
wire n_3875;
wire n_5370;
wire n_6391;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_5594;
wire n_4301;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_6471;
wire n_3777;
wire n_6627;
wire n_5761;
wire n_4784;
wire n_7203;
wire n_2999;
wire n_7512;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_7215;
wire n_3080;
wire n_6636;
wire n_4199;
wire n_2701;
wire n_5929;
wire n_3362;
wire n_5559;
wire n_3105;
wire n_5478;
wire n_7388;
wire n_6243;
wire n_6488;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_6022;
wire n_6457;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_3913;
wire n_6867;
wire n_3417;
wire n_5868;
wire n_6230;
wire n_4034;
wire n_6538;
wire n_6633;
wire n_6187;
wire n_3327;
wire n_6172;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_7311;
wire n_2755;
wire n_5989;
wire n_3237;
wire n_6574;
wire n_1992;
wire n_6395;
wire n_4402;
wire n_4239;
wire n_6854;
wire n_3400;
wire n_6233;
wire n_4550;
wire n_6456;
wire n_3382;
wire n_7488;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_7198;
wire n_4201;
wire n_6784;
wire n_6168;
wire n_3316;
wire n_6766;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_3603;
wire n_4123;
wire n_6330;
wire n_2192;
wire n_5520;
wire n_3633;
wire n_4479;
wire n_7249;
wire n_2670;
wire n_5947;
wire n_7336;
wire n_4416;
wire n_3372;
wire n_7031;
wire n_4539;
wire n_2707;
wire n_6799;
wire n_5920;
wire n_6672;
wire n_2471;
wire n_6149;
wire n_7142;
wire n_3230;
wire n_5808;
wire n_3342;
wire n_6054;
wire n_7089;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_6450;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_7042;
wire n_3780;
wire n_1928;
wire n_5244;
wire n_6523;
wire n_5382;
wire n_6107;
wire n_3957;
wire n_6775;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_6232;
wire n_6445;
wire n_7181;
wire n_6134;
wire n_5384;
wire n_3608;
wire n_6056;
wire n_6932;
wire n_7036;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_5587;
wire n_2619;
wire n_6855;
wire n_2444;
wire n_5789;
wire n_3123;
wire n_5787;
wire n_6585;
wire n_6369;
wire n_5056;
wire n_5249;
wire n_3393;
wire n_7447;
wire n_5198;
wire n_5360;
wire n_7455;
wire n_5233;
wire n_4887;
wire n_5829;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_6252;
wire n_5866;
wire n_6493;
wire n_4005;
wire n_4904;
wire n_5899;
wire n_7629;
wire n_4792;
wire n_7104;
wire n_3578;
wire n_3812;
wire n_7601;
wire n_4980;
wire n_6026;
wire n_4290;
wire n_5247;
wire n_5865;
wire n_3727;
wire n_5317;
wire n_6544;
wire n_3774;
wire n_3093;
wire n_3061;
wire n_7138;
wire n_7290;
wire n_2431;
wire n_6679;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_5924;
wire n_3182;
wire n_7625;
wire n_5822;
wire n_2564;
wire n_6259;
wire n_4947;
wire n_7284;
wire n_4656;
wire n_3896;
wire n_3958;
wire n_6390;
wire n_3450;
wire n_4729;
wire n_5786;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_2000;
wire n_2074;
wire n_3174;
wire n_2217;
wire n_6630;
wire n_3398;
wire n_5658;
wire n_2307;
wire n_3408;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_3432;
wire n_6279;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_6813;
wire n_5564;
wire n_2445;
wire n_1988;
wire n_7106;
wire n_6042;
wire n_7644;
wire n_6057;
wire n_4137;
wire n_7529;
wire n_6675;
wire n_2634;
wire n_4529;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_6476;
wire n_3972;
wire n_6207;
wire n_5539;
wire n_6268;
wire n_6878;
wire n_6286;
wire n_3308;
wire n_6524;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_6225;
wire n_4322;
wire n_7297;
wire n_6291;
wire n_2830;
wire n_5893;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_7199;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_5261;
wire n_6520;
wire n_7648;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_2245;
wire n_4909;
wire n_2965;
wire n_3635;
wire n_6024;
wire n_5022;
wire n_5005;
wire n_2814;
wire n_3882;
wire n_3046;
wire n_7487;
wire n_2213;
wire n_6425;
wire n_5993;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_7638;
wire n_5703;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_6432;
wire n_5534;
wire n_3204;
wire n_7259;
wire n_2136;
wire n_6540;
wire n_6955;
wire n_5174;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_4380;
wire n_3129;
wire n_4126;
wire n_7237;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_6388;
wire n_5904;
wire n_4880;
wire n_6760;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_5061;
wire n_5572;
wire n_5750;
wire n_7063;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_7576;
wire n_3023;
wire n_6795;
wire n_5881;
wire n_6664;
wire n_5815;
wire n_6261;
wire n_4193;
wire n_5873;
wire n_4075;
wire n_3104;
wire n_6487;
wire n_4737;
wire n_6729;
wire n_3647;
wire n_5755;
wire n_2819;
wire n_5949;
wire n_5195;
wire n_7483;
wire n_3609;
wire n_4136;
wire n_6608;
wire n_1952;
wire n_4393;
wire n_7385;
wire n_3720;
wire n_4535;
wire n_7668;
wire n_2560;
wire n_4522;
wire n_6663;
wire n_4794;
wire n_5955;
wire n_7476;
wire n_3959;
wire n_7327;
wire n_5763;
wire n_6656;
wire n_6843;
wire n_3140;
wire n_5246;
wire n_5964;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_7266;
wire n_5164;
wire n_4196;
wire n_6969;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_5665;
wire n_6485;
wire n_3069;
wire n_5498;
wire n_7100;
wire n_4370;
wire n_5783;
wire n_5183;
wire n_6075;
wire n_7082;
wire n_3084;
wire n_6120;
wire n_6659;
wire n_2735;
wire n_6750;
wire n_3412;
wire n_2497;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_3761;
wire n_4889;
wire n_7132;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_5739;
wire n_3184;
wire n_4828;
wire n_6003;
wire n_5385;
wire n_4558;
wire n_6478;
wire n_2172;
wire n_6066;
wire n_7034;
wire n_6086;
wire n_4722;
wire n_6650;
wire n_6224;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_2250;
wire n_7084;
wire n_5845;
wire n_7293;
wire n_4092;
wire n_5990;
wire n_3908;
wire n_6175;
wire n_6060;
wire n_7253;
wire n_2423;
wire n_3671;
wire n_6891;
wire n_5663;
wire n_6410;
wire n_3344;
wire n_2194;
wire n_4465;
wire n_5973;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_2680;
wire n_6059;
wire n_5130;
wire n_7520;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_6103;
wire n_6809;
wire n_3265;
wire n_4482;
wire n_2041;
wire n_6267;
wire n_2957;
wire n_5855;
wire n_2357;
wire n_5757;
wire n_6437;
wire n_3309;
wire n_7331;
wire n_6610;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_4116;
wire n_6957;
wire n_5704;
wire n_7514;
wire n_7163;
wire n_7620;
wire n_2570;
wire n_2815;
wire n_5473;
wire n_3754;
wire n_4612;
wire n_5946;
wire n_2744;
wire n_6711;
wire n_4287;
wire n_2397;
wire n_7445;
wire n_2208;
wire n_6847;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_7123;
wire n_6384;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_7563;
wire n_6298;
wire n_2591;
wire n_3384;
wire n_7361;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_7322;
wire n_5710;
wire n_7453;
wire n_6067;
wire n_5070;
wire n_6377;
wire n_4445;
wire n_5566;
wire n_5414;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_6348;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_6129;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_6834;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_6136;
wire n_7261;
wire n_6723;
wire n_5834;
wire n_2823;
wire n_5874;
wire n_7508;
wire n_7021;
wire n_5270;
wire n_5956;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_6078;
wire n_7000;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_7130;
wire n_5823;
wire n_3997;
wire n_5465;
wire n_4032;
wire n_3582;
wire n_7538;
wire n_7517;
wire n_5853;
wire n_2826;
wire n_3539;
wire n_7077;
wire n_4343;
wire n_4212;
wire n_6642;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_7346;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_7333;
wire n_4364;
wire n_4245;
wire n_4928;
wire n_2225;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_7546;
wire n_3853;
wire n_4216;
wire n_5934;
wire n_6942;
wire n_2019;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_6511;
wire n_3721;
wire n_6507;
wire n_2026;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_2614;
wire n_7319;
wire n_2991;
wire n_6497;
wire n_6001;
wire n_6007;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_6606;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_5395;
wire n_2237;
wire n_7078;
wire n_3463;
wire n_7047;
wire n_3699;
wire n_5067;
wire n_7107;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_7469;
wire n_3857;
wire n_2728;

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1785),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1707),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_512),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1502),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1303),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_160),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_1803),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_903),
.Y(n_1931)
);

INVx2_ASAP7_75t_SL g1932 ( 
.A(n_1374),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1709),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_460),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1672),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_122),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_966),
.Y(n_1937)
);

BUFx5_ASAP7_75t_L g1938 ( 
.A(n_1037),
.Y(n_1938)
);

CKINVDCx20_ASAP7_75t_R g1939 ( 
.A(n_495),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1476),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_227),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_488),
.Y(n_1942)
);

CKINVDCx14_ASAP7_75t_R g1943 ( 
.A(n_10),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_852),
.Y(n_1944)
);

BUFx6f_ASAP7_75t_L g1945 ( 
.A(n_470),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1586),
.Y(n_1946)
);

CKINVDCx20_ASAP7_75t_R g1947 ( 
.A(n_264),
.Y(n_1947)
);

CKINVDCx20_ASAP7_75t_R g1948 ( 
.A(n_275),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1897),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_490),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1220),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1250),
.Y(n_1952)
);

CKINVDCx16_ASAP7_75t_R g1953 ( 
.A(n_974),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1906),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_944),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1058),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1877),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_409),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_263),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_46),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1429),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_57),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1757),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1805),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_323),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_1457),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1526),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_724),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1499),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_162),
.Y(n_1970)
);

CKINVDCx20_ASAP7_75t_R g1971 ( 
.A(n_1537),
.Y(n_1971)
);

CKINVDCx20_ASAP7_75t_R g1972 ( 
.A(n_598),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1775),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_91),
.Y(n_1974)
);

BUFx6f_ASAP7_75t_L g1975 ( 
.A(n_1627),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1272),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_962),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1864),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1244),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_880),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_478),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_670),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_644),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1721),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_676),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_801),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_555),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_1696),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_1712),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1593),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_30),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1797),
.Y(n_1992)
);

INVx1_ASAP7_75t_SL g1993 ( 
.A(n_1026),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1341),
.Y(n_1994)
);

BUFx2_ASAP7_75t_SL g1995 ( 
.A(n_742),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1387),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1233),
.Y(n_1997)
);

INVxp67_ASAP7_75t_SL g1998 ( 
.A(n_865),
.Y(n_1998)
);

INVx1_ASAP7_75t_SL g1999 ( 
.A(n_1301),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1751),
.Y(n_2000)
);

CKINVDCx20_ASAP7_75t_R g2001 ( 
.A(n_44),
.Y(n_2001)
);

BUFx2_ASAP7_75t_SL g2002 ( 
.A(n_1802),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1649),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_39),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1425),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1830),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1108),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1685),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1624),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1875),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1913),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_896),
.Y(n_2012)
);

BUFx3_ASAP7_75t_L g2013 ( 
.A(n_631),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_603),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_169),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1736),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1114),
.Y(n_2017)
);

CKINVDCx20_ASAP7_75t_R g2018 ( 
.A(n_443),
.Y(n_2018)
);

BUFx6f_ASAP7_75t_L g2019 ( 
.A(n_1574),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1292),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1631),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_845),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1237),
.Y(n_2023)
);

BUFx6f_ASAP7_75t_L g2024 ( 
.A(n_1703),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1691),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_614),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_332),
.Y(n_2027)
);

CKINVDCx20_ASAP7_75t_R g2028 ( 
.A(n_1823),
.Y(n_2028)
);

CKINVDCx20_ASAP7_75t_R g2029 ( 
.A(n_398),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_SL g2030 ( 
.A(n_1588),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1143),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1069),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1637),
.Y(n_2033)
);

INVx4_ASAP7_75t_R g2034 ( 
.A(n_234),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1299),
.Y(n_2035)
);

CKINVDCx20_ASAP7_75t_R g2036 ( 
.A(n_1722),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1613),
.Y(n_2037)
);

CKINVDCx16_ASAP7_75t_R g2038 ( 
.A(n_239),
.Y(n_2038)
);

BUFx3_ASAP7_75t_L g2039 ( 
.A(n_134),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_101),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1756),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_937),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1170),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_1768),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_208),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1518),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1219),
.Y(n_2047)
);

INVx2_ASAP7_75t_SL g2048 ( 
.A(n_1175),
.Y(n_2048)
);

CKINVDCx20_ASAP7_75t_R g2049 ( 
.A(n_960),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_773),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_199),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1908),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1415),
.Y(n_2053)
);

BUFx5_ASAP7_75t_L g2054 ( 
.A(n_1598),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_619),
.Y(n_2055)
);

CKINVDCx5p33_ASAP7_75t_R g2056 ( 
.A(n_1663),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_812),
.Y(n_2057)
);

BUFx2_ASAP7_75t_L g2058 ( 
.A(n_1732),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_31),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_177),
.Y(n_2060)
);

CKINVDCx20_ASAP7_75t_R g2061 ( 
.A(n_616),
.Y(n_2061)
);

CKINVDCx20_ASAP7_75t_R g2062 ( 
.A(n_1138),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1559),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_1451),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1670),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1915),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1563),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_774),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1800),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_696),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_475),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_1889),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_582),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1827),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1792),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1249),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_1417),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_813),
.Y(n_2078)
);

CKINVDCx20_ASAP7_75t_R g2079 ( 
.A(n_613),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1790),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1312),
.Y(n_2081)
);

BUFx3_ASAP7_75t_L g2082 ( 
.A(n_1911),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1494),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_34),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1687),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_829),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_1509),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1719),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_179),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_857),
.Y(n_2090)
);

INVx1_ASAP7_75t_SL g2091 ( 
.A(n_1921),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1005),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1857),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1435),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_393),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_504),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1887),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_401),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_900),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1434),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_1920),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_265),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1391),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_410),
.Y(n_2104)
);

CKINVDCx16_ASAP7_75t_R g2105 ( 
.A(n_477),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1227),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1383),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_611),
.Y(n_2108)
);

BUFx10_ASAP7_75t_L g2109 ( 
.A(n_1717),
.Y(n_2109)
);

CKINVDCx20_ASAP7_75t_R g2110 ( 
.A(n_1539),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1755),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_1261),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1680),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_154),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_278),
.Y(n_2115)
);

CKINVDCx20_ASAP7_75t_R g2116 ( 
.A(n_1308),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1584),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_401),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1738),
.Y(n_2119)
);

CKINVDCx16_ASAP7_75t_R g2120 ( 
.A(n_1490),
.Y(n_2120)
);

CKINVDCx16_ASAP7_75t_R g2121 ( 
.A(n_893),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_155),
.Y(n_2122)
);

CKINVDCx20_ASAP7_75t_R g2123 ( 
.A(n_15),
.Y(n_2123)
);

CKINVDCx20_ASAP7_75t_R g2124 ( 
.A(n_888),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1506),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_462),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1873),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1335),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_1104),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1798),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_1757),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_14),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1788),
.Y(n_2133)
);

INVx1_ASAP7_75t_SL g2134 ( 
.A(n_1643),
.Y(n_2134)
);

CKINVDCx16_ASAP7_75t_R g2135 ( 
.A(n_1736),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_164),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_572),
.Y(n_2137)
);

INVx2_ASAP7_75t_SL g2138 ( 
.A(n_1746),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_669),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_456),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1790),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_1590),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_887),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1103),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_1008),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_752),
.Y(n_2146)
);

CKINVDCx20_ASAP7_75t_R g2147 ( 
.A(n_1161),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_921),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_492),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_301),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1316),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_24),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_446),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_543),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_82),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_1763),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_1639),
.Y(n_2157)
);

INVx1_ASAP7_75t_SL g2158 ( 
.A(n_1712),
.Y(n_2158)
);

BUFx2_ASAP7_75t_L g2159 ( 
.A(n_737),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_1302),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_320),
.Y(n_2161)
);

BUFx10_ASAP7_75t_L g2162 ( 
.A(n_1287),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_754),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_196),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_830),
.Y(n_2165)
);

CKINVDCx5p33_ASAP7_75t_R g2166 ( 
.A(n_1629),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_1555),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_670),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_1513),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_1010),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_90),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_1507),
.Y(n_2172)
);

BUFx2_ASAP7_75t_SL g2173 ( 
.A(n_965),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1764),
.Y(n_2174)
);

CKINVDCx16_ASAP7_75t_R g2175 ( 
.A(n_858),
.Y(n_2175)
);

BUFx3_ASAP7_75t_L g2176 ( 
.A(n_506),
.Y(n_2176)
);

BUFx10_ASAP7_75t_L g2177 ( 
.A(n_280),
.Y(n_2177)
);

CKINVDCx5p33_ASAP7_75t_R g2178 ( 
.A(n_1265),
.Y(n_2178)
);

INVx2_ASAP7_75t_SL g2179 ( 
.A(n_1316),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_643),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_651),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_1723),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1721),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_215),
.Y(n_2184)
);

CKINVDCx16_ASAP7_75t_R g2185 ( 
.A(n_1413),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1795),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_1648),
.Y(n_2187)
);

BUFx6f_ASAP7_75t_L g2188 ( 
.A(n_1744),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_14),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_241),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_121),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_499),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_1759),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_209),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_968),
.Y(n_2195)
);

CKINVDCx5p33_ASAP7_75t_R g2196 ( 
.A(n_32),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_479),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_408),
.Y(n_2198)
);

INVx1_ASAP7_75t_SL g2199 ( 
.A(n_25),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_1149),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_572),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_259),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_326),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_1539),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_782),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1633),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_1112),
.Y(n_2208)
);

BUFx3_ASAP7_75t_L g2209 ( 
.A(n_1080),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_606),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1570),
.Y(n_2211)
);

BUFx10_ASAP7_75t_L g2212 ( 
.A(n_262),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_545),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_565),
.Y(n_2214)
);

INVx1_ASAP7_75t_SL g2215 ( 
.A(n_903),
.Y(n_2215)
);

BUFx3_ASAP7_75t_L g2216 ( 
.A(n_1190),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_429),
.Y(n_2217)
);

CKINVDCx20_ASAP7_75t_R g2218 ( 
.A(n_852),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_1458),
.Y(n_2219)
);

BUFx10_ASAP7_75t_L g2220 ( 
.A(n_559),
.Y(n_2220)
);

CKINVDCx20_ASAP7_75t_R g2221 ( 
.A(n_666),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_1718),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_733),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_245),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_1064),
.Y(n_2225)
);

CKINVDCx14_ASAP7_75t_R g2226 ( 
.A(n_1682),
.Y(n_2226)
);

CKINVDCx20_ASAP7_75t_R g2227 ( 
.A(n_359),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_677),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1829),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_28),
.Y(n_2230)
);

CKINVDCx20_ASAP7_75t_R g2231 ( 
.A(n_1333),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_1105),
.Y(n_2232)
);

CKINVDCx20_ASAP7_75t_R g2233 ( 
.A(n_1391),
.Y(n_2233)
);

CKINVDCx20_ASAP7_75t_R g2234 ( 
.A(n_1778),
.Y(n_2234)
);

CKINVDCx14_ASAP7_75t_R g2235 ( 
.A(n_1789),
.Y(n_2235)
);

CKINVDCx16_ASAP7_75t_R g2236 ( 
.A(n_600),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_1677),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_1401),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_892),
.Y(n_2239)
);

BUFx6f_ASAP7_75t_L g2240 ( 
.A(n_301),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1710),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_432),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_1656),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_487),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_L g2245 ( 
.A(n_747),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_195),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1825),
.Y(n_2247)
);

INVx2_ASAP7_75t_SL g2248 ( 
.A(n_1294),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1311),
.Y(n_2249)
);

BUFx8_ASAP7_75t_SL g2250 ( 
.A(n_1619),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_943),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_1730),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_665),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1384),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_829),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_643),
.Y(n_2256)
);

INVx2_ASAP7_75t_SL g2257 ( 
.A(n_942),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_1212),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_672),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_594),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_1550),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_1106),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1551),
.Y(n_2263)
);

INVx2_ASAP7_75t_SL g2264 ( 
.A(n_1589),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1733),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_640),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_193),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_859),
.Y(n_2268)
);

CKINVDCx5p33_ASAP7_75t_R g2269 ( 
.A(n_1503),
.Y(n_2269)
);

CKINVDCx5p33_ASAP7_75t_R g2270 ( 
.A(n_969),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1659),
.Y(n_2271)
);

HB1xp67_ASAP7_75t_L g2272 ( 
.A(n_297),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_4),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1401),
.Y(n_2274)
);

BUFx6f_ASAP7_75t_L g2275 ( 
.A(n_1660),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_1227),
.Y(n_2276)
);

BUFx10_ASAP7_75t_L g2277 ( 
.A(n_1705),
.Y(n_2277)
);

CKINVDCx5p33_ASAP7_75t_R g2278 ( 
.A(n_1618),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_203),
.Y(n_2279)
);

BUFx3_ASAP7_75t_L g2280 ( 
.A(n_1601),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_19),
.Y(n_2281)
);

CKINVDCx5p33_ASAP7_75t_R g2282 ( 
.A(n_1427),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_434),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_1797),
.Y(n_2284)
);

INVx1_ASAP7_75t_SL g2285 ( 
.A(n_925),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_977),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_810),
.Y(n_2287)
);

CKINVDCx20_ASAP7_75t_R g2288 ( 
.A(n_1221),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_727),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_223),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_989),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_1728),
.Y(n_2292)
);

CKINVDCx20_ASAP7_75t_R g2293 ( 
.A(n_1922),
.Y(n_2293)
);

CKINVDCx5p33_ASAP7_75t_R g2294 ( 
.A(n_1655),
.Y(n_2294)
);

BUFx3_ASAP7_75t_L g2295 ( 
.A(n_1657),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1654),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_22),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_503),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1674),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_1784),
.Y(n_2300)
);

HB1xp67_ASAP7_75t_L g2301 ( 
.A(n_1796),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_1146),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_1340),
.Y(n_2303)
);

CKINVDCx5p33_ASAP7_75t_R g2304 ( 
.A(n_1371),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_526),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_827),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_809),
.Y(n_2307)
);

INVx1_ASAP7_75t_SL g2308 ( 
.A(n_138),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_527),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1344),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_438),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_502),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1918),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_1200),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_409),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_91),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_429),
.Y(n_2317)
);

CKINVDCx5p33_ASAP7_75t_R g2318 ( 
.A(n_1641),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1554),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_835),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_1739),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1632),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_523),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_1623),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_209),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_394),
.Y(n_2326)
);

CKINVDCx5p33_ASAP7_75t_R g2327 ( 
.A(n_368),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_1530),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_78),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_1139),
.Y(n_2330)
);

CKINVDCx5p33_ASAP7_75t_R g2331 ( 
.A(n_1907),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1672),
.Y(n_2332)
);

CKINVDCx14_ASAP7_75t_R g2333 ( 
.A(n_664),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_1680),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1169),
.Y(n_2335)
);

CKINVDCx14_ASAP7_75t_R g2336 ( 
.A(n_931),
.Y(n_2336)
);

CKINVDCx5p33_ASAP7_75t_R g2337 ( 
.A(n_806),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1020),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_397),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_1683),
.Y(n_2340)
);

INVx1_ASAP7_75t_SL g2341 ( 
.A(n_1695),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_586),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_967),
.Y(n_2343)
);

CKINVDCx5p33_ASAP7_75t_R g2344 ( 
.A(n_947),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_1268),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_482),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_258),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_789),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_1917),
.Y(n_2349)
);

CKINVDCx16_ASAP7_75t_R g2350 ( 
.A(n_445),
.Y(n_2350)
);

INVx1_ASAP7_75t_SL g2351 ( 
.A(n_1163),
.Y(n_2351)
);

CKINVDCx5p33_ASAP7_75t_R g2352 ( 
.A(n_1780),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1660),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_1765),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_1904),
.Y(n_2355)
);

CKINVDCx20_ASAP7_75t_R g2356 ( 
.A(n_1448),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_129),
.Y(n_2357)
);

INVxp67_ASAP7_75t_L g2358 ( 
.A(n_1441),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_105),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_702),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_714),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_930),
.Y(n_2362)
);

CKINVDCx20_ASAP7_75t_R g2363 ( 
.A(n_1874),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_711),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_150),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_888),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1551),
.Y(n_2367)
);

CKINVDCx5p33_ASAP7_75t_R g2368 ( 
.A(n_838),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_624),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_1049),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_432),
.Y(n_2371)
);

CKINVDCx5p33_ASAP7_75t_R g2372 ( 
.A(n_1358),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_1741),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1762),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_157),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_1619),
.Y(n_2376)
);

CKINVDCx20_ASAP7_75t_R g2377 ( 
.A(n_99),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_1437),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_1615),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_636),
.Y(n_2380)
);

CKINVDCx5p33_ASAP7_75t_R g2381 ( 
.A(n_578),
.Y(n_2381)
);

CKINVDCx20_ASAP7_75t_R g2382 ( 
.A(n_1096),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1252),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_1822),
.Y(n_2384)
);

CKINVDCx5p33_ASAP7_75t_R g2385 ( 
.A(n_1146),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_493),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_815),
.Y(n_2387)
);

CKINVDCx20_ASAP7_75t_R g2388 ( 
.A(n_1676),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_1711),
.Y(n_2389)
);

INVx1_ASAP7_75t_SL g2390 ( 
.A(n_221),
.Y(n_2390)
);

INVxp67_ASAP7_75t_L g2391 ( 
.A(n_1064),
.Y(n_2391)
);

BUFx3_ASAP7_75t_L g2392 ( 
.A(n_907),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_1713),
.Y(n_2393)
);

BUFx3_ASAP7_75t_L g2394 ( 
.A(n_1811),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_865),
.Y(n_2395)
);

INVx1_ASAP7_75t_SL g2396 ( 
.A(n_1017),
.Y(n_2396)
);

INVx2_ASAP7_75t_SL g2397 ( 
.A(n_1175),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_1295),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_L g2399 ( 
.A(n_263),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_1169),
.Y(n_2400)
);

CKINVDCx20_ASAP7_75t_R g2401 ( 
.A(n_962),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_1303),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_1642),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_1506),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_754),
.Y(n_2405)
);

CKINVDCx5p33_ASAP7_75t_R g2406 ( 
.A(n_1474),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_742),
.Y(n_2407)
);

CKINVDCx5p33_ASAP7_75t_R g2408 ( 
.A(n_1701),
.Y(n_2408)
);

CKINVDCx16_ASAP7_75t_R g2409 ( 
.A(n_1870),
.Y(n_2409)
);

CKINVDCx5p33_ASAP7_75t_R g2410 ( 
.A(n_80),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1411),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_69),
.Y(n_2412)
);

CKINVDCx5p33_ASAP7_75t_R g2413 ( 
.A(n_266),
.Y(n_2413)
);

BUFx6f_ASAP7_75t_L g2414 ( 
.A(n_890),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_1831),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1653),
.Y(n_2416)
);

BUFx2_ASAP7_75t_L g2417 ( 
.A(n_1471),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_1249),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_1919),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_102),
.Y(n_2420)
);

BUFx10_ASAP7_75t_L g2421 ( 
.A(n_284),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_1299),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_41),
.Y(n_2423)
);

CKINVDCx5p33_ASAP7_75t_R g2424 ( 
.A(n_1260),
.Y(n_2424)
);

HB1xp67_ASAP7_75t_L g2425 ( 
.A(n_1794),
.Y(n_2425)
);

INVx1_ASAP7_75t_SL g2426 ( 
.A(n_1774),
.Y(n_2426)
);

BUFx10_ASAP7_75t_L g2427 ( 
.A(n_1914),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_1620),
.Y(n_2428)
);

CKINVDCx20_ASAP7_75t_R g2429 ( 
.A(n_1766),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_1662),
.Y(n_2430)
);

CKINVDCx5p33_ASAP7_75t_R g2431 ( 
.A(n_90),
.Y(n_2431)
);

CKINVDCx5p33_ASAP7_75t_R g2432 ( 
.A(n_188),
.Y(n_2432)
);

INVx1_ASAP7_75t_SL g2433 ( 
.A(n_1668),
.Y(n_2433)
);

CKINVDCx5p33_ASAP7_75t_R g2434 ( 
.A(n_701),
.Y(n_2434)
);

CKINVDCx16_ASAP7_75t_R g2435 ( 
.A(n_1802),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_321),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_483),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1795),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_816),
.Y(n_2439)
);

BUFx2_ASAP7_75t_L g2440 ( 
.A(n_1690),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_1071),
.Y(n_2441)
);

CKINVDCx5p33_ASAP7_75t_R g2442 ( 
.A(n_1315),
.Y(n_2442)
);

INVx1_ASAP7_75t_SL g2443 ( 
.A(n_570),
.Y(n_2443)
);

INVx1_ASAP7_75t_SL g2444 ( 
.A(n_1379),
.Y(n_2444)
);

INVx2_ASAP7_75t_SL g2445 ( 
.A(n_1812),
.Y(n_2445)
);

BUFx6f_ASAP7_75t_L g2446 ( 
.A(n_1695),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_7),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_1503),
.Y(n_2448)
);

CKINVDCx5p33_ASAP7_75t_R g2449 ( 
.A(n_375),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_633),
.Y(n_2450)
);

CKINVDCx20_ASAP7_75t_R g2451 ( 
.A(n_1637),
.Y(n_2451)
);

BUFx6f_ASAP7_75t_L g2452 ( 
.A(n_782),
.Y(n_2452)
);

INVx1_ASAP7_75t_SL g2453 ( 
.A(n_688),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_21),
.Y(n_2454)
);

HB1xp67_ASAP7_75t_L g2455 ( 
.A(n_1468),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_1362),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_1258),
.Y(n_2457)
);

CKINVDCx5p33_ASAP7_75t_R g2458 ( 
.A(n_564),
.Y(n_2458)
);

CKINVDCx5p33_ASAP7_75t_R g2459 ( 
.A(n_764),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_1510),
.Y(n_2460)
);

INVx1_ASAP7_75t_SL g2461 ( 
.A(n_981),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_1107),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_319),
.Y(n_2463)
);

INVx2_ASAP7_75t_SL g2464 ( 
.A(n_1792),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_98),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_1626),
.Y(n_2466)
);

INVxp67_ASAP7_75t_L g2467 ( 
.A(n_318),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_1791),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_159),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_1923),
.Y(n_2470)
);

CKINVDCx20_ASAP7_75t_R g2471 ( 
.A(n_317),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_1675),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1304),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_391),
.Y(n_2474)
);

BUFx10_ASAP7_75t_L g2475 ( 
.A(n_1773),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_302),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_691),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_1611),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_890),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_1252),
.Y(n_2480)
);

CKINVDCx5p33_ASAP7_75t_R g2481 ( 
.A(n_282),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_632),
.Y(n_2482)
);

INVx1_ASAP7_75t_SL g2483 ( 
.A(n_259),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_128),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_1731),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_637),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_1681),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_873),
.Y(n_2488)
);

BUFx5_ASAP7_75t_L g2489 ( 
.A(n_1120),
.Y(n_2489)
);

INVx2_ASAP7_75t_SL g2490 ( 
.A(n_1060),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_1364),
.Y(n_2491)
);

CKINVDCx5p33_ASAP7_75t_R g2492 ( 
.A(n_336),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_334),
.Y(n_2493)
);

CKINVDCx5p33_ASAP7_75t_R g2494 ( 
.A(n_1351),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_1731),
.Y(n_2495)
);

CKINVDCx16_ASAP7_75t_R g2496 ( 
.A(n_1258),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_1073),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_368),
.Y(n_2498)
);

CKINVDCx5p33_ASAP7_75t_R g2499 ( 
.A(n_148),
.Y(n_2499)
);

CKINVDCx5p33_ASAP7_75t_R g2500 ( 
.A(n_1666),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_812),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_1494),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_631),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_1785),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_1854),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_35),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_710),
.Y(n_2507)
);

CKINVDCx5p33_ASAP7_75t_R g2508 ( 
.A(n_874),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_1678),
.Y(n_2509)
);

CKINVDCx5p33_ASAP7_75t_R g2510 ( 
.A(n_1142),
.Y(n_2510)
);

CKINVDCx5p33_ASAP7_75t_R g2511 ( 
.A(n_1020),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_1224),
.Y(n_2512)
);

CKINVDCx20_ASAP7_75t_R g2513 ( 
.A(n_482),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_1027),
.Y(n_2514)
);

CKINVDCx20_ASAP7_75t_R g2515 ( 
.A(n_1443),
.Y(n_2515)
);

BUFx2_ASAP7_75t_L g2516 ( 
.A(n_1807),
.Y(n_2516)
);

CKINVDCx20_ASAP7_75t_R g2517 ( 
.A(n_1758),
.Y(n_2517)
);

INVxp67_ASAP7_75t_L g2518 ( 
.A(n_690),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_1592),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_707),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_303),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_564),
.Y(n_2522)
);

CKINVDCx5p33_ASAP7_75t_R g2523 ( 
.A(n_1708),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_949),
.Y(n_2524)
);

INVx2_ASAP7_75t_SL g2525 ( 
.A(n_1650),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_1240),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_611),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_1220),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_1603),
.Y(n_2529)
);

CKINVDCx5p33_ASAP7_75t_R g2530 ( 
.A(n_1692),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_1241),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_344),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_82),
.Y(n_2533)
);

CKINVDCx5p33_ASAP7_75t_R g2534 ( 
.A(n_1118),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_950),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_703),
.Y(n_2536)
);

BUFx6f_ASAP7_75t_L g2537 ( 
.A(n_795),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_1418),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_915),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_1184),
.Y(n_2540)
);

CKINVDCx16_ASAP7_75t_R g2541 ( 
.A(n_510),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_302),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_128),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_867),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_1652),
.Y(n_2545)
);

CKINVDCx5p33_ASAP7_75t_R g2546 ( 
.A(n_264),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_623),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_1661),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_1034),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_1124),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_879),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_503),
.Y(n_2552)
);

CKINVDCx5p33_ASAP7_75t_R g2553 ( 
.A(n_1916),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_975),
.Y(n_2554)
);

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_1745),
.Y(n_2555)
);

INVx1_ASAP7_75t_SL g2556 ( 
.A(n_1748),
.Y(n_2556)
);

BUFx6f_ASAP7_75t_L g2557 ( 
.A(n_945),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_1653),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_877),
.Y(n_2559)
);

CKINVDCx5p33_ASAP7_75t_R g2560 ( 
.A(n_1479),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_1625),
.Y(n_2561)
);

CKINVDCx5p33_ASAP7_75t_R g2562 ( 
.A(n_578),
.Y(n_2562)
);

CKINVDCx20_ASAP7_75t_R g2563 ( 
.A(n_935),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_950),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_1749),
.Y(n_2565)
);

CKINVDCx5p33_ASAP7_75t_R g2566 ( 
.A(n_1694),
.Y(n_2566)
);

BUFx2_ASAP7_75t_L g2567 ( 
.A(n_722),
.Y(n_2567)
);

CKINVDCx5p33_ASAP7_75t_R g2568 ( 
.A(n_1595),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_309),
.Y(n_2569)
);

CKINVDCx5p33_ASAP7_75t_R g2570 ( 
.A(n_1697),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_222),
.Y(n_2571)
);

BUFx3_ASAP7_75t_L g2572 ( 
.A(n_219),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_837),
.Y(n_2573)
);

INVx1_ASAP7_75t_SL g2574 ( 
.A(n_1479),
.Y(n_2574)
);

CKINVDCx20_ASAP7_75t_R g2575 ( 
.A(n_1437),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_1777),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_1467),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_504),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_1086),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_1729),
.Y(n_2580)
);

CKINVDCx5p33_ASAP7_75t_R g2581 ( 
.A(n_526),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_686),
.Y(n_2582)
);

CKINVDCx5p33_ASAP7_75t_R g2583 ( 
.A(n_535),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_990),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_1535),
.Y(n_2585)
);

CKINVDCx5p33_ASAP7_75t_R g2586 ( 
.A(n_1257),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_1123),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_1651),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_1593),
.Y(n_2589)
);

CKINVDCx5p33_ASAP7_75t_R g2590 ( 
.A(n_1718),
.Y(n_2590)
);

CKINVDCx5p33_ASAP7_75t_R g2591 ( 
.A(n_1029),
.Y(n_2591)
);

BUFx6f_ASAP7_75t_L g2592 ( 
.A(n_1314),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_464),
.Y(n_2593)
);

BUFx10_ASAP7_75t_L g2594 ( 
.A(n_1684),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_1772),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_396),
.Y(n_2596)
);

INVx1_ASAP7_75t_SL g2597 ( 
.A(n_644),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_1090),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_592),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_1344),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_333),
.Y(n_2601)
);

CKINVDCx5p33_ASAP7_75t_R g2602 ( 
.A(n_757),
.Y(n_2602)
);

CKINVDCx5p33_ASAP7_75t_R g2603 ( 
.A(n_230),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_849),
.Y(n_2604)
);

INVxp67_ASAP7_75t_L g2605 ( 
.A(n_926),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_1642),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_560),
.Y(n_2607)
);

BUFx6f_ASAP7_75t_L g2608 ( 
.A(n_613),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_390),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_1706),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_1858),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_1603),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_468),
.Y(n_2613)
);

CKINVDCx5p33_ASAP7_75t_R g2614 ( 
.A(n_156),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_1760),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_1486),
.Y(n_2616)
);

BUFx10_ASAP7_75t_L g2617 ( 
.A(n_1788),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_1646),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_1400),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_1678),
.Y(n_2620)
);

BUFx5_ASAP7_75t_L g2621 ( 
.A(n_622),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_94),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_215),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_1267),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_786),
.Y(n_2625)
);

CKINVDCx5p33_ASAP7_75t_R g2626 ( 
.A(n_1665),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_1767),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_1617),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_1700),
.Y(n_2629)
);

CKINVDCx16_ASAP7_75t_R g2630 ( 
.A(n_566),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_565),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_1519),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_1752),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_1658),
.Y(n_2634)
);

BUFx6f_ASAP7_75t_L g2635 ( 
.A(n_193),
.Y(n_2635)
);

CKINVDCx5p33_ASAP7_75t_R g2636 ( 
.A(n_1586),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_804),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_1632),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_362),
.Y(n_2639)
);

CKINVDCx5p33_ASAP7_75t_R g2640 ( 
.A(n_1819),
.Y(n_2640)
);

BUFx6f_ASAP7_75t_L g2641 ( 
.A(n_1724),
.Y(n_2641)
);

CKINVDCx5p33_ASAP7_75t_R g2642 ( 
.A(n_1119),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_931),
.Y(n_2643)
);

CKINVDCx20_ASAP7_75t_R g2644 ( 
.A(n_392),
.Y(n_2644)
);

CKINVDCx5p33_ASAP7_75t_R g2645 ( 
.A(n_375),
.Y(n_2645)
);

INVxp67_ASAP7_75t_L g2646 ( 
.A(n_1688),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_1028),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_1629),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_441),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_1686),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_915),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_808),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_898),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_845),
.Y(n_2654)
);

INVxp67_ASAP7_75t_SL g2655 ( 
.A(n_1246),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_309),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_1782),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_183),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_1847),
.Y(n_2659)
);

CKINVDCx5p33_ASAP7_75t_R g2660 ( 
.A(n_1164),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_1487),
.Y(n_2661)
);

INVx1_ASAP7_75t_SL g2662 ( 
.A(n_1901),
.Y(n_2662)
);

BUFx2_ASAP7_75t_L g2663 ( 
.A(n_1622),
.Y(n_2663)
);

CKINVDCx5p33_ASAP7_75t_R g2664 ( 
.A(n_1912),
.Y(n_2664)
);

CKINVDCx5p33_ASAP7_75t_R g2665 ( 
.A(n_1225),
.Y(n_2665)
);

BUFx6f_ASAP7_75t_L g2666 ( 
.A(n_19),
.Y(n_2666)
);

CKINVDCx5p33_ASAP7_75t_R g2667 ( 
.A(n_1150),
.Y(n_2667)
);

CKINVDCx5p33_ASAP7_75t_R g2668 ( 
.A(n_1113),
.Y(n_2668)
);

CKINVDCx5p33_ASAP7_75t_R g2669 ( 
.A(n_442),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_608),
.Y(n_2670)
);

BUFx10_ASAP7_75t_L g2671 ( 
.A(n_1282),
.Y(n_2671)
);

HB1xp67_ASAP7_75t_L g2672 ( 
.A(n_384),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_907),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_440),
.Y(n_2674)
);

BUFx10_ASAP7_75t_L g2675 ( 
.A(n_374),
.Y(n_2675)
);

CKINVDCx5p33_ASAP7_75t_R g2676 ( 
.A(n_886),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_719),
.Y(n_2677)
);

CKINVDCx5p33_ASAP7_75t_R g2678 ( 
.A(n_554),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_1098),
.Y(n_2679)
);

BUFx8_ASAP7_75t_SL g2680 ( 
.A(n_321),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_417),
.Y(n_2681)
);

CKINVDCx5p33_ASAP7_75t_R g2682 ( 
.A(n_1888),
.Y(n_2682)
);

CKINVDCx5p33_ASAP7_75t_R g2683 ( 
.A(n_1567),
.Y(n_2683)
);

CKINVDCx5p33_ASAP7_75t_R g2684 ( 
.A(n_1621),
.Y(n_2684)
);

CKINVDCx5p33_ASAP7_75t_R g2685 ( 
.A(n_1112),
.Y(n_2685)
);

INVx2_ASAP7_75t_SL g2686 ( 
.A(n_1628),
.Y(n_2686)
);

CKINVDCx5p33_ASAP7_75t_R g2687 ( 
.A(n_778),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_1716),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_1796),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_698),
.Y(n_2690)
);

CKINVDCx5p33_ASAP7_75t_R g2691 ( 
.A(n_179),
.Y(n_2691)
);

CKINVDCx5p33_ASAP7_75t_R g2692 ( 
.A(n_65),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_917),
.Y(n_2693)
);

CKINVDCx5p33_ASAP7_75t_R g2694 ( 
.A(n_1370),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_1761),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_1905),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_1625),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_1132),
.Y(n_2698)
);

CKINVDCx5p33_ASAP7_75t_R g2699 ( 
.A(n_560),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_1029),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_663),
.Y(n_2701)
);

CKINVDCx20_ASAP7_75t_R g2702 ( 
.A(n_663),
.Y(n_2702)
);

BUFx5_ASAP7_75t_L g2703 ( 
.A(n_1159),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_933),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_152),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_1649),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_222),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_98),
.Y(n_2708)
);

CKINVDCx16_ASAP7_75t_R g2709 ( 
.A(n_627),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_1727),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_610),
.Y(n_2711)
);

CKINVDCx5p33_ASAP7_75t_R g2712 ( 
.A(n_807),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_703),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_1200),
.Y(n_2714)
);

CKINVDCx5p33_ASAP7_75t_R g2715 ( 
.A(n_790),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_169),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_166),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_1715),
.Y(n_2718)
);

INVx1_ASAP7_75t_SL g2719 ( 
.A(n_473),
.Y(n_2719)
);

CKINVDCx5p33_ASAP7_75t_R g2720 ( 
.A(n_1028),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_682),
.Y(n_2721)
);

BUFx5_ASAP7_75t_L g2722 ( 
.A(n_1063),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_107),
.Y(n_2723)
);

CKINVDCx20_ASAP7_75t_R g2724 ( 
.A(n_1853),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_1720),
.Y(n_2725)
);

BUFx5_ASAP7_75t_L g2726 ( 
.A(n_163),
.Y(n_2726)
);

CKINVDCx20_ASAP7_75t_R g2727 ( 
.A(n_774),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_896),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_1636),
.Y(n_2729)
);

CKINVDCx5p33_ASAP7_75t_R g2730 ( 
.A(n_765),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_809),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_273),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_539),
.Y(n_2733)
);

CKINVDCx20_ASAP7_75t_R g2734 ( 
.A(n_1635),
.Y(n_2734)
);

CKINVDCx5p33_ASAP7_75t_R g2735 ( 
.A(n_94),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_1424),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_797),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_66),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_1749),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_236),
.Y(n_2740)
);

CKINVDCx5p33_ASAP7_75t_R g2741 ( 
.A(n_1743),
.Y(n_2741)
);

BUFx3_ASAP7_75t_L g2742 ( 
.A(n_1076),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_1261),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_1448),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_403),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_152),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_1063),
.Y(n_2747)
);

INVx1_ASAP7_75t_SL g2748 ( 
.A(n_622),
.Y(n_2748)
);

CKINVDCx14_ASAP7_75t_R g2749 ( 
.A(n_120),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_1059),
.Y(n_2750)
);

CKINVDCx5p33_ASAP7_75t_R g2751 ( 
.A(n_1616),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_1645),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_1155),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_883),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_1793),
.Y(n_2755)
);

CKINVDCx5p33_ASAP7_75t_R g2756 ( 
.A(n_1036),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_1633),
.Y(n_2757)
);

CKINVDCx5p33_ASAP7_75t_R g2758 ( 
.A(n_777),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_1067),
.Y(n_2759)
);

BUFx10_ASAP7_75t_L g2760 ( 
.A(n_1030),
.Y(n_2760)
);

BUFx3_ASAP7_75t_L g2761 ( 
.A(n_1570),
.Y(n_2761)
);

CKINVDCx5p33_ASAP7_75t_R g2762 ( 
.A(n_1154),
.Y(n_2762)
);

CKINVDCx5p33_ASAP7_75t_R g2763 ( 
.A(n_1801),
.Y(n_2763)
);

INVxp67_ASAP7_75t_L g2764 ( 
.A(n_1744),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_336),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_985),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_1233),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_1445),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_117),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_1647),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_1734),
.Y(n_2771)
);

CKINVDCx5p33_ASAP7_75t_R g2772 ( 
.A(n_1791),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_1289),
.Y(n_2773)
);

CKINVDCx14_ASAP7_75t_R g2774 ( 
.A(n_1320),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_1346),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_455),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_1492),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_187),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_1674),
.Y(n_2779)
);

INVx1_ASAP7_75t_SL g2780 ( 
.A(n_489),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_1775),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_1419),
.Y(n_2782)
);

CKINVDCx20_ASAP7_75t_R g2783 ( 
.A(n_1726),
.Y(n_2783)
);

CKINVDCx5p33_ASAP7_75t_R g2784 ( 
.A(n_1052),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_1828),
.Y(n_2785)
);

CKINVDCx5p33_ASAP7_75t_R g2786 ( 
.A(n_1016),
.Y(n_2786)
);

CKINVDCx5p33_ASAP7_75t_R g2787 ( 
.A(n_853),
.Y(n_2787)
);

CKINVDCx5p33_ASAP7_75t_R g2788 ( 
.A(n_1762),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_688),
.Y(n_2789)
);

CKINVDCx5p33_ASAP7_75t_R g2790 ( 
.A(n_1781),
.Y(n_2790)
);

CKINVDCx5p33_ASAP7_75t_R g2791 ( 
.A(n_45),
.Y(n_2791)
);

BUFx2_ASAP7_75t_L g2792 ( 
.A(n_1770),
.Y(n_2792)
);

CKINVDCx5p33_ASAP7_75t_R g2793 ( 
.A(n_558),
.Y(n_2793)
);

CKINVDCx20_ASAP7_75t_R g2794 ( 
.A(n_1409),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_598),
.Y(n_2795)
);

CKINVDCx20_ASAP7_75t_R g2796 ( 
.A(n_1899),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_944),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_1671),
.Y(n_2798)
);

CKINVDCx5p33_ASAP7_75t_R g2799 ( 
.A(n_637),
.Y(n_2799)
);

CKINVDCx5p33_ASAP7_75t_R g2800 ( 
.A(n_1786),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_1747),
.Y(n_2801)
);

BUFx6f_ASAP7_75t_L g2802 ( 
.A(n_438),
.Y(n_2802)
);

CKINVDCx5p33_ASAP7_75t_R g2803 ( 
.A(n_1129),
.Y(n_2803)
);

CKINVDCx5p33_ASAP7_75t_R g2804 ( 
.A(n_685),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_1347),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_414),
.Y(n_2806)
);

INVxp67_ASAP7_75t_L g2807 ( 
.A(n_1799),
.Y(n_2807)
);

CKINVDCx5p33_ASAP7_75t_R g2808 ( 
.A(n_108),
.Y(n_2808)
);

CKINVDCx5p33_ASAP7_75t_R g2809 ( 
.A(n_379),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_1699),
.Y(n_2810)
);

INVx2_ASAP7_75t_SL g2811 ( 
.A(n_906),
.Y(n_2811)
);

CKINVDCx20_ASAP7_75t_R g2812 ( 
.A(n_279),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_748),
.Y(n_2813)
);

CKINVDCx5p33_ASAP7_75t_R g2814 ( 
.A(n_981),
.Y(n_2814)
);

CKINVDCx5p33_ASAP7_75t_R g2815 ( 
.A(n_396),
.Y(n_2815)
);

CKINVDCx5p33_ASAP7_75t_R g2816 ( 
.A(n_769),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_143),
.Y(n_2817)
);

CKINVDCx14_ASAP7_75t_R g2818 ( 
.A(n_454),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_1903),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_1813),
.Y(n_2820)
);

INVx1_ASAP7_75t_SL g2821 ( 
.A(n_548),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_1610),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_1042),
.Y(n_2823)
);

BUFx10_ASAP7_75t_L g2824 ( 
.A(n_1748),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_118),
.Y(n_2825)
);

CKINVDCx5p33_ASAP7_75t_R g2826 ( 
.A(n_510),
.Y(n_2826)
);

CKINVDCx5p33_ASAP7_75t_R g2827 ( 
.A(n_166),
.Y(n_2827)
);

CKINVDCx5p33_ASAP7_75t_R g2828 ( 
.A(n_1251),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_1753),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_799),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_1607),
.Y(n_2831)
);

CKINVDCx5p33_ASAP7_75t_R g2832 ( 
.A(n_608),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_1702),
.Y(n_2833)
);

CKINVDCx5p33_ASAP7_75t_R g2834 ( 
.A(n_610),
.Y(n_2834)
);

CKINVDCx5p33_ASAP7_75t_R g2835 ( 
.A(n_1170),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_418),
.Y(n_2836)
);

CKINVDCx5p33_ASAP7_75t_R g2837 ( 
.A(n_505),
.Y(n_2837)
);

CKINVDCx5p33_ASAP7_75t_R g2838 ( 
.A(n_1453),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_913),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_1754),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_1910),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_464),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_56),
.Y(n_2843)
);

CKINVDCx5p33_ASAP7_75t_R g2844 ( 
.A(n_1634),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_1771),
.Y(n_2845)
);

CKINVDCx5p33_ASAP7_75t_R g2846 ( 
.A(n_1349),
.Y(n_2846)
);

CKINVDCx5p33_ASAP7_75t_R g2847 ( 
.A(n_1215),
.Y(n_2847)
);

CKINVDCx5p33_ASAP7_75t_R g2848 ( 
.A(n_922),
.Y(n_2848)
);

INVx1_ASAP7_75t_SL g2849 ( 
.A(n_450),
.Y(n_2849)
);

CKINVDCx5p33_ASAP7_75t_R g2850 ( 
.A(n_1234),
.Y(n_2850)
);

CKINVDCx5p33_ASAP7_75t_R g2851 ( 
.A(n_32),
.Y(n_2851)
);

CKINVDCx20_ASAP7_75t_R g2852 ( 
.A(n_1776),
.Y(n_2852)
);

CKINVDCx5p33_ASAP7_75t_R g2853 ( 
.A(n_908),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_1758),
.Y(n_2854)
);

BUFx6f_ASAP7_75t_L g2855 ( 
.A(n_618),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_505),
.Y(n_2856)
);

CKINVDCx5p33_ASAP7_75t_R g2857 ( 
.A(n_1172),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_615),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_1576),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_1534),
.Y(n_2860)
);

CKINVDCx5p33_ASAP7_75t_R g2861 ( 
.A(n_1234),
.Y(n_2861)
);

CKINVDCx20_ASAP7_75t_R g2862 ( 
.A(n_1751),
.Y(n_2862)
);

CKINVDCx5p33_ASAP7_75t_R g2863 ( 
.A(n_1041),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_825),
.Y(n_2864)
);

CKINVDCx5p33_ASAP7_75t_R g2865 ( 
.A(n_1692),
.Y(n_2865)
);

CKINVDCx5p33_ASAP7_75t_R g2866 ( 
.A(n_1160),
.Y(n_2866)
);

CKINVDCx5p33_ASAP7_75t_R g2867 ( 
.A(n_1157),
.Y(n_2867)
);

CKINVDCx5p33_ASAP7_75t_R g2868 ( 
.A(n_50),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_361),
.Y(n_2869)
);

BUFx3_ASAP7_75t_L g2870 ( 
.A(n_201),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_1519),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_755),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_969),
.Y(n_2873)
);

BUFx2_ASAP7_75t_L g2874 ( 
.A(n_356),
.Y(n_2874)
);

CKINVDCx5p33_ASAP7_75t_R g2875 ( 
.A(n_1669),
.Y(n_2875)
);

INVx1_ASAP7_75t_SL g2876 ( 
.A(n_893),
.Y(n_2876)
);

CKINVDCx5p33_ASAP7_75t_R g2877 ( 
.A(n_1630),
.Y(n_2877)
);

CKINVDCx20_ASAP7_75t_R g2878 ( 
.A(n_1579),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_1388),
.Y(n_2879)
);

INVx1_ASAP7_75t_SL g2880 ( 
.A(n_1793),
.Y(n_2880)
);

CKINVDCx5p33_ASAP7_75t_R g2881 ( 
.A(n_1909),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_423),
.Y(n_2882)
);

CKINVDCx5p33_ASAP7_75t_R g2883 ( 
.A(n_1575),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_1688),
.Y(n_2884)
);

CKINVDCx5p33_ASAP7_75t_R g2885 ( 
.A(n_1403),
.Y(n_2885)
);

CKINVDCx20_ASAP7_75t_R g2886 ( 
.A(n_1246),
.Y(n_2886)
);

CKINVDCx20_ASAP7_75t_R g2887 ( 
.A(n_1644),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_1467),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_786),
.Y(n_2889)
);

CKINVDCx5p33_ASAP7_75t_R g2890 ( 
.A(n_1059),
.Y(n_2890)
);

BUFx2_ASAP7_75t_SL g2891 ( 
.A(n_919),
.Y(n_2891)
);

CKINVDCx5p33_ASAP7_75t_R g2892 ( 
.A(n_1826),
.Y(n_2892)
);

CKINVDCx5p33_ASAP7_75t_R g2893 ( 
.A(n_418),
.Y(n_2893)
);

CKINVDCx5p33_ASAP7_75t_R g2894 ( 
.A(n_1504),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_1890),
.Y(n_2895)
);

CKINVDCx5p33_ASAP7_75t_R g2896 ( 
.A(n_466),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_1281),
.Y(n_2897)
);

CKINVDCx5p33_ASAP7_75t_R g2898 ( 
.A(n_1664),
.Y(n_2898)
);

CKINVDCx5p33_ASAP7_75t_R g2899 ( 
.A(n_1300),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_1598),
.Y(n_2900)
);

CKINVDCx5p33_ASAP7_75t_R g2901 ( 
.A(n_1379),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_676),
.Y(n_2902)
);

CKINVDCx5p33_ASAP7_75t_R g2903 ( 
.A(n_1047),
.Y(n_2903)
);

CKINVDCx20_ASAP7_75t_R g2904 ( 
.A(n_1560),
.Y(n_2904)
);

BUFx2_ASAP7_75t_L g2905 ( 
.A(n_1209),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_415),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_1320),
.Y(n_2907)
);

CKINVDCx5p33_ASAP7_75t_R g2908 ( 
.A(n_1735),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_1483),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_1066),
.Y(n_2910)
);

CKINVDCx5p33_ASAP7_75t_R g2911 ( 
.A(n_835),
.Y(n_2911)
);

CKINVDCx5p33_ASAP7_75t_R g2912 ( 
.A(n_1560),
.Y(n_2912)
);

CKINVDCx5p33_ASAP7_75t_R g2913 ( 
.A(n_743),
.Y(n_2913)
);

CKINVDCx5p33_ASAP7_75t_R g2914 ( 
.A(n_272),
.Y(n_2914)
);

CKINVDCx5p33_ASAP7_75t_R g2915 ( 
.A(n_371),
.Y(n_2915)
);

INVx2_ASAP7_75t_SL g2916 ( 
.A(n_885),
.Y(n_2916)
);

BUFx3_ASAP7_75t_L g2917 ( 
.A(n_1693),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_330),
.Y(n_2918)
);

CKINVDCx20_ASAP7_75t_R g2919 ( 
.A(n_1346),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_662),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_1787),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_1667),
.Y(n_2922)
);

CKINVDCx20_ASAP7_75t_R g2923 ( 
.A(n_1634),
.Y(n_2923)
);

CKINVDCx5p33_ASAP7_75t_R g2924 ( 
.A(n_496),
.Y(n_2924)
);

CKINVDCx5p33_ASAP7_75t_R g2925 ( 
.A(n_997),
.Y(n_2925)
);

CKINVDCx5p33_ASAP7_75t_R g2926 ( 
.A(n_281),
.Y(n_2926)
);

CKINVDCx5p33_ASAP7_75t_R g2927 ( 
.A(n_1487),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_344),
.Y(n_2928)
);

BUFx2_ASAP7_75t_L g2929 ( 
.A(n_1145),
.Y(n_2929)
);

CKINVDCx5p33_ASAP7_75t_R g2930 ( 
.A(n_1740),
.Y(n_2930)
);

CKINVDCx5p33_ASAP7_75t_R g2931 ( 
.A(n_1125),
.Y(n_2931)
);

CKINVDCx20_ASAP7_75t_R g2932 ( 
.A(n_1779),
.Y(n_2932)
);

CKINVDCx5p33_ASAP7_75t_R g2933 ( 
.A(n_569),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_1606),
.Y(n_2934)
);

CKINVDCx5p33_ASAP7_75t_R g2935 ( 
.A(n_252),
.Y(n_2935)
);

BUFx6f_ASAP7_75t_L g2936 ( 
.A(n_1195),
.Y(n_2936)
);

BUFx6f_ASAP7_75t_L g2937 ( 
.A(n_1651),
.Y(n_2937)
);

CKINVDCx5p33_ASAP7_75t_R g2938 ( 
.A(n_468),
.Y(n_2938)
);

CKINVDCx5p33_ASAP7_75t_R g2939 ( 
.A(n_1033),
.Y(n_2939)
);

CKINVDCx20_ASAP7_75t_R g2940 ( 
.A(n_1580),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_1698),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_1707),
.Y(n_2942)
);

CKINVDCx5p33_ASAP7_75t_R g2943 ( 
.A(n_186),
.Y(n_2943)
);

CKINVDCx5p33_ASAP7_75t_R g2944 ( 
.A(n_171),
.Y(n_2944)
);

CKINVDCx20_ASAP7_75t_R g2945 ( 
.A(n_1750),
.Y(n_2945)
);

INVx2_ASAP7_75t_SL g2946 ( 
.A(n_1335),
.Y(n_2946)
);

CKINVDCx5p33_ASAP7_75t_R g2947 ( 
.A(n_1705),
.Y(n_2947)
);

CKINVDCx5p33_ASAP7_75t_R g2948 ( 
.A(n_1640),
.Y(n_2948)
);

CKINVDCx5p33_ASAP7_75t_R g2949 ( 
.A(n_1742),
.Y(n_2949)
);

CKINVDCx5p33_ASAP7_75t_R g2950 ( 
.A(n_694),
.Y(n_2950)
);

CKINVDCx5p33_ASAP7_75t_R g2951 ( 
.A(n_1455),
.Y(n_2951)
);

CKINVDCx5p33_ASAP7_75t_R g2952 ( 
.A(n_246),
.Y(n_2952)
);

BUFx3_ASAP7_75t_L g2953 ( 
.A(n_492),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_487),
.Y(n_2954)
);

CKINVDCx5p33_ASAP7_75t_R g2955 ( 
.A(n_1099),
.Y(n_2955)
);

CKINVDCx5p33_ASAP7_75t_R g2956 ( 
.A(n_1184),
.Y(n_2956)
);

CKINVDCx5p33_ASAP7_75t_R g2957 ( 
.A(n_1443),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_743),
.Y(n_2958)
);

CKINVDCx5p33_ASAP7_75t_R g2959 ( 
.A(n_1725),
.Y(n_2959)
);

CKINVDCx5p33_ASAP7_75t_R g2960 ( 
.A(n_1555),
.Y(n_2960)
);

CKINVDCx5p33_ASAP7_75t_R g2961 ( 
.A(n_1367),
.Y(n_2961)
);

CKINVDCx5p33_ASAP7_75t_R g2962 ( 
.A(n_440),
.Y(n_2962)
);

BUFx3_ASAP7_75t_L g2963 ( 
.A(n_470),
.Y(n_2963)
);

CKINVDCx5p33_ASAP7_75t_R g2964 ( 
.A(n_1767),
.Y(n_2964)
);

CKINVDCx5p33_ASAP7_75t_R g2965 ( 
.A(n_249),
.Y(n_2965)
);

CKINVDCx5p33_ASAP7_75t_R g2966 ( 
.A(n_1673),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_465),
.Y(n_2967)
);

CKINVDCx5p33_ASAP7_75t_R g2968 ( 
.A(n_815),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_937),
.Y(n_2969)
);

CKINVDCx5p33_ASAP7_75t_R g2970 ( 
.A(n_1704),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_1021),
.Y(n_2971)
);

CKINVDCx20_ASAP7_75t_R g2972 ( 
.A(n_1737),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_1689),
.Y(n_2973)
);

BUFx2_ASAP7_75t_L g2974 ( 
.A(n_1264),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_272),
.Y(n_2975)
);

CKINVDCx5p33_ASAP7_75t_R g2976 ( 
.A(n_1679),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_473),
.Y(n_2977)
);

CKINVDCx5p33_ASAP7_75t_R g2978 ( 
.A(n_1783),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_87),
.Y(n_2979)
);

CKINVDCx5p33_ASAP7_75t_R g2980 ( 
.A(n_4),
.Y(n_2980)
);

CKINVDCx5p33_ASAP7_75t_R g2981 ( 
.A(n_727),
.Y(n_2981)
);

CKINVDCx5p33_ASAP7_75t_R g2982 ( 
.A(n_62),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_291),
.Y(n_2983)
);

CKINVDCx5p33_ASAP7_75t_R g2984 ( 
.A(n_405),
.Y(n_2984)
);

CKINVDCx5p33_ASAP7_75t_R g2985 ( 
.A(n_394),
.Y(n_2985)
);

CKINVDCx5p33_ASAP7_75t_R g2986 ( 
.A(n_1833),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_1153),
.Y(n_2987)
);

CKINVDCx5p33_ASAP7_75t_R g2988 ( 
.A(n_475),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_799),
.Y(n_2989)
);

CKINVDCx5p33_ASAP7_75t_R g2990 ( 
.A(n_1708),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_1),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_1638),
.Y(n_2992)
);

CKINVDCx5p33_ASAP7_75t_R g2993 ( 
.A(n_1610),
.Y(n_2993)
);

CKINVDCx5p33_ASAP7_75t_R g2994 ( 
.A(n_1769),
.Y(n_2994)
);

CKINVDCx5p33_ASAP7_75t_R g2995 ( 
.A(n_993),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_239),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_256),
.Y(n_2997)
);

CKINVDCx5p33_ASAP7_75t_R g2998 ( 
.A(n_1714),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_265),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_1631),
.Y(n_3000)
);

CKINVDCx5p33_ASAP7_75t_R g3001 ( 
.A(n_1818),
.Y(n_3001)
);

CKINVDCx16_ASAP7_75t_R g3002 ( 
.A(n_949),
.Y(n_3002)
);

CKINVDCx20_ASAP7_75t_R g3003 ( 
.A(n_402),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_1938),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_1931),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_1938),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_1938),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_1938),
.Y(n_3008)
);

BUFx2_ASAP7_75t_SL g3009 ( 
.A(n_2006),
.Y(n_3009)
);

CKINVDCx20_ASAP7_75t_R g3010 ( 
.A(n_2028),
.Y(n_3010)
);

INVxp33_ASAP7_75t_SL g3011 ( 
.A(n_2245),
.Y(n_3011)
);

BUFx6f_ASAP7_75t_L g3012 ( 
.A(n_1931),
.Y(n_3012)
);

CKINVDCx5p33_ASAP7_75t_R g3013 ( 
.A(n_2250),
.Y(n_3013)
);

BUFx3_ASAP7_75t_L g3014 ( 
.A(n_2427),
.Y(n_3014)
);

CKINVDCx5p33_ASAP7_75t_R g3015 ( 
.A(n_2680),
.Y(n_3015)
);

CKINVDCx20_ASAP7_75t_R g3016 ( 
.A(n_2293),
.Y(n_3016)
);

CKINVDCx14_ASAP7_75t_R g3017 ( 
.A(n_1943),
.Y(n_3017)
);

CKINVDCx5p33_ASAP7_75t_R g3018 ( 
.A(n_1930),
.Y(n_3018)
);

INVxp67_ASAP7_75t_SL g3019 ( 
.A(n_2516),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_1938),
.Y(n_3020)
);

CKINVDCx5p33_ASAP7_75t_R g3021 ( 
.A(n_1949),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2054),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2054),
.Y(n_3023)
);

HB1xp67_ASAP7_75t_L g3024 ( 
.A(n_3002),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2054),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2054),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2054),
.Y(n_3027)
);

CKINVDCx5p33_ASAP7_75t_R g3028 ( 
.A(n_1954),
.Y(n_3028)
);

INVxp67_ASAP7_75t_SL g3029 ( 
.A(n_2082),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2489),
.Y(n_3030)
);

INVxp67_ASAP7_75t_SL g3031 ( 
.A(n_2394),
.Y(n_3031)
);

INVxp67_ASAP7_75t_L g3032 ( 
.A(n_2058),
.Y(n_3032)
);

INVxp67_ASAP7_75t_SL g3033 ( 
.A(n_1980),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2489),
.Y(n_3034)
);

BUFx6f_ASAP7_75t_L g3035 ( 
.A(n_1931),
.Y(n_3035)
);

CKINVDCx16_ASAP7_75t_R g3036 ( 
.A(n_1953),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2489),
.Y(n_3037)
);

CKINVDCx20_ASAP7_75t_R g3038 ( 
.A(n_2363),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2489),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2489),
.Y(n_3040)
);

CKINVDCx16_ASAP7_75t_R g3041 ( 
.A(n_2038),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2621),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2621),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2621),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2621),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2621),
.Y(n_3046)
);

INVxp33_ASAP7_75t_SL g3047 ( 
.A(n_2272),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2703),
.Y(n_3048)
);

BUFx3_ASAP7_75t_L g3049 ( 
.A(n_2427),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2703),
.Y(n_3050)
);

INVxp67_ASAP7_75t_L g3051 ( 
.A(n_2159),
.Y(n_3051)
);

INVxp67_ASAP7_75t_SL g3052 ( 
.A(n_2301),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2703),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2703),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2703),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2722),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2722),
.Y(n_3057)
);

HB1xp67_ASAP7_75t_L g3058 ( 
.A(n_2105),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2722),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2722),
.Y(n_3060)
);

BUFx3_ASAP7_75t_L g3061 ( 
.A(n_2013),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2722),
.Y(n_3062)
);

CKINVDCx20_ASAP7_75t_R g3063 ( 
.A(n_2724),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2726),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2726),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2726),
.Y(n_3066)
);

CKINVDCx16_ASAP7_75t_R g3067 ( 
.A(n_2120),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2726),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2726),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_1945),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_1945),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_1945),
.Y(n_3072)
);

BUFx2_ASAP7_75t_L g3073 ( 
.A(n_2417),
.Y(n_3073)
);

CKINVDCx16_ASAP7_75t_R g3074 ( 
.A(n_2121),
.Y(n_3074)
);

INVxp67_ASAP7_75t_L g3075 ( 
.A(n_2440),
.Y(n_3075)
);

HB1xp67_ASAP7_75t_L g3076 ( 
.A(n_2135),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_1975),
.Y(n_3077)
);

CKINVDCx20_ASAP7_75t_R g3078 ( 
.A(n_2796),
.Y(n_3078)
);

BUFx2_ASAP7_75t_SL g3079 ( 
.A(n_2445),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_1975),
.Y(n_3080)
);

CKINVDCx5p33_ASAP7_75t_R g3081 ( 
.A(n_1957),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_1975),
.Y(n_3082)
);

INVxp67_ASAP7_75t_SL g3083 ( 
.A(n_2425),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_1985),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_1985),
.Y(n_3085)
);

BUFx3_ASAP7_75t_L g3086 ( 
.A(n_2039),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_1985),
.Y(n_3087)
);

HB1xp67_ASAP7_75t_L g3088 ( 
.A(n_2175),
.Y(n_3088)
);

CKINVDCx5p33_ASAP7_75t_R g3089 ( 
.A(n_1964),
.Y(n_3089)
);

CKINVDCx14_ASAP7_75t_R g3090 ( 
.A(n_2226),
.Y(n_3090)
);

INVxp67_ASAP7_75t_L g3091 ( 
.A(n_2567),
.Y(n_3091)
);

CKINVDCx5p33_ASAP7_75t_R g3092 ( 
.A(n_1978),
.Y(n_3092)
);

CKINVDCx20_ASAP7_75t_R g3093 ( 
.A(n_2409),
.Y(n_3093)
);

CKINVDCx5p33_ASAP7_75t_R g3094 ( 
.A(n_2052),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2019),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2019),
.Y(n_3096)
);

INVxp67_ASAP7_75t_SL g3097 ( 
.A(n_2455),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2019),
.Y(n_3098)
);

BUFx3_ASAP7_75t_L g3099 ( 
.A(n_2096),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2024),
.Y(n_3100)
);

CKINVDCx16_ASAP7_75t_R g3101 ( 
.A(n_2185),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2024),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2024),
.Y(n_3103)
);

BUFx10_ASAP7_75t_L g3104 ( 
.A(n_2610),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2076),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2076),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2076),
.Y(n_3107)
);

INVxp33_ASAP7_75t_SL g3108 ( 
.A(n_2672),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2145),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2145),
.Y(n_3110)
);

CKINVDCx5p33_ASAP7_75t_R g3111 ( 
.A(n_2066),
.Y(n_3111)
);

INVxp67_ASAP7_75t_SL g3112 ( 
.A(n_2145),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2152),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2152),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2152),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2188),
.Y(n_3116)
);

CKINVDCx20_ASAP7_75t_R g3117 ( 
.A(n_2235),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2188),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2188),
.Y(n_3119)
);

CKINVDCx5p33_ASAP7_75t_R g3120 ( 
.A(n_2072),
.Y(n_3120)
);

INVxp33_ASAP7_75t_SL g3121 ( 
.A(n_2663),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2240),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2240),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2240),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2275),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2275),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2275),
.Y(n_3127)
);

CKINVDCx5p33_ASAP7_75t_R g3128 ( 
.A(n_2093),
.Y(n_3128)
);

INVxp67_ASAP7_75t_SL g3129 ( 
.A(n_2399),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_2399),
.Y(n_3130)
);

NOR2xp33_ASAP7_75t_L g3131 ( 
.A(n_2333),
.B(n_0),
.Y(n_3131)
);

INVxp67_ASAP7_75t_L g3132 ( 
.A(n_2792),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2399),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2414),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2414),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2414),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2437),
.Y(n_3137)
);

BUFx6f_ASAP7_75t_L g3138 ( 
.A(n_2437),
.Y(n_3138)
);

CKINVDCx14_ASAP7_75t_R g3139 ( 
.A(n_2336),
.Y(n_3139)
);

BUFx6f_ASAP7_75t_L g3140 ( 
.A(n_2437),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2446),
.Y(n_3141)
);

INVx1_ASAP7_75t_SL g3142 ( 
.A(n_2874),
.Y(n_3142)
);

CKINVDCx20_ASAP7_75t_R g3143 ( 
.A(n_2749),
.Y(n_3143)
);

CKINVDCx16_ASAP7_75t_R g3144 ( 
.A(n_2236),
.Y(n_3144)
);

CKINVDCx5p33_ASAP7_75t_R g3145 ( 
.A(n_2097),
.Y(n_3145)
);

HB1xp67_ASAP7_75t_L g3146 ( 
.A(n_2350),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2446),
.Y(n_3147)
);

INVxp33_ASAP7_75t_SL g3148 ( 
.A(n_2905),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2446),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2452),
.Y(n_3150)
);

CKINVDCx5p33_ASAP7_75t_R g3151 ( 
.A(n_2101),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2452),
.Y(n_3152)
);

CKINVDCx16_ASAP7_75t_R g3153 ( 
.A(n_2435),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2452),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_2537),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2537),
.Y(n_3156)
);

CKINVDCx5p33_ASAP7_75t_R g3157 ( 
.A(n_2331),
.Y(n_3157)
);

BUFx2_ASAP7_75t_SL g3158 ( 
.A(n_2349),
.Y(n_3158)
);

INVxp33_ASAP7_75t_SL g3159 ( 
.A(n_2929),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2537),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2557),
.Y(n_3161)
);

INVxp67_ASAP7_75t_L g3162 ( 
.A(n_2974),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2557),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2557),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2592),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2592),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2592),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2608),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2608),
.Y(n_3169)
);

CKINVDCx20_ASAP7_75t_R g3170 ( 
.A(n_2774),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2608),
.Y(n_3171)
);

CKINVDCx5p33_ASAP7_75t_R g3172 ( 
.A(n_2415),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2635),
.Y(n_3173)
);

NOR2xp33_ASAP7_75t_L g3174 ( 
.A(n_2818),
.B(n_0),
.Y(n_3174)
);

INVxp67_ASAP7_75t_SL g3175 ( 
.A(n_2635),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2635),
.Y(n_3176)
);

CKINVDCx20_ASAP7_75t_R g3177 ( 
.A(n_3001),
.Y(n_3177)
);

CKINVDCx20_ASAP7_75t_R g3178 ( 
.A(n_2419),
.Y(n_3178)
);

CKINVDCx20_ASAP7_75t_R g3179 ( 
.A(n_2470),
.Y(n_3179)
);

INVx2_ASAP7_75t_SL g3180 ( 
.A(n_2109),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2641),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2641),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2641),
.Y(n_3183)
);

INVx2_ASAP7_75t_SL g3184 ( 
.A(n_2109),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2666),
.Y(n_3185)
);

INVxp67_ASAP7_75t_SL g3186 ( 
.A(n_2666),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2666),
.Y(n_3187)
);

INVxp67_ASAP7_75t_L g3188 ( 
.A(n_2030),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2802),
.Y(n_3189)
);

INVxp67_ASAP7_75t_SL g3190 ( 
.A(n_2802),
.Y(n_3190)
);

INVxp33_ASAP7_75t_SL g3191 ( 
.A(n_1926),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2802),
.Y(n_3192)
);

CKINVDCx16_ASAP7_75t_R g3193 ( 
.A(n_2496),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2855),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2855),
.Y(n_3195)
);

CKINVDCx5p33_ASAP7_75t_R g3196 ( 
.A(n_2553),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_2855),
.Y(n_3197)
);

BUFx3_ASAP7_75t_L g3198 ( 
.A(n_2176),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2936),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2936),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2936),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2937),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2937),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2937),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2979),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2979),
.Y(n_3206)
);

CKINVDCx5p33_ASAP7_75t_R g3207 ( 
.A(n_2611),
.Y(n_3207)
);

INVxp67_ASAP7_75t_SL g3208 ( 
.A(n_2979),
.Y(n_3208)
);

CKINVDCx5p33_ASAP7_75t_R g3209 ( 
.A(n_2640),
.Y(n_3209)
);

INVxp67_ASAP7_75t_L g3210 ( 
.A(n_2162),
.Y(n_3210)
);

INVxp67_ASAP7_75t_SL g3211 ( 
.A(n_2209),
.Y(n_3211)
);

CKINVDCx16_ASAP7_75t_R g3212 ( 
.A(n_2541),
.Y(n_3212)
);

INVxp33_ASAP7_75t_SL g3213 ( 
.A(n_1933),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2216),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2280),
.Y(n_3215)
);

INVx1_ASAP7_75t_SL g3216 ( 
.A(n_1947),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2295),
.Y(n_3217)
);

INVxp67_ASAP7_75t_L g3218 ( 
.A(n_2162),
.Y(n_3218)
);

BUFx2_ASAP7_75t_L g3219 ( 
.A(n_2392),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2491),
.Y(n_3220)
);

CKINVDCx5p33_ASAP7_75t_R g3221 ( 
.A(n_2664),
.Y(n_3221)
);

CKINVDCx5p33_ASAP7_75t_R g3222 ( 
.A(n_2682),
.Y(n_3222)
);

INVx4_ASAP7_75t_R g3223 ( 
.A(n_2091),
.Y(n_3223)
);

CKINVDCx16_ASAP7_75t_R g3224 ( 
.A(n_2630),
.Y(n_3224)
);

CKINVDCx5p33_ASAP7_75t_R g3225 ( 
.A(n_2696),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2572),
.Y(n_3226)
);

HB1xp67_ASAP7_75t_L g3227 ( 
.A(n_2709),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2742),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2761),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2870),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2917),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2953),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_2963),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_1925),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_1928),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_1929),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2996),
.Y(n_3237)
);

BUFx3_ASAP7_75t_L g3238 ( 
.A(n_2881),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2997),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3000),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_1934),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_1936),
.Y(n_3242)
);

BUFx3_ASAP7_75t_L g3243 ( 
.A(n_2892),
.Y(n_3243)
);

INVx2_ASAP7_75t_L g3244 ( 
.A(n_1941),
.Y(n_3244)
);

INVx4_ASAP7_75t_R g3245 ( 
.A(n_2662),
.Y(n_3245)
);

INVxp67_ASAP7_75t_SL g3246 ( 
.A(n_2010),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2989),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2991),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2992),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_1944),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_1955),
.Y(n_3251)
);

CKINVDCx5p33_ASAP7_75t_R g3252 ( 
.A(n_2986),
.Y(n_3252)
);

INVxp33_ASAP7_75t_SL g3253 ( 
.A(n_1937),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_1956),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_1961),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_1963),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_1965),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_1974),
.Y(n_3258)
);

CKINVDCx5p33_ASAP7_75t_R g3259 ( 
.A(n_2999),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_1981),
.Y(n_3260)
);

CKINVDCx20_ASAP7_75t_R g3261 ( 
.A(n_1939),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2983),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_1983),
.Y(n_3263)
);

BUFx3_ASAP7_75t_L g3264 ( 
.A(n_2177),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_3070),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_3084),
.Y(n_3266)
);

OA21x2_ASAP7_75t_L g3267 ( 
.A1(n_3004),
.A2(n_2074),
.B(n_2011),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_3109),
.Y(n_3268)
);

INVx3_ASAP7_75t_L g3269 ( 
.A(n_3005),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3112),
.Y(n_3270)
);

BUFx6f_ASAP7_75t_L g3271 ( 
.A(n_3005),
.Y(n_3271)
);

AND2x4_ASAP7_75t_L g3272 ( 
.A(n_3238),
.B(n_2127),
.Y(n_3272)
);

AOI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_3121),
.A2(n_2655),
.B1(n_1998),
.B2(n_1940),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3129),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3123),
.Y(n_3275)
);

INVx2_ASAP7_75t_SL g3276 ( 
.A(n_3104),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_3012),
.Y(n_3277)
);

OAI21x1_ASAP7_75t_L g3278 ( 
.A1(n_3023),
.A2(n_2505),
.B(n_2384),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3130),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3175),
.Y(n_3280)
);

BUFx6f_ASAP7_75t_L g3281 ( 
.A(n_3012),
.Y(n_3281)
);

BUFx6f_ASAP7_75t_L g3282 ( 
.A(n_3035),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_3018),
.B(n_2785),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_3135),
.Y(n_3284)
);

BUFx6f_ASAP7_75t_L g3285 ( 
.A(n_3035),
.Y(n_3285)
);

AND2x4_ASAP7_75t_L g3286 ( 
.A(n_3243),
.B(n_2229),
.Y(n_3286)
);

INVx5_ASAP7_75t_L g3287 ( 
.A(n_3180),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3186),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3190),
.Y(n_3289)
);

AOI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_3148),
.A2(n_1946),
.B1(n_1951),
.B2(n_1950),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3155),
.Y(n_3291)
);

OA21x2_ASAP7_75t_L g3292 ( 
.A1(n_3006),
.A2(n_2313),
.B(n_2247),
.Y(n_3292)
);

BUFx6f_ASAP7_75t_L g3293 ( 
.A(n_3138),
.Y(n_3293)
);

BUFx6f_ASAP7_75t_L g3294 ( 
.A(n_3138),
.Y(n_3294)
);

BUFx8_ASAP7_75t_L g3295 ( 
.A(n_3073),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_SL g3296 ( 
.A(n_3036),
.B(n_2177),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3021),
.B(n_2659),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3208),
.Y(n_3298)
);

INVx4_ASAP7_75t_L g3299 ( 
.A(n_3028),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_3017),
.B(n_1932),
.Y(n_3300)
);

BUFx6f_ASAP7_75t_L g3301 ( 
.A(n_3140),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3140),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_3164),
.Y(n_3303)
);

INVx5_ASAP7_75t_L g3304 ( 
.A(n_3184),
.Y(n_3304)
);

OAI22x1_ASAP7_75t_L g3305 ( 
.A1(n_3142),
.A2(n_1968),
.B1(n_1993),
.B2(n_1924),
.Y(n_3305)
);

AOI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_3159),
.A2(n_1952),
.B1(n_1959),
.B2(n_1958),
.Y(n_3306)
);

INVx3_ASAP7_75t_L g3307 ( 
.A(n_3061),
.Y(n_3307)
);

INVx3_ASAP7_75t_L g3308 ( 
.A(n_3086),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3081),
.B(n_2819),
.Y(n_3309)
);

BUFx8_ASAP7_75t_L g3310 ( 
.A(n_3219),
.Y(n_3310)
);

BUFx6f_ASAP7_75t_L g3311 ( 
.A(n_3166),
.Y(n_3311)
);

BUFx6f_ASAP7_75t_L g3312 ( 
.A(n_3168),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_3191),
.B(n_2820),
.Y(n_3313)
);

AND2x4_ASAP7_75t_L g3314 ( 
.A(n_3014),
.B(n_2841),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3089),
.B(n_2895),
.Y(n_3315)
);

BUFx12f_ASAP7_75t_L g3316 ( 
.A(n_3013),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_3183),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3195),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3092),
.B(n_2355),
.Y(n_3319)
);

BUFx6f_ASAP7_75t_L g3320 ( 
.A(n_3202),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_3071),
.Y(n_3321)
);

BUFx12f_ASAP7_75t_L g3322 ( 
.A(n_3015),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3072),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_3041),
.B(n_2212),
.Y(n_3324)
);

INVx3_ASAP7_75t_L g3325 ( 
.A(n_3099),
.Y(n_3325)
);

CKINVDCx5p33_ASAP7_75t_R g3326 ( 
.A(n_3094),
.Y(n_3326)
);

BUFx6f_ASAP7_75t_L g3327 ( 
.A(n_3198),
.Y(n_3327)
);

BUFx6f_ASAP7_75t_L g3328 ( 
.A(n_3077),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3080),
.Y(n_3329)
);

INVx3_ASAP7_75t_L g3330 ( 
.A(n_3233),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_3082),
.Y(n_3331)
);

BUFx6f_ASAP7_75t_L g3332 ( 
.A(n_3085),
.Y(n_3332)
);

INVx3_ASAP7_75t_L g3333 ( 
.A(n_3087),
.Y(n_3333)
);

AOI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_3011),
.A2(n_1960),
.B1(n_1967),
.B2(n_1962),
.Y(n_3334)
);

BUFx6f_ASAP7_75t_L g3335 ( 
.A(n_3095),
.Y(n_3335)
);

CKINVDCx6p67_ASAP7_75t_R g3336 ( 
.A(n_3117),
.Y(n_3336)
);

OA21x2_ASAP7_75t_L g3337 ( 
.A1(n_3007),
.A2(n_1935),
.B(n_1927),
.Y(n_3337)
);

CKINVDCx5p33_ASAP7_75t_R g3338 ( 
.A(n_3111),
.Y(n_3338)
);

HB1xp67_ASAP7_75t_L g3339 ( 
.A(n_3188),
.Y(n_3339)
);

AND2x4_ASAP7_75t_L g3340 ( 
.A(n_3049),
.B(n_2048),
.Y(n_3340)
);

BUFx6f_ASAP7_75t_L g3341 ( 
.A(n_3096),
.Y(n_3341)
);

BUFx6f_ASAP7_75t_L g3342 ( 
.A(n_3098),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_3100),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3102),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3103),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3105),
.Y(n_3346)
);

OAI21x1_ASAP7_75t_L g3347 ( 
.A1(n_3042),
.A2(n_1976),
.B(n_1942),
.Y(n_3347)
);

OAI21x1_ASAP7_75t_L g3348 ( 
.A1(n_3056),
.A2(n_2020),
.B(n_1986),
.Y(n_3348)
);

OR2x6_ASAP7_75t_L g3349 ( 
.A(n_3009),
.B(n_1995),
.Y(n_3349)
);

AOI22xp5_ASAP7_75t_L g3350 ( 
.A1(n_3047),
.A2(n_1970),
.B1(n_1973),
.B2(n_1969),
.Y(n_3350)
);

AND2x6_ASAP7_75t_L g3351 ( 
.A(n_3131),
.B(n_1999),
.Y(n_3351)
);

INVx3_ASAP7_75t_L g3352 ( 
.A(n_3106),
.Y(n_3352)
);

XNOR2x1_ASAP7_75t_L g3353 ( 
.A(n_3216),
.B(n_1977),
.Y(n_3353)
);

OAI21x1_ASAP7_75t_L g3354 ( 
.A1(n_3065),
.A2(n_2099),
.B(n_2080),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3107),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_3110),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3113),
.Y(n_3357)
);

BUFx6f_ASAP7_75t_L g3358 ( 
.A(n_3114),
.Y(n_3358)
);

CKINVDCx16_ASAP7_75t_R g3359 ( 
.A(n_3143),
.Y(n_3359)
);

INVx3_ASAP7_75t_L g3360 ( 
.A(n_3115),
.Y(n_3360)
);

CKINVDCx16_ASAP7_75t_R g3361 ( 
.A(n_3170),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_3067),
.B(n_2212),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3120),
.B(n_2355),
.Y(n_3363)
);

AND2x6_ASAP7_75t_L g3364 ( 
.A(n_3174),
.B(n_2134),
.Y(n_3364)
);

INVx5_ASAP7_75t_L g3365 ( 
.A(n_3264),
.Y(n_3365)
);

CKINVDCx16_ASAP7_75t_R g3366 ( 
.A(n_3074),
.Y(n_3366)
);

BUFx6f_ASAP7_75t_L g3367 ( 
.A(n_3116),
.Y(n_3367)
);

BUFx6f_ASAP7_75t_L g3368 ( 
.A(n_3118),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3119),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3122),
.Y(n_3370)
);

INVxp67_ASAP7_75t_L g3371 ( 
.A(n_3024),
.Y(n_3371)
);

AOI22xp5_ASAP7_75t_L g3372 ( 
.A1(n_3108),
.A2(n_3093),
.B1(n_3144),
.B2(n_3101),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3128),
.B(n_2355),
.Y(n_3373)
);

BUFx3_ASAP7_75t_L g3374 ( 
.A(n_3177),
.Y(n_3374)
);

OAI22x1_ASAP7_75t_SL g3375 ( 
.A1(n_3261),
.A2(n_1966),
.B1(n_1971),
.B2(n_1948),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3124),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3125),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_3126),
.Y(n_3378)
);

NOR2xp33_ASAP7_75t_L g3379 ( 
.A(n_3213),
.B(n_2138),
.Y(n_3379)
);

BUFx3_ASAP7_75t_L g3380 ( 
.A(n_3178),
.Y(n_3380)
);

BUFx6f_ASAP7_75t_L g3381 ( 
.A(n_3127),
.Y(n_3381)
);

BUFx6f_ASAP7_75t_L g3382 ( 
.A(n_3133),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3145),
.B(n_2179),
.Y(n_3383)
);

AND2x4_ASAP7_75t_L g3384 ( 
.A(n_3019),
.B(n_2248),
.Y(n_3384)
);

OAI22xp5_ASAP7_75t_L g3385 ( 
.A1(n_3032),
.A2(n_2391),
.B1(n_2467),
.B2(n_2358),
.Y(n_3385)
);

OAI22x1_ASAP7_75t_SL g3386 ( 
.A1(n_3010),
.A2(n_2001),
.B1(n_2018),
.B2(n_1972),
.Y(n_3386)
);

BUFx8_ASAP7_75t_L g3387 ( 
.A(n_3214),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_L g3388 ( 
.A(n_3253),
.B(n_2257),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3134),
.Y(n_3389)
);

OAI22x1_ASAP7_75t_L g3390 ( 
.A1(n_3210),
.A2(n_2199),
.B1(n_2215),
.B2(n_2158),
.Y(n_3390)
);

BUFx2_ASAP7_75t_L g3391 ( 
.A(n_3259),
.Y(n_3391)
);

BUFx12f_ASAP7_75t_L g3392 ( 
.A(n_3151),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3136),
.Y(n_3393)
);

AND2x6_ASAP7_75t_L g3394 ( 
.A(n_3215),
.B(n_2285),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3137),
.Y(n_3395)
);

BUFx3_ASAP7_75t_L g3396 ( 
.A(n_3179),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_3141),
.Y(n_3397)
);

BUFx3_ASAP7_75t_L g3398 ( 
.A(n_3217),
.Y(n_3398)
);

BUFx2_ASAP7_75t_L g3399 ( 
.A(n_3090),
.Y(n_3399)
);

OAI21x1_ASAP7_75t_L g3400 ( 
.A1(n_3008),
.A2(n_2125),
.B(n_2111),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3139),
.B(n_3029),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3147),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3157),
.B(n_2264),
.Y(n_3403)
);

BUFx2_ASAP7_75t_L g3404 ( 
.A(n_3058),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3149),
.Y(n_3405)
);

BUFx6f_ASAP7_75t_L g3406 ( 
.A(n_3150),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3172),
.B(n_2397),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3152),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3154),
.Y(n_3409)
);

INVx2_ASAP7_75t_L g3410 ( 
.A(n_3156),
.Y(n_3410)
);

BUFx6f_ASAP7_75t_L g3411 ( 
.A(n_3160),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3161),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3196),
.B(n_2464),
.Y(n_3413)
);

BUFx6f_ASAP7_75t_L g3414 ( 
.A(n_3163),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_3079),
.B(n_2490),
.Y(n_3415)
);

AOI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3153),
.A2(n_1982),
.B1(n_1988),
.B2(n_1979),
.Y(n_3416)
);

INVx5_ASAP7_75t_L g3417 ( 
.A(n_3193),
.Y(n_3417)
);

BUFx6f_ASAP7_75t_L g3418 ( 
.A(n_3165),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_3167),
.Y(n_3419)
);

INVx2_ASAP7_75t_SL g3420 ( 
.A(n_3220),
.Y(n_3420)
);

AND2x2_ASAP7_75t_SL g3421 ( 
.A(n_3212),
.B(n_2144),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3169),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_3171),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_3173),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3031),
.B(n_2525),
.Y(n_3425)
);

BUFx6f_ASAP7_75t_L g3426 ( 
.A(n_3176),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3181),
.Y(n_3427)
);

INVx5_ASAP7_75t_L g3428 ( 
.A(n_3224),
.Y(n_3428)
);

OA21x2_ASAP7_75t_L g3429 ( 
.A1(n_3020),
.A2(n_3025),
.B(n_3022),
.Y(n_3429)
);

INVx4_ASAP7_75t_L g3430 ( 
.A(n_3207),
.Y(n_3430)
);

INVx3_ASAP7_75t_L g3431 ( 
.A(n_3182),
.Y(n_3431)
);

BUFx6f_ASAP7_75t_L g3432 ( 
.A(n_3185),
.Y(n_3432)
);

OAI22x1_ASAP7_75t_R g3433 ( 
.A1(n_3016),
.A2(n_2036),
.B1(n_2049),
.B2(n_2029),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3187),
.Y(n_3434)
);

INVx3_ASAP7_75t_L g3435 ( 
.A(n_3189),
.Y(n_3435)
);

OAI22xp5_ASAP7_75t_SL g3436 ( 
.A1(n_3038),
.A2(n_2062),
.B1(n_2079),
.B2(n_2061),
.Y(n_3436)
);

AND2x4_ASAP7_75t_L g3437 ( 
.A(n_3033),
.B(n_2686),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_3192),
.Y(n_3438)
);

OA21x2_ASAP7_75t_L g3439 ( 
.A1(n_3026),
.A2(n_2224),
.B(n_2183),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3209),
.B(n_2689),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_3194),
.Y(n_3441)
);

BUFx2_ASAP7_75t_L g3442 ( 
.A(n_3076),
.Y(n_3442)
);

BUFx8_ASAP7_75t_L g3443 ( 
.A(n_3226),
.Y(n_3443)
);

INVx2_ASAP7_75t_L g3444 ( 
.A(n_3197),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3199),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3200),
.Y(n_3446)
);

OAI21x1_ASAP7_75t_L g3447 ( 
.A1(n_3027),
.A2(n_2254),
.B(n_2241),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3201),
.Y(n_3448)
);

INVx5_ASAP7_75t_L g3449 ( 
.A(n_3234),
.Y(n_3449)
);

BUFx8_ASAP7_75t_L g3450 ( 
.A(n_3228),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3203),
.Y(n_3451)
);

AND2x2_ASAP7_75t_L g3452 ( 
.A(n_3211),
.B(n_2811),
.Y(n_3452)
);

INVx3_ASAP7_75t_L g3453 ( 
.A(n_3204),
.Y(n_3453)
);

BUFx8_ASAP7_75t_L g3454 ( 
.A(n_3229),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3205),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3206),
.Y(n_3456)
);

BUFx6f_ASAP7_75t_L g3457 ( 
.A(n_3235),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3052),
.B(n_3083),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_L g3459 ( 
.A(n_3221),
.B(n_2916),
.Y(n_3459)
);

OAI21x1_ASAP7_75t_L g3460 ( 
.A1(n_3030),
.A2(n_2287),
.B(n_2281),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3222),
.B(n_2946),
.Y(n_3461)
);

AND2x2_ASAP7_75t_L g3462 ( 
.A(n_3097),
.B(n_2220),
.Y(n_3462)
);

INVx4_ASAP7_75t_L g3463 ( 
.A(n_3225),
.Y(n_3463)
);

AND2x2_ASAP7_75t_SL g3464 ( 
.A(n_3088),
.B(n_2290),
.Y(n_3464)
);

OAI21x1_ASAP7_75t_L g3465 ( 
.A1(n_3034),
.A2(n_2334),
.B(n_2329),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3037),
.Y(n_3466)
);

BUFx8_ASAP7_75t_L g3467 ( 
.A(n_3230),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_3039),
.Y(n_3468)
);

AND2x4_ASAP7_75t_L g3469 ( 
.A(n_3051),
.B(n_2353),
.Y(n_3469)
);

BUFx2_ASAP7_75t_L g3470 ( 
.A(n_3146),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3252),
.B(n_2220),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3040),
.Y(n_3472)
);

INVx3_ASAP7_75t_L g3473 ( 
.A(n_3236),
.Y(n_3473)
);

BUFx3_ASAP7_75t_L g3474 ( 
.A(n_3231),
.Y(n_3474)
);

OA21x2_ASAP7_75t_L g3475 ( 
.A1(n_3043),
.A2(n_2380),
.B(n_2359),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3044),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3045),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3466),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3476),
.Y(n_3479)
);

HB1xp67_ASAP7_75t_L g3480 ( 
.A(n_3307),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_SL g3481 ( 
.A(n_3366),
.B(n_3063),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3319),
.B(n_3246),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3477),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3311),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3468),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3472),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3398),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3474),
.Y(n_3488)
);

INVx3_ASAP7_75t_L g3489 ( 
.A(n_3327),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3312),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3457),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3363),
.B(n_3158),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3320),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3330),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3270),
.Y(n_3495)
);

AND2x6_ASAP7_75t_L g3496 ( 
.A(n_3300),
.B(n_3232),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3274),
.Y(n_3497)
);

BUFx8_ASAP7_75t_L g3498 ( 
.A(n_3404),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3265),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3280),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3288),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3289),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_3266),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3298),
.Y(n_3504)
);

NAND3xp33_ASAP7_75t_L g3505 ( 
.A(n_3379),
.B(n_3091),
.C(n_3075),
.Y(n_3505)
);

NAND2x1p5_ASAP7_75t_L g3506 ( 
.A(n_3308),
.B(n_3237),
.Y(n_3506)
);

AND2x4_ASAP7_75t_L g3507 ( 
.A(n_3272),
.B(n_3286),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3337),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3439),
.Y(n_3509)
);

BUFx8_ASAP7_75t_L g3510 ( 
.A(n_3442),
.Y(n_3510)
);

BUFx2_ASAP7_75t_L g3511 ( 
.A(n_3470),
.Y(n_3511)
);

NAND3xp33_ASAP7_75t_L g3512 ( 
.A(n_3388),
.B(n_3162),
.C(n_3132),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3373),
.B(n_3046),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_SL g3514 ( 
.A(n_3421),
.B(n_3227),
.Y(n_3514)
);

INVx3_ASAP7_75t_L g3515 ( 
.A(n_3271),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3475),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3268),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3400),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3447),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3460),
.Y(n_3520)
);

INVx3_ASAP7_75t_L g3521 ( 
.A(n_3281),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3465),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3323),
.Y(n_3523)
);

INVxp67_ASAP7_75t_L g3524 ( 
.A(n_3353),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3283),
.B(n_3048),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3329),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3344),
.Y(n_3527)
);

BUFx2_ASAP7_75t_L g3528 ( 
.A(n_3310),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3355),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3297),
.B(n_3050),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3357),
.Y(n_3531)
);

NAND2xp33_ASAP7_75t_SL g3532 ( 
.A(n_3305),
.B(n_2110),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3369),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3275),
.Y(n_3534)
);

OA21x2_ASAP7_75t_L g3535 ( 
.A1(n_3278),
.A2(n_3054),
.B(n_3053),
.Y(n_3535)
);

OA21x2_ASAP7_75t_L g3536 ( 
.A1(n_3347),
.A2(n_3057),
.B(n_3055),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3370),
.Y(n_3537)
);

BUFx6f_ASAP7_75t_L g3538 ( 
.A(n_3282),
.Y(n_3538)
);

AND2x2_ASAP7_75t_L g3539 ( 
.A(n_3339),
.B(n_3218),
.Y(n_3539)
);

HB1xp67_ASAP7_75t_L g3540 ( 
.A(n_3325),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3376),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3377),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3389),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3279),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3395),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3402),
.Y(n_3546)
);

INVx3_ASAP7_75t_L g3547 ( 
.A(n_3285),
.Y(n_3547)
);

BUFx6f_ASAP7_75t_L g3548 ( 
.A(n_3293),
.Y(n_3548)
);

BUFx6f_ASAP7_75t_L g3549 ( 
.A(n_3294),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3405),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3409),
.Y(n_3551)
);

BUFx6f_ASAP7_75t_L g3552 ( 
.A(n_3301),
.Y(n_3552)
);

BUFx6f_ASAP7_75t_L g3553 ( 
.A(n_3328),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3422),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3427),
.Y(n_3555)
);

OAI21x1_ASAP7_75t_L g3556 ( 
.A1(n_3348),
.A2(n_3060),
.B(n_3059),
.Y(n_3556)
);

OAI21x1_ASAP7_75t_L g3557 ( 
.A1(n_3354),
.A2(n_3064),
.B(n_3062),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3456),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3284),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3458),
.B(n_3244),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3291),
.Y(n_3561)
);

AOI22xp5_ASAP7_75t_L g3562 ( 
.A1(n_3351),
.A2(n_3078),
.B1(n_2341),
.B2(n_2351),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3401),
.B(n_3239),
.Y(n_3563)
);

AND2x2_ASAP7_75t_L g3564 ( 
.A(n_3425),
.B(n_3240),
.Y(n_3564)
);

INVxp67_ASAP7_75t_L g3565 ( 
.A(n_3415),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3303),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3317),
.Y(n_3567)
);

AND2x2_ASAP7_75t_L g3568 ( 
.A(n_3462),
.B(n_3241),
.Y(n_3568)
);

OA21x2_ASAP7_75t_L g3569 ( 
.A1(n_3309),
.A2(n_3068),
.B(n_3066),
.Y(n_3569)
);

BUFx6f_ASAP7_75t_L g3570 ( 
.A(n_3332),
.Y(n_3570)
);

NOR2xp33_ASAP7_75t_L g3571 ( 
.A(n_3315),
.B(n_3383),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3321),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3302),
.Y(n_3573)
);

AND2x6_ASAP7_75t_L g3574 ( 
.A(n_3471),
.B(n_3242),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3331),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3473),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3420),
.Y(n_3577)
);

BUFx6f_ASAP7_75t_L g3578 ( 
.A(n_3335),
.Y(n_3578)
);

INVx2_ASAP7_75t_L g3579 ( 
.A(n_3343),
.Y(n_3579)
);

AND2x4_ASAP7_75t_L g3580 ( 
.A(n_3314),
.B(n_3247),
.Y(n_3580)
);

BUFx6f_ASAP7_75t_L g3581 ( 
.A(n_3341),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3429),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3313),
.B(n_3459),
.Y(n_3583)
);

BUFx6f_ASAP7_75t_L g3584 ( 
.A(n_3342),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3333),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3352),
.Y(n_3586)
);

INVx4_ASAP7_75t_L g3587 ( 
.A(n_3392),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3452),
.B(n_3403),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3360),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3407),
.B(n_3069),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3345),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3431),
.Y(n_3592)
);

NAND2x1p5_ASAP7_75t_L g3593 ( 
.A(n_3417),
.B(n_3248),
.Y(n_3593)
);

AND2x4_ASAP7_75t_L g3594 ( 
.A(n_3349),
.B(n_3249),
.Y(n_3594)
);

BUFx8_ASAP7_75t_L g3595 ( 
.A(n_3316),
.Y(n_3595)
);

BUFx2_ASAP7_75t_L g3596 ( 
.A(n_3295),
.Y(n_3596)
);

CKINVDCx5p33_ASAP7_75t_R g3597 ( 
.A(n_3326),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3435),
.Y(n_3598)
);

NAND2xp33_ASAP7_75t_SL g3599 ( 
.A(n_3390),
.B(n_2116),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3453),
.Y(n_3600)
);

INVx3_ASAP7_75t_L g3601 ( 
.A(n_3269),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3346),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_3356),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3378),
.Y(n_3604)
);

OAI22xp5_ASAP7_75t_L g3605 ( 
.A1(n_3273),
.A2(n_2605),
.B1(n_2646),
.B2(n_2518),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3393),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_SL g3607 ( 
.A(n_3464),
.B(n_3223),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_3397),
.Y(n_3608)
);

AND3x1_ASAP7_75t_L g3609 ( 
.A(n_3334),
.B(n_1987),
.C(n_1984),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3408),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3410),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_3412),
.Y(n_3612)
);

INVx2_ASAP7_75t_L g3613 ( 
.A(n_3419),
.Y(n_3613)
);

OAI21x1_ASAP7_75t_L g3614 ( 
.A1(n_3267),
.A2(n_3251),
.B(n_3250),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_L g3615 ( 
.A(n_3413),
.B(n_3254),
.Y(n_3615)
);

HB1xp67_ASAP7_75t_L g3616 ( 
.A(n_3371),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_L g3617 ( 
.A(n_3440),
.B(n_3255),
.Y(n_3617)
);

BUFx6f_ASAP7_75t_L g3618 ( 
.A(n_3358),
.Y(n_3618)
);

OA21x2_ASAP7_75t_L g3619 ( 
.A1(n_3461),
.A2(n_3257),
.B(n_3256),
.Y(n_3619)
);

AND2x4_ASAP7_75t_L g3620 ( 
.A(n_3340),
.B(n_3258),
.Y(n_3620)
);

INVx2_ASAP7_75t_L g3621 ( 
.A(n_3423),
.Y(n_3621)
);

AND2x6_ASAP7_75t_L g3622 ( 
.A(n_3384),
.B(n_3260),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3424),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3434),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_3287),
.B(n_3245),
.Y(n_3625)
);

BUFx6f_ASAP7_75t_L g3626 ( 
.A(n_3367),
.Y(n_3626)
);

BUFx6f_ASAP7_75t_L g3627 ( 
.A(n_3368),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3438),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3441),
.Y(n_3629)
);

BUFx6f_ASAP7_75t_L g3630 ( 
.A(n_3381),
.Y(n_3630)
);

NAND2x1_ASAP7_75t_L g3631 ( 
.A(n_3292),
.B(n_2034),
.Y(n_3631)
);

BUFx6f_ASAP7_75t_L g3632 ( 
.A(n_3382),
.Y(n_3632)
);

INVxp67_ASAP7_75t_L g3633 ( 
.A(n_3351),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3444),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3445),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3446),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3448),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3451),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3455),
.Y(n_3639)
);

INVx2_ASAP7_75t_L g3640 ( 
.A(n_3406),
.Y(n_3640)
);

AND2x6_ASAP7_75t_L g3641 ( 
.A(n_3437),
.B(n_3262),
.Y(n_3641)
);

CKINVDCx5p33_ASAP7_75t_R g3642 ( 
.A(n_3338),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3277),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3318),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3411),
.Y(n_3645)
);

OA21x2_ASAP7_75t_L g3646 ( 
.A1(n_3416),
.A2(n_3263),
.B(n_2807),
.Y(n_3646)
);

BUFx2_ASAP7_75t_L g3647 ( 
.A(n_3394),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3414),
.Y(n_3648)
);

OAI22xp5_ASAP7_75t_L g3649 ( 
.A1(n_3290),
.A2(n_2764),
.B1(n_1991),
.B2(n_1992),
.Y(n_3649)
);

INVx3_ASAP7_75t_L g3650 ( 
.A(n_3418),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3426),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3432),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3449),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3469),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_SL g3655 ( 
.A(n_3304),
.B(n_1989),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3394),
.Y(n_3656)
);

CKINVDCx5p33_ASAP7_75t_R g3657 ( 
.A(n_3322),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3299),
.Y(n_3658)
);

OA21x2_ASAP7_75t_L g3659 ( 
.A1(n_3306),
.A2(n_1996),
.B(n_1990),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_SL g3660 ( 
.A(n_3428),
.B(n_1994),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3430),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3463),
.B(n_2457),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3364),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3364),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3391),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3365),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_SL g3667 ( 
.A(n_3350),
.B(n_1997),
.Y(n_3667)
);

INVxp33_ASAP7_75t_L g3668 ( 
.A(n_3433),
.Y(n_3668)
);

BUFx6f_ASAP7_75t_L g3669 ( 
.A(n_3399),
.Y(n_3669)
);

AND2x2_ASAP7_75t_SL g3670 ( 
.A(n_3359),
.B(n_2460),
.Y(n_3670)
);

AND2x4_ASAP7_75t_L g3671 ( 
.A(n_3296),
.B(n_2000),
.Y(n_3671)
);

INVx2_ASAP7_75t_L g3672 ( 
.A(n_3385),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3324),
.B(n_2463),
.Y(n_3673)
);

BUFx6f_ASAP7_75t_L g3674 ( 
.A(n_3362),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3467),
.Y(n_3675)
);

BUFx3_ASAP7_75t_L g3676 ( 
.A(n_3374),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3454),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3387),
.Y(n_3678)
);

OAI22xp5_ASAP7_75t_L g3679 ( 
.A1(n_3372),
.A2(n_2003),
.B1(n_2007),
.B2(n_2005),
.Y(n_3679)
);

XNOR2x2_ASAP7_75t_L g3680 ( 
.A(n_3436),
.B(n_2308),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3450),
.Y(n_3681)
);

NOR2xp33_ASAP7_75t_SL g3682 ( 
.A(n_3276),
.B(n_2123),
.Y(n_3682)
);

BUFx6f_ASAP7_75t_L g3683 ( 
.A(n_3380),
.Y(n_3683)
);

OR2x2_ASAP7_75t_L g3684 ( 
.A(n_3361),
.B(n_2390),
.Y(n_3684)
);

INVx2_ASAP7_75t_L g3685 ( 
.A(n_3443),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3396),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3336),
.B(n_2501),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3386),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3375),
.Y(n_3689)
);

BUFx6f_ASAP7_75t_L g3690 ( 
.A(n_3271),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3466),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3466),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3466),
.Y(n_3693)
);

BUFx6f_ASAP7_75t_L g3694 ( 
.A(n_3271),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3466),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3466),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3466),
.Y(n_3697)
);

BUFx2_ASAP7_75t_L g3698 ( 
.A(n_3404),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3466),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3466),
.Y(n_3700)
);

BUFx6f_ASAP7_75t_L g3701 ( 
.A(n_3271),
.Y(n_3701)
);

AOI22xp5_ASAP7_75t_L g3702 ( 
.A1(n_3421),
.A2(n_2426),
.B1(n_2433),
.B2(n_2396),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3466),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3466),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3523),
.Y(n_3705)
);

INVx3_ASAP7_75t_L g3706 ( 
.A(n_3538),
.Y(n_3706)
);

AND2x4_ASAP7_75t_L g3707 ( 
.A(n_3489),
.B(n_2004),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3571),
.B(n_2008),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3499),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3503),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_3517),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3534),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3583),
.B(n_2012),
.Y(n_3713)
);

NOR2xp33_ASAP7_75t_L g3714 ( 
.A(n_3565),
.B(n_2443),
.Y(n_3714)
);

BUFx3_ASAP7_75t_L g3715 ( 
.A(n_3683),
.Y(n_3715)
);

BUFx6f_ASAP7_75t_L g3716 ( 
.A(n_3538),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3544),
.Y(n_3717)
);

NOR2xp33_ASAP7_75t_L g3718 ( 
.A(n_3588),
.B(n_2444),
.Y(n_3718)
);

NOR2xp33_ASAP7_75t_L g3719 ( 
.A(n_3482),
.B(n_2453),
.Y(n_3719)
);

NOR2xp33_ASAP7_75t_SL g3720 ( 
.A(n_3587),
.B(n_2124),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_SL g3721 ( 
.A(n_3663),
.B(n_2014),
.Y(n_3721)
);

INVx5_ASAP7_75t_L g3722 ( 
.A(n_3669),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_L g3723 ( 
.A(n_3664),
.B(n_2461),
.Y(n_3723)
);

INVx5_ASAP7_75t_L g3724 ( 
.A(n_3669),
.Y(n_3724)
);

BUFx4f_ASAP7_75t_L g3725 ( 
.A(n_3683),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3526),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3527),
.Y(n_3727)
);

CKINVDCx5p33_ASAP7_75t_R g3728 ( 
.A(n_3597),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3525),
.B(n_2015),
.Y(n_3729)
);

INVx2_ASAP7_75t_SL g3730 ( 
.A(n_3511),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3529),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3530),
.B(n_2016),
.Y(n_3732)
);

INVx5_ASAP7_75t_L g3733 ( 
.A(n_3548),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3633),
.B(n_2483),
.Y(n_3734)
);

INVx4_ASAP7_75t_L g3735 ( 
.A(n_3553),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_SL g3736 ( 
.A(n_3656),
.B(n_2017),
.Y(n_3736)
);

NOR2xp33_ASAP7_75t_L g3737 ( 
.A(n_3607),
.B(n_2556),
.Y(n_3737)
);

NOR2x1p5_ASAP7_75t_L g3738 ( 
.A(n_3685),
.B(n_2021),
.Y(n_3738)
);

BUFx3_ASAP7_75t_L g3739 ( 
.A(n_3548),
.Y(n_3739)
);

INVxp33_ASAP7_75t_L g3740 ( 
.A(n_3539),
.Y(n_3740)
);

BUFx10_ASAP7_75t_L g3741 ( 
.A(n_3657),
.Y(n_3741)
);

AND3x1_ASAP7_75t_L g3742 ( 
.A(n_3562),
.B(n_2025),
.C(n_2009),
.Y(n_3742)
);

BUFx2_ASAP7_75t_L g3743 ( 
.A(n_3698),
.Y(n_3743)
);

BUFx6f_ASAP7_75t_L g3744 ( 
.A(n_3549),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3531),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3533),
.Y(n_3746)
);

INVx1_ASAP7_75t_SL g3747 ( 
.A(n_3684),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3537),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3541),
.Y(n_3749)
);

INVx1_ASAP7_75t_SL g3750 ( 
.A(n_3616),
.Y(n_3750)
);

INVx1_ASAP7_75t_SL g3751 ( 
.A(n_3647),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3542),
.Y(n_3752)
);

CKINVDCx5p33_ASAP7_75t_R g3753 ( 
.A(n_3642),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3563),
.B(n_2277),
.Y(n_3754)
);

NAND2xp33_ASAP7_75t_L g3755 ( 
.A(n_3496),
.B(n_2022),
.Y(n_3755)
);

BUFx10_ASAP7_75t_L g3756 ( 
.A(n_3671),
.Y(n_3756)
);

BUFx10_ASAP7_75t_L g3757 ( 
.A(n_3594),
.Y(n_3757)
);

INVx3_ASAP7_75t_L g3758 ( 
.A(n_3549),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3543),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_SL g3760 ( 
.A(n_3615),
.B(n_2023),
.Y(n_3760)
);

NOR2xp33_ASAP7_75t_L g3761 ( 
.A(n_3590),
.B(n_3514),
.Y(n_3761)
);

BUFx4f_ASAP7_75t_L g3762 ( 
.A(n_3674),
.Y(n_3762)
);

BUFx10_ASAP7_75t_L g3763 ( 
.A(n_3675),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3545),
.Y(n_3764)
);

BUFx6f_ASAP7_75t_SL g3765 ( 
.A(n_3670),
.Y(n_3765)
);

NOR2xp33_ASAP7_75t_L g3766 ( 
.A(n_3492),
.B(n_2574),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3567),
.Y(n_3767)
);

BUFx8_ASAP7_75t_SL g3768 ( 
.A(n_3596),
.Y(n_3768)
);

INVx3_ASAP7_75t_L g3769 ( 
.A(n_3552),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3546),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3513),
.B(n_2026),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3550),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_SL g3773 ( 
.A(n_3568),
.B(n_2027),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_SL g3774 ( 
.A(n_3560),
.B(n_2031),
.Y(n_3774)
);

AOI22xp33_ASAP7_75t_L g3775 ( 
.A1(n_3582),
.A2(n_2173),
.B1(n_2891),
.B2(n_2002),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3564),
.B(n_2277),
.Y(n_3776)
);

INVx8_ASAP7_75t_L g3777 ( 
.A(n_3496),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_SL g3778 ( 
.A(n_3617),
.B(n_2032),
.Y(n_3778)
);

AND2x4_ASAP7_75t_L g3779 ( 
.A(n_3601),
.B(n_2033),
.Y(n_3779)
);

INVx1_ASAP7_75t_SL g3780 ( 
.A(n_3687),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3572),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3575),
.Y(n_3782)
);

INVx1_ASAP7_75t_SL g3783 ( 
.A(n_3625),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3478),
.B(n_2037),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3662),
.B(n_2040),
.Y(n_3785)
);

INVx2_ASAP7_75t_SL g3786 ( 
.A(n_3654),
.Y(n_3786)
);

INVxp67_ASAP7_75t_L g3787 ( 
.A(n_3505),
.Y(n_3787)
);

HB1xp67_ASAP7_75t_L g3788 ( 
.A(n_3659),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3551),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3479),
.B(n_2041),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3704),
.B(n_3483),
.Y(n_3791)
);

INVx4_ASAP7_75t_L g3792 ( 
.A(n_3553),
.Y(n_3792)
);

AND2x2_ASAP7_75t_L g3793 ( 
.A(n_3620),
.B(n_2421),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3703),
.B(n_3691),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3554),
.Y(n_3795)
);

INVx4_ASAP7_75t_L g3796 ( 
.A(n_3570),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3692),
.B(n_2042),
.Y(n_3797)
);

NOR2xp33_ASAP7_75t_L g3798 ( 
.A(n_3667),
.B(n_2597),
.Y(n_3798)
);

BUFx8_ASAP7_75t_SL g3799 ( 
.A(n_3528),
.Y(n_3799)
);

INVx2_ASAP7_75t_SL g3800 ( 
.A(n_3580),
.Y(n_3800)
);

INVx4_ASAP7_75t_L g3801 ( 
.A(n_3570),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3555),
.Y(n_3802)
);

NOR2xp33_ASAP7_75t_L g3803 ( 
.A(n_3512),
.B(n_2719),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3693),
.B(n_2043),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3695),
.B(n_2044),
.Y(n_3805)
);

NAND2xp33_ASAP7_75t_SL g3806 ( 
.A(n_3674),
.B(n_2147),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3558),
.Y(n_3807)
);

INVx2_ASAP7_75t_SL g3808 ( 
.A(n_3646),
.Y(n_3808)
);

AND2x4_ASAP7_75t_L g3809 ( 
.A(n_3484),
.B(n_2035),
.Y(n_3809)
);

OAI22xp33_ASAP7_75t_L g3810 ( 
.A1(n_3702),
.A2(n_2780),
.B1(n_2821),
.B2(n_2748),
.Y(n_3810)
);

NOR2x1p5_ASAP7_75t_L g3811 ( 
.A(n_3677),
.B(n_2045),
.Y(n_3811)
);

BUFx2_ASAP7_75t_L g3812 ( 
.A(n_3498),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_SL g3813 ( 
.A(n_3658),
.B(n_2046),
.Y(n_3813)
);

INVx2_ASAP7_75t_L g3814 ( 
.A(n_3579),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3576),
.Y(n_3815)
);

NOR2xp33_ASAP7_75t_L g3816 ( 
.A(n_3495),
.B(n_2849),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3696),
.B(n_2055),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3559),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3591),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3603),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_SL g3821 ( 
.A(n_3661),
.B(n_3507),
.Y(n_3821)
);

NOR2xp33_ASAP7_75t_L g3822 ( 
.A(n_3497),
.B(n_2876),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3561),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3697),
.B(n_2056),
.Y(n_3824)
);

INVx3_ASAP7_75t_L g3825 ( 
.A(n_3552),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3604),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3608),
.Y(n_3827)
);

BUFx10_ASAP7_75t_L g3828 ( 
.A(n_3678),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3566),
.Y(n_3829)
);

INVxp33_ASAP7_75t_L g3830 ( 
.A(n_3481),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3699),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3700),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3500),
.B(n_2057),
.Y(n_3833)
);

NAND2xp33_ASAP7_75t_L g3834 ( 
.A(n_3574),
.B(n_2060),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3644),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_SL g3836 ( 
.A(n_3673),
.B(n_2063),
.Y(n_3836)
);

AOI22xp33_ASAP7_75t_L g3837 ( 
.A1(n_3569),
.A2(n_3509),
.B1(n_3516),
.B2(n_3508),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3494),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3611),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_SL g3840 ( 
.A(n_3487),
.B(n_2064),
.Y(n_3840)
);

NOR2xp33_ASAP7_75t_L g3841 ( 
.A(n_3501),
.B(n_2880),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_SL g3842 ( 
.A(n_3488),
.B(n_2068),
.Y(n_3842)
);

HB1xp67_ASAP7_75t_L g3843 ( 
.A(n_3619),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_SL g3844 ( 
.A(n_3577),
.B(n_2069),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3612),
.Y(n_3845)
);

NOR2xp33_ASAP7_75t_SL g3846 ( 
.A(n_3682),
.B(n_2218),
.Y(n_3846)
);

NAND3xp33_ASAP7_75t_L g3847 ( 
.A(n_3649),
.B(n_2073),
.C(n_2071),
.Y(n_3847)
);

NOR2xp33_ASAP7_75t_L g3848 ( 
.A(n_3502),
.B(n_2075),
.Y(n_3848)
);

AND3x2_ASAP7_75t_L g3849 ( 
.A(n_3524),
.B(n_2604),
.C(n_2579),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3613),
.Y(n_3850)
);

NOR2xp33_ASAP7_75t_L g3851 ( 
.A(n_3504),
.B(n_2077),
.Y(n_3851)
);

AOI22xp33_ASAP7_75t_L g3852 ( 
.A1(n_3672),
.A2(n_2637),
.B1(n_2649),
.B2(n_2627),
.Y(n_3852)
);

INVx4_ASAP7_75t_L g3853 ( 
.A(n_3578),
.Y(n_3853)
);

BUFx6f_ASAP7_75t_L g3854 ( 
.A(n_3690),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3621),
.Y(n_3855)
);

INVx3_ASAP7_75t_L g3856 ( 
.A(n_3690),
.Y(n_3856)
);

INVx5_ASAP7_75t_L g3857 ( 
.A(n_3694),
.Y(n_3857)
);

INVx3_ASAP7_75t_L g3858 ( 
.A(n_3694),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3623),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_SL g3860 ( 
.A(n_3609),
.B(n_2078),
.Y(n_3860)
);

INVx3_ASAP7_75t_L g3861 ( 
.A(n_3701),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3628),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3635),
.Y(n_3863)
);

BUFx3_ASAP7_75t_L g3864 ( 
.A(n_3701),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3485),
.B(n_2081),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_SL g3866 ( 
.A(n_3665),
.B(n_3585),
.Y(n_3866)
);

BUFx6f_ASAP7_75t_L g3867 ( 
.A(n_3578),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_SL g3868 ( 
.A(n_3586),
.B(n_2083),
.Y(n_3868)
);

INVx2_ASAP7_75t_SL g3869 ( 
.A(n_3480),
.Y(n_3869)
);

BUFx10_ASAP7_75t_L g3870 ( 
.A(n_3681),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_3486),
.B(n_2085),
.Y(n_3871)
);

BUFx10_ASAP7_75t_L g3872 ( 
.A(n_3689),
.Y(n_3872)
);

AND2x4_ASAP7_75t_L g3873 ( 
.A(n_3490),
.B(n_2047),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3602),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3606),
.Y(n_3875)
);

BUFx10_ASAP7_75t_L g3876 ( 
.A(n_3491),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3610),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3624),
.Y(n_3878)
);

AND2x4_ASAP7_75t_L g3879 ( 
.A(n_3493),
.B(n_2050),
.Y(n_3879)
);

INVx1_ASAP7_75t_SL g3880 ( 
.A(n_3676),
.Y(n_3880)
);

BUFx3_ASAP7_75t_L g3881 ( 
.A(n_3581),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_SL g3882 ( 
.A(n_3589),
.B(n_2087),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3629),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3634),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3614),
.B(n_2090),
.Y(n_3885)
);

NOR2xp33_ASAP7_75t_L g3886 ( 
.A(n_3540),
.B(n_2094),
.Y(n_3886)
);

INVx3_ASAP7_75t_L g3887 ( 
.A(n_3581),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3641),
.B(n_2100),
.Y(n_3888)
);

AND2x6_ASAP7_75t_L g3889 ( 
.A(n_3518),
.B(n_2051),
.Y(n_3889)
);

INVx3_ASAP7_75t_L g3890 ( 
.A(n_3584),
.Y(n_3890)
);

INVx5_ASAP7_75t_L g3891 ( 
.A(n_3584),
.Y(n_3891)
);

BUFx6f_ASAP7_75t_L g3892 ( 
.A(n_3618),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3636),
.Y(n_3893)
);

BUFx6f_ASAP7_75t_L g3894 ( 
.A(n_3618),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_SL g3895 ( 
.A(n_3592),
.B(n_3598),
.Y(n_3895)
);

OR2x2_ASAP7_75t_L g3896 ( 
.A(n_3679),
.B(n_2102),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_3641),
.B(n_2103),
.Y(n_3897)
);

AND2x4_ASAP7_75t_L g3898 ( 
.A(n_3640),
.B(n_2053),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3637),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_3638),
.Y(n_3900)
);

AOI22xp5_ASAP7_75t_L g3901 ( 
.A1(n_3574),
.A2(n_2227),
.B1(n_2231),
.B2(n_2221),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_SL g3902 ( 
.A(n_3600),
.B(n_2104),
.Y(n_3902)
);

INVx1_ASAP7_75t_SL g3903 ( 
.A(n_3593),
.Y(n_3903)
);

BUFx2_ASAP7_75t_L g3904 ( 
.A(n_3510),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3639),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3622),
.B(n_2108),
.Y(n_3906)
);

INVx3_ASAP7_75t_L g3907 ( 
.A(n_3626),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3536),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3622),
.B(n_2112),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_3573),
.Y(n_3910)
);

INVx2_ASAP7_75t_SL g3911 ( 
.A(n_3645),
.Y(n_3911)
);

INVx2_ASAP7_75t_L g3912 ( 
.A(n_3556),
.Y(n_3912)
);

INVx2_ASAP7_75t_SL g3913 ( 
.A(n_3643),
.Y(n_3913)
);

INVx4_ASAP7_75t_L g3914 ( 
.A(n_3626),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_SL g3915 ( 
.A(n_3627),
.B(n_2115),
.Y(n_3915)
);

INVx1_ASAP7_75t_SL g3916 ( 
.A(n_3532),
.Y(n_3916)
);

INVx2_ASAP7_75t_SL g3917 ( 
.A(n_3506),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3519),
.Y(n_3918)
);

NAND2xp33_ASAP7_75t_L g3919 ( 
.A(n_3520),
.B(n_2122),
.Y(n_3919)
);

OAI21xp33_ASAP7_75t_SL g3920 ( 
.A1(n_3522),
.A2(n_2065),
.B(n_2059),
.Y(n_3920)
);

INVx4_ASAP7_75t_L g3921 ( 
.A(n_3627),
.Y(n_3921)
);

CKINVDCx20_ASAP7_75t_R g3922 ( 
.A(n_3595),
.Y(n_3922)
);

HB1xp67_ASAP7_75t_L g3923 ( 
.A(n_3686),
.Y(n_3923)
);

NOR2xp33_ASAP7_75t_L g3924 ( 
.A(n_3660),
.B(n_2129),
.Y(n_3924)
);

INVx2_ASAP7_75t_SL g3925 ( 
.A(n_3515),
.Y(n_3925)
);

NOR2xp33_ASAP7_75t_L g3926 ( 
.A(n_3605),
.B(n_2131),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3557),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3631),
.B(n_2136),
.Y(n_3928)
);

BUFx6f_ASAP7_75t_L g3929 ( 
.A(n_3630),
.Y(n_3929)
);

INVx2_ASAP7_75t_SL g3930 ( 
.A(n_3521),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3535),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_3648),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3651),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3652),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3630),
.Y(n_3935)
);

AND2x6_ASAP7_75t_L g3936 ( 
.A(n_3688),
.B(n_2067),
.Y(n_3936)
);

BUFx3_ASAP7_75t_L g3937 ( 
.A(n_3632),
.Y(n_3937)
);

BUFx6f_ASAP7_75t_SL g3938 ( 
.A(n_3632),
.Y(n_3938)
);

INVxp33_ASAP7_75t_L g3939 ( 
.A(n_3668),
.Y(n_3939)
);

NOR2xp33_ASAP7_75t_L g3940 ( 
.A(n_3655),
.B(n_2137),
.Y(n_3940)
);

INVx3_ASAP7_75t_L g3941 ( 
.A(n_3547),
.Y(n_3941)
);

BUFx3_ASAP7_75t_L g3942 ( 
.A(n_3650),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3653),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3666),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3680),
.Y(n_3945)
);

INVx1_ASAP7_75t_SL g3946 ( 
.A(n_3599),
.Y(n_3946)
);

INVx2_ASAP7_75t_L g3947 ( 
.A(n_3499),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3523),
.Y(n_3948)
);

INVx5_ASAP7_75t_L g3949 ( 
.A(n_3669),
.Y(n_3949)
);

NOR2xp33_ASAP7_75t_L g3950 ( 
.A(n_3583),
.B(n_2139),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3523),
.Y(n_3951)
);

OR2x2_ASAP7_75t_L g3952 ( 
.A(n_3583),
.B(n_2140),
.Y(n_3952)
);

INVx3_ASAP7_75t_L g3953 ( 
.A(n_3538),
.Y(n_3953)
);

AOI22xp33_ASAP7_75t_L g3954 ( 
.A1(n_3583),
.A2(n_2717),
.B1(n_2736),
.B2(n_2708),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_3499),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3563),
.B(n_2421),
.Y(n_3956)
);

AOI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3571),
.A2(n_2234),
.B1(n_2288),
.B2(n_2233),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3499),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3571),
.B(n_2142),
.Y(n_3959)
);

INVx3_ASAP7_75t_L g3960 ( 
.A(n_3538),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3523),
.Y(n_3961)
);

INVx3_ASAP7_75t_L g3962 ( 
.A(n_3538),
.Y(n_3962)
);

INVx3_ASAP7_75t_L g3963 ( 
.A(n_3538),
.Y(n_3963)
);

AND2x4_ASAP7_75t_L g3964 ( 
.A(n_3489),
.B(n_2070),
.Y(n_3964)
);

NOR2xp33_ASAP7_75t_L g3965 ( 
.A(n_3583),
.B(n_2148),
.Y(n_3965)
);

NAND2xp33_ASAP7_75t_L g3966 ( 
.A(n_3583),
.B(n_2149),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3571),
.B(n_2150),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3523),
.Y(n_3968)
);

BUFx3_ASAP7_75t_L g3969 ( 
.A(n_3683),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3523),
.Y(n_3970)
);

AND2x6_ASAP7_75t_L g3971 ( 
.A(n_3582),
.B(n_2084),
.Y(n_3971)
);

INVx1_ASAP7_75t_SL g3972 ( 
.A(n_3511),
.Y(n_3972)
);

AOI22xp33_ASAP7_75t_L g3973 ( 
.A1(n_3583),
.A2(n_2771),
.B1(n_2776),
.B2(n_2755),
.Y(n_3973)
);

INVx4_ASAP7_75t_SL g3974 ( 
.A(n_3669),
.Y(n_3974)
);

INVx3_ASAP7_75t_L g3975 ( 
.A(n_3538),
.Y(n_3975)
);

INVx4_ASAP7_75t_SL g3976 ( 
.A(n_3669),
.Y(n_3976)
);

BUFx4f_ASAP7_75t_L g3977 ( 
.A(n_3669),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3499),
.Y(n_3978)
);

INVx1_ASAP7_75t_SL g3979 ( 
.A(n_3511),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3523),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3523),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3499),
.Y(n_3982)
);

INVx3_ASAP7_75t_L g3983 ( 
.A(n_3538),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3571),
.B(n_2156),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3571),
.B(n_2157),
.Y(n_3985)
);

AOI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_3571),
.A2(n_2377),
.B1(n_2382),
.B2(n_2356),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3571),
.B(n_2160),
.Y(n_3987)
);

OR2x2_ASAP7_75t_L g3988 ( 
.A(n_3583),
.B(n_2161),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_3499),
.Y(n_3989)
);

BUFx6f_ASAP7_75t_L g3990 ( 
.A(n_3538),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3571),
.B(n_2165),
.Y(n_3991)
);

INVx2_ASAP7_75t_SL g3992 ( 
.A(n_3511),
.Y(n_3992)
);

BUFx10_ASAP7_75t_L g3993 ( 
.A(n_3669),
.Y(n_3993)
);

BUFx3_ASAP7_75t_L g3994 ( 
.A(n_3683),
.Y(n_3994)
);

INVx2_ASAP7_75t_L g3995 ( 
.A(n_3499),
.Y(n_3995)
);

BUFx4f_ASAP7_75t_L g3996 ( 
.A(n_3669),
.Y(n_3996)
);

OR2x2_ASAP7_75t_L g3997 ( 
.A(n_3583),
.B(n_2166),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3523),
.Y(n_3998)
);

BUFx6f_ASAP7_75t_L g3999 ( 
.A(n_3538),
.Y(n_3999)
);

INVxp67_ASAP7_75t_SL g4000 ( 
.A(n_3508),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3523),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3523),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3523),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3571),
.B(n_2167),
.Y(n_4004)
);

INVx3_ASAP7_75t_L g4005 ( 
.A(n_3538),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3705),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_3950),
.B(n_3965),
.Y(n_4007)
);

INVxp67_ASAP7_75t_L g4008 ( 
.A(n_3754),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3719),
.B(n_2168),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3708),
.B(n_2169),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3714),
.B(n_2475),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3959),
.B(n_2170),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3967),
.B(n_2171),
.Y(n_4013)
);

NOR2xp33_ASAP7_75t_L g4014 ( 
.A(n_3780),
.B(n_2388),
.Y(n_4014)
);

OAI22xp5_ASAP7_75t_L g4015 ( 
.A1(n_3837),
.A2(n_2429),
.B1(n_2451),
.B2(n_2401),
.Y(n_4015)
);

AOI22xp33_ASAP7_75t_L g4016 ( 
.A1(n_3798),
.A2(n_2513),
.B1(n_2515),
.B2(n_2471),
.Y(n_4016)
);

NOR3xp33_ASAP7_75t_L g4017 ( 
.A(n_3806),
.B(n_2174),
.C(n_2172),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3726),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3984),
.B(n_2178),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3709),
.Y(n_4020)
);

BUFx6f_ASAP7_75t_SL g4021 ( 
.A(n_3993),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3985),
.B(n_2180),
.Y(n_4022)
);

AOI22xp33_ASAP7_75t_L g4023 ( 
.A1(n_3945),
.A2(n_2563),
.B1(n_2575),
.B2(n_2517),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3987),
.B(n_3991),
.Y(n_4024)
);

NOR2x1p5_ASAP7_75t_L g4025 ( 
.A(n_3715),
.B(n_3969),
.Y(n_4025)
);

OAI221xp5_ASAP7_75t_L g4026 ( 
.A1(n_4004),
.A2(n_2089),
.B1(n_2092),
.B2(n_2088),
.C(n_2086),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_L g4027 ( 
.A(n_3718),
.B(n_2181),
.Y(n_4027)
);

BUFx2_ASAP7_75t_L g4028 ( 
.A(n_3743),
.Y(n_4028)
);

NOR2xp33_ASAP7_75t_L g4029 ( 
.A(n_3740),
.B(n_2644),
.Y(n_4029)
);

INVx5_ASAP7_75t_L g4030 ( 
.A(n_3777),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3761),
.B(n_2182),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3710),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_4000),
.B(n_2187),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3713),
.B(n_2189),
.Y(n_4034)
);

AOI22xp5_ASAP7_75t_L g4035 ( 
.A1(n_3808),
.A2(n_2727),
.B1(n_2734),
.B2(n_2702),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3727),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_3711),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3712),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_3717),
.Y(n_4039)
);

AND2x4_ASAP7_75t_L g4040 ( 
.A(n_3974),
.B(n_2095),
.Y(n_4040)
);

NOR2xp33_ASAP7_75t_L g4041 ( 
.A(n_3747),
.B(n_3787),
.Y(n_4041)
);

NOR3xp33_ASAP7_75t_L g4042 ( 
.A(n_3926),
.B(n_2193),
.C(n_2191),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3731),
.Y(n_4043)
);

NOR3xp33_ASAP7_75t_L g4044 ( 
.A(n_3810),
.B(n_2195),
.C(n_2194),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3766),
.B(n_2196),
.Y(n_4045)
);

BUFx6f_ASAP7_75t_L g4046 ( 
.A(n_3716),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3745),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3746),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_3732),
.B(n_2198),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_SL g4050 ( 
.A(n_3750),
.B(n_2783),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3729),
.B(n_2200),
.Y(n_4051)
);

AOI21xp5_ASAP7_75t_L g4052 ( 
.A1(n_3908),
.A2(n_2106),
.B(n_2098),
.Y(n_4052)
);

HB1xp67_ASAP7_75t_L g4053 ( 
.A(n_3730),
.Y(n_4053)
);

AOI22xp5_ASAP7_75t_L g4054 ( 
.A1(n_3788),
.A2(n_2812),
.B1(n_2852),
.B2(n_2794),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_SL g4055 ( 
.A(n_3725),
.B(n_2862),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_SL g4056 ( 
.A(n_3846),
.B(n_2878),
.Y(n_4056)
);

INVx2_ASAP7_75t_L g4057 ( 
.A(n_3767),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_3947),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3771),
.B(n_3816),
.Y(n_4059)
);

INVx2_ASAP7_75t_L g4060 ( 
.A(n_3955),
.Y(n_4060)
);

NOR2xp33_ASAP7_75t_SL g4061 ( 
.A(n_3728),
.B(n_2886),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_SL g4062 ( 
.A(n_3762),
.B(n_2887),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3822),
.B(n_3841),
.Y(n_4063)
);

CKINVDCx20_ASAP7_75t_R g4064 ( 
.A(n_3753),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3952),
.B(n_2203),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_SL g4066 ( 
.A(n_3988),
.B(n_2904),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_3748),
.Y(n_4067)
);

NAND3xp33_ASAP7_75t_L g4068 ( 
.A(n_3966),
.B(n_2205),
.C(n_2204),
.Y(n_4068)
);

AOI22xp33_ASAP7_75t_L g4069 ( 
.A1(n_3971),
.A2(n_2923),
.B1(n_2932),
.B2(n_2919),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_3958),
.Y(n_4070)
);

INVxp67_ASAP7_75t_L g4071 ( 
.A(n_3956),
.Y(n_4071)
);

NOR2xp33_ASAP7_75t_L g4072 ( 
.A(n_3997),
.B(n_2940),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_SL g4073 ( 
.A(n_3992),
.B(n_2945),
.Y(n_4073)
);

INVx2_ASAP7_75t_L g4074 ( 
.A(n_3978),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3749),
.Y(n_4075)
);

A2O1A1Ixp33_ASAP7_75t_L g4076 ( 
.A1(n_3803),
.A2(n_2113),
.B(n_2114),
.C(n_2107),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_3752),
.B(n_2206),
.Y(n_4077)
);

INVx8_ASAP7_75t_L g4078 ( 
.A(n_3722),
.Y(n_4078)
);

INVx3_ASAP7_75t_L g4079 ( 
.A(n_3867),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3759),
.Y(n_4080)
);

CKINVDCx5p33_ASAP7_75t_R g4081 ( 
.A(n_3768),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3764),
.B(n_2208),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3770),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3772),
.B(n_2210),
.Y(n_4084)
);

INVxp67_ASAP7_75t_L g4085 ( 
.A(n_3776),
.Y(n_4085)
);

OAI21xp5_ASAP7_75t_L g4086 ( 
.A1(n_3931),
.A2(n_2118),
.B(n_2117),
.Y(n_4086)
);

NOR2xp33_ASAP7_75t_L g4087 ( 
.A(n_3957),
.B(n_3986),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_L g4088 ( 
.A(n_3789),
.B(n_2213),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_SL g4089 ( 
.A(n_3722),
.B(n_2972),
.Y(n_4089)
);

NOR2xp33_ASAP7_75t_L g4090 ( 
.A(n_3734),
.B(n_3003),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3795),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3802),
.Y(n_4092)
);

OR2x2_ASAP7_75t_L g4093 ( 
.A(n_3972),
.B(n_3979),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3724),
.B(n_2475),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3807),
.Y(n_4095)
);

INVx2_ASAP7_75t_L g4096 ( 
.A(n_3982),
.Y(n_4096)
);

NOR2xp33_ASAP7_75t_L g4097 ( 
.A(n_3880),
.B(n_2217),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3989),
.Y(n_4098)
);

INVx2_ASAP7_75t_SL g4099 ( 
.A(n_3724),
.Y(n_4099)
);

INVx2_ASAP7_75t_L g4100 ( 
.A(n_3995),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_3831),
.B(n_2219),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_3832),
.B(n_2222),
.Y(n_4102)
);

INVxp33_ASAP7_75t_L g4103 ( 
.A(n_3977),
.Y(n_4103)
);

NOR3xp33_ASAP7_75t_L g4104 ( 
.A(n_3847),
.B(n_2225),
.C(n_2223),
.Y(n_4104)
);

O2A1O1Ixp5_ASAP7_75t_L g4105 ( 
.A1(n_3885),
.A2(n_2830),
.B(n_2842),
.C(n_2789),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_3781),
.Y(n_4106)
);

NOR2xp33_ASAP7_75t_L g4107 ( 
.A(n_3737),
.B(n_3946),
.Y(n_4107)
);

CKINVDCx16_ASAP7_75t_R g4108 ( 
.A(n_3741),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3948),
.B(n_2228),
.Y(n_4109)
);

NOR2xp33_ASAP7_75t_L g4110 ( 
.A(n_3916),
.B(n_2230),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_3951),
.B(n_2232),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_SL g4112 ( 
.A(n_3949),
.B(n_2237),
.Y(n_4112)
);

NOR2xp33_ASAP7_75t_L g4113 ( 
.A(n_3896),
.B(n_2238),
.Y(n_4113)
);

O2A1O1Ixp33_ASAP7_75t_L g4114 ( 
.A1(n_3920),
.A2(n_2126),
.B(n_2128),
.C(n_2119),
.Y(n_4114)
);

INVx2_ASAP7_75t_L g4115 ( 
.A(n_3782),
.Y(n_4115)
);

BUFx12f_ASAP7_75t_L g4116 ( 
.A(n_3757),
.Y(n_4116)
);

NAND3xp33_ASAP7_75t_SL g4117 ( 
.A(n_3901),
.B(n_2244),
.C(n_2243),
.Y(n_4117)
);

CKINVDCx5p33_ASAP7_75t_R g4118 ( 
.A(n_3799),
.Y(n_4118)
);

BUFx5_ASAP7_75t_L g4119 ( 
.A(n_3927),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_SL g4120 ( 
.A(n_3949),
.B(n_2246),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3961),
.B(n_2249),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3968),
.Y(n_4122)
);

NOR3xp33_ASAP7_75t_L g4123 ( 
.A(n_3860),
.B(n_2253),
.C(n_2252),
.Y(n_4123)
);

INVx2_ASAP7_75t_L g4124 ( 
.A(n_3814),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_3819),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_3970),
.B(n_2255),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_3820),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_3980),
.B(n_2258),
.Y(n_4128)
);

AND2x2_ASAP7_75t_L g4129 ( 
.A(n_3723),
.B(n_2594),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3981),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3998),
.B(n_2259),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_4001),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_4002),
.B(n_2261),
.Y(n_4133)
);

INVx3_ASAP7_75t_L g4134 ( 
.A(n_3867),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4003),
.B(n_2262),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_SL g4136 ( 
.A(n_3996),
.B(n_2268),
.Y(n_4136)
);

AO22x2_ASAP7_75t_L g4137 ( 
.A1(n_3751),
.A2(n_2132),
.B1(n_2133),
.B2(n_2130),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3791),
.B(n_2269),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_SL g4139 ( 
.A(n_3756),
.B(n_2270),
.Y(n_4139)
);

INVxp67_ASAP7_75t_SL g4140 ( 
.A(n_3923),
.Y(n_4140)
);

INVx3_ASAP7_75t_L g4141 ( 
.A(n_3892),
.Y(n_4141)
);

NOR2xp33_ASAP7_75t_L g4142 ( 
.A(n_3830),
.B(n_2276),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3794),
.B(n_2278),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_3826),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3835),
.Y(n_4145)
);

OR2x2_ASAP7_75t_L g4146 ( 
.A(n_3774),
.B(n_3773),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_3848),
.B(n_2279),
.Y(n_4147)
);

INVxp33_ASAP7_75t_L g4148 ( 
.A(n_3793),
.Y(n_4148)
);

INVx2_ASAP7_75t_L g4149 ( 
.A(n_3827),
.Y(n_4149)
);

INVx5_ASAP7_75t_L g4150 ( 
.A(n_3777),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_3851),
.B(n_2282),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_3918),
.B(n_2283),
.Y(n_4152)
);

NOR2xp33_ASAP7_75t_L g4153 ( 
.A(n_3760),
.B(n_2284),
.Y(n_4153)
);

INVx2_ASAP7_75t_L g4154 ( 
.A(n_3845),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_3775),
.B(n_3862),
.Y(n_4155)
);

NOR2xp67_ASAP7_75t_L g4156 ( 
.A(n_3891),
.B(n_1804),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_3971),
.B(n_3843),
.Y(n_4157)
);

NOR2xp33_ASAP7_75t_L g4158 ( 
.A(n_3886),
.B(n_2291),
.Y(n_4158)
);

NOR2xp33_ASAP7_75t_L g4159 ( 
.A(n_3869),
.B(n_2292),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_3971),
.B(n_3839),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_3786),
.B(n_2294),
.Y(n_4161)
);

NOR3xp33_ASAP7_75t_L g4162 ( 
.A(n_3888),
.B(n_2298),
.C(n_2296),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_SL g4163 ( 
.A(n_3833),
.B(n_3994),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_3850),
.B(n_2300),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_3818),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_3855),
.B(n_2302),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_SL g4167 ( 
.A(n_3910),
.B(n_3917),
.Y(n_4167)
);

INVx2_ASAP7_75t_L g4168 ( 
.A(n_3859),
.Y(n_4168)
);

NOR2xp33_ASAP7_75t_L g4169 ( 
.A(n_3783),
.B(n_2303),
.Y(n_4169)
);

CKINVDCx5p33_ASAP7_75t_R g4170 ( 
.A(n_3765),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_SL g4171 ( 
.A(n_3928),
.B(n_2304),
.Y(n_4171)
);

NOR3xp33_ASAP7_75t_L g4172 ( 
.A(n_3897),
.B(n_2306),
.C(n_2305),
.Y(n_4172)
);

AND2x2_ASAP7_75t_L g4173 ( 
.A(n_3976),
.B(n_2594),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_SL g4174 ( 
.A(n_3924),
.B(n_2307),
.Y(n_4174)
);

NOR2xp33_ASAP7_75t_L g4175 ( 
.A(n_3939),
.B(n_2309),
.Y(n_4175)
);

NOR2xp33_ASAP7_75t_L g4176 ( 
.A(n_3778),
.B(n_2312),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3823),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_3863),
.B(n_2314),
.Y(n_4178)
);

A2O1A1Ixp33_ASAP7_75t_L g4179 ( 
.A1(n_3940),
.A2(n_2143),
.B(n_2146),
.C(n_2141),
.Y(n_4179)
);

INVx2_ASAP7_75t_L g4180 ( 
.A(n_3878),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_3829),
.B(n_2316),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_SL g4182 ( 
.A(n_3884),
.B(n_2318),
.Y(n_4182)
);

INVx4_ASAP7_75t_L g4183 ( 
.A(n_3891),
.Y(n_4183)
);

BUFx6f_ASAP7_75t_L g4184 ( 
.A(n_3716),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_3874),
.B(n_2320),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3875),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_SL g4187 ( 
.A(n_3893),
.B(n_2321),
.Y(n_4187)
);

INVx2_ASAP7_75t_L g4188 ( 
.A(n_3900),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_SL g4189 ( 
.A(n_3784),
.B(n_3790),
.Y(n_4189)
);

NOR2xp33_ASAP7_75t_L g4190 ( 
.A(n_3785),
.B(n_2324),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_3877),
.B(n_2327),
.Y(n_4191)
);

HB1xp67_ASAP7_75t_L g4192 ( 
.A(n_3744),
.Y(n_4192)
);

AND2x2_ASAP7_75t_L g4193 ( 
.A(n_3800),
.B(n_2617),
.Y(n_4193)
);

AOI22xp33_ASAP7_75t_L g4194 ( 
.A1(n_3889),
.A2(n_2872),
.B1(n_2888),
.B2(n_2845),
.Y(n_4194)
);

INVxp67_ASAP7_75t_L g4195 ( 
.A(n_3892),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_3903),
.B(n_2617),
.Y(n_4196)
);

OAI22xp5_ASAP7_75t_L g4197 ( 
.A1(n_3912),
.A2(n_2330),
.B1(n_2337),
.B2(n_2328),
.Y(n_4197)
);

O2A1O1Ixp33_ASAP7_75t_L g4198 ( 
.A1(n_3919),
.A2(n_2153),
.B(n_2154),
.C(n_2151),
.Y(n_4198)
);

HB1xp67_ASAP7_75t_L g4199 ( 
.A(n_3744),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_3883),
.B(n_2340),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_3899),
.B(n_2343),
.Y(n_4201)
);

NOR2xp33_ASAP7_75t_L g4202 ( 
.A(n_3797),
.B(n_2344),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_3905),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_3815),
.Y(n_4204)
);

INVx8_ASAP7_75t_L g4205 ( 
.A(n_3733),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_3838),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_3944),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_3889),
.B(n_2345),
.Y(n_4208)
);

AOI22xp33_ASAP7_75t_L g4209 ( 
.A1(n_3889),
.A2(n_2907),
.B1(n_2934),
.B2(n_2902),
.Y(n_4209)
);

NOR2xp33_ASAP7_75t_L g4210 ( 
.A(n_3804),
.B(n_2346),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_3805),
.B(n_2347),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_3817),
.B(n_2348),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_SL g4213 ( 
.A(n_3824),
.B(n_2352),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_3865),
.B(n_2354),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_3871),
.B(n_2357),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_SL g4216 ( 
.A(n_3906),
.B(n_2361),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_3895),
.B(n_2365),
.Y(n_4217)
);

INVx2_ASAP7_75t_SL g4218 ( 
.A(n_3894),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_3913),
.Y(n_4219)
);

NAND3xp33_ASAP7_75t_L g4220 ( 
.A(n_3954),
.B(n_3973),
.C(n_3755),
.Y(n_4220)
);

BUFx2_ASAP7_75t_L g4221 ( 
.A(n_3854),
.Y(n_4221)
);

AOI221xp5_ASAP7_75t_L g4222 ( 
.A1(n_3742),
.A2(n_2164),
.B1(n_2184),
.B2(n_2163),
.C(n_2155),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_3852),
.B(n_2366),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_3932),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3809),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_3866),
.B(n_2368),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_3836),
.B(n_2370),
.Y(n_4227)
);

OR2x2_ASAP7_75t_L g4228 ( 
.A(n_3909),
.B(n_2371),
.Y(n_4228)
);

INVx2_ASAP7_75t_L g4229 ( 
.A(n_3933),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_3821),
.B(n_2372),
.Y(n_4230)
);

OAI221xp5_ASAP7_75t_L g4231 ( 
.A1(n_3840),
.A2(n_2192),
.B1(n_2197),
.B2(n_2190),
.C(n_2186),
.Y(n_4231)
);

CKINVDCx5p33_ASAP7_75t_R g4232 ( 
.A(n_3938),
.Y(n_4232)
);

INVx2_ASAP7_75t_SL g4233 ( 
.A(n_3894),
.Y(n_4233)
);

AOI22xp5_ASAP7_75t_L g4234 ( 
.A1(n_3721),
.A2(n_2378),
.B1(n_2379),
.B2(n_2376),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_3813),
.B(n_2381),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_3736),
.B(n_3868),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_SL g4237 ( 
.A(n_3720),
.B(n_2385),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_SL g4238 ( 
.A(n_3929),
.B(n_2389),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_3873),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_3879),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_3882),
.B(n_2398),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_SL g4242 ( 
.A(n_3929),
.B(n_2400),
.Y(n_4242)
);

INVx2_ASAP7_75t_L g4243 ( 
.A(n_3898),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_3934),
.B(n_2402),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3943),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_3881),
.B(n_2671),
.Y(n_4246)
);

NOR2xp33_ASAP7_75t_R g4247 ( 
.A(n_3922),
.B(n_3834),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_3911),
.Y(n_4248)
);

INVx2_ASAP7_75t_L g4249 ( 
.A(n_3779),
.Y(n_4249)
);

BUFx5_ASAP7_75t_L g4250 ( 
.A(n_3876),
.Y(n_4250)
);

BUFx2_ASAP7_75t_L g4251 ( 
.A(n_3854),
.Y(n_4251)
);

INVx2_ASAP7_75t_L g4252 ( 
.A(n_3935),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_3707),
.Y(n_4253)
);

NOR2xp33_ASAP7_75t_L g4254 ( 
.A(n_3842),
.B(n_2403),
.Y(n_4254)
);

NOR2xp67_ASAP7_75t_L g4255 ( 
.A(n_3735),
.B(n_3792),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_3902),
.B(n_2405),
.Y(n_4256)
);

INVx2_ASAP7_75t_L g4257 ( 
.A(n_3964),
.Y(n_4257)
);

INVx2_ASAP7_75t_L g4258 ( 
.A(n_3941),
.Y(n_4258)
);

NAND2xp5_ASAP7_75t_L g4259 ( 
.A(n_3844),
.B(n_2406),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3925),
.Y(n_4260)
);

CKINVDCx14_ASAP7_75t_R g4261 ( 
.A(n_3812),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_3887),
.B(n_2407),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_3890),
.B(n_2408),
.Y(n_4263)
);

AOI22xp33_ASAP7_75t_L g4264 ( 
.A1(n_3936),
.A2(n_3811),
.B1(n_3915),
.B2(n_3738),
.Y(n_4264)
);

NAND3x1_ASAP7_75t_L g4265 ( 
.A(n_3706),
.B(n_2202),
.C(n_2201),
.Y(n_4265)
);

INVx3_ASAP7_75t_L g4266 ( 
.A(n_3990),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_3930),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_3907),
.B(n_2410),
.Y(n_4268)
);

NOR2xp33_ASAP7_75t_L g4269 ( 
.A(n_3796),
.B(n_2412),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_SL g4270 ( 
.A(n_3801),
.B(n_2413),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_3853),
.B(n_2418),
.Y(n_4271)
);

INVxp67_ASAP7_75t_L g4272 ( 
.A(n_3990),
.Y(n_4272)
);

NOR2xp33_ASAP7_75t_L g4273 ( 
.A(n_3914),
.B(n_2420),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_3921),
.B(n_2422),
.Y(n_4274)
);

NOR2xp33_ASAP7_75t_L g4275 ( 
.A(n_3937),
.B(n_2424),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3942),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_3999),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_3758),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_3999),
.Y(n_4279)
);

NAND2x1p5_ASAP7_75t_L g4280 ( 
.A(n_3733),
.B(n_2207),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_3769),
.B(n_2431),
.Y(n_4281)
);

INVx2_ASAP7_75t_SL g4282 ( 
.A(n_3857),
.Y(n_4282)
);

INVx2_ASAP7_75t_L g4283 ( 
.A(n_3825),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_SL g4284 ( 
.A(n_3857),
.B(n_2432),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_3856),
.B(n_2434),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_3858),
.B(n_2436),
.Y(n_4286)
);

NOR3xp33_ASAP7_75t_L g4287 ( 
.A(n_3861),
.B(n_2442),
.C(n_2441),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_3953),
.B(n_2448),
.Y(n_4288)
);

BUFx6f_ASAP7_75t_L g4289 ( 
.A(n_3739),
.Y(n_4289)
);

AND2x2_ASAP7_75t_L g4290 ( 
.A(n_3864),
.B(n_2671),
.Y(n_4290)
);

INVxp67_ASAP7_75t_L g4291 ( 
.A(n_3936),
.Y(n_4291)
);

AOI22xp5_ASAP7_75t_L g4292 ( 
.A1(n_3936),
.A2(n_2454),
.B1(n_2458),
.B2(n_2449),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_SL g4293 ( 
.A(n_3960),
.B(n_3962),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_3963),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_3975),
.B(n_2459),
.Y(n_4295)
);

AND2x6_ASAP7_75t_L g4296 ( 
.A(n_3983),
.B(n_2211),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_SL g4297 ( 
.A(n_4005),
.B(n_2465),
.Y(n_4297)
);

INVx2_ASAP7_75t_L g4298 ( 
.A(n_3849),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_3872),
.B(n_2466),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_3763),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_3828),
.B(n_2476),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_SL g4302 ( 
.A(n_3870),
.B(n_2477),
.Y(n_4302)
);

AND2x4_ASAP7_75t_L g4303 ( 
.A(n_3904),
.B(n_2214),
.Y(n_4303)
);

NAND3xp33_ASAP7_75t_L g4304 ( 
.A(n_3950),
.B(n_2480),
.C(n_2479),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_3950),
.B(n_2481),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_3709),
.Y(n_4306)
);

HB1xp67_ASAP7_75t_L g4307 ( 
.A(n_3743),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_3950),
.B(n_2484),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_3950),
.B(n_2485),
.Y(n_4309)
);

AOI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_4000),
.A2(n_2242),
.B(n_2239),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_3714),
.B(n_2675),
.Y(n_4311)
);

INVx2_ASAP7_75t_SL g4312 ( 
.A(n_3722),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_3950),
.B(n_2486),
.Y(n_4313)
);

AOI22xp5_ASAP7_75t_L g4314 ( 
.A1(n_3950),
.A2(n_2492),
.B1(n_2493),
.B2(n_2488),
.Y(n_4314)
);

AND2x6_ASAP7_75t_L g4315 ( 
.A(n_3918),
.B(n_2251),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_L g4316 ( 
.A(n_3950),
.B(n_2494),
.Y(n_4316)
);

AOI22xp5_ASAP7_75t_L g4317 ( 
.A1(n_3950),
.A2(n_2499),
.B1(n_2500),
.B2(n_2495),
.Y(n_4317)
);

INVx4_ASAP7_75t_L g4318 ( 
.A(n_3722),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_SL g4319 ( 
.A(n_3761),
.B(n_2503),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_3705),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_3709),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_3950),
.B(n_2506),
.Y(n_4322)
);

NAND3xp33_ASAP7_75t_L g4323 ( 
.A(n_3950),
.B(n_2510),
.C(n_2508),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_3705),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_3950),
.B(n_2511),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_SL g4326 ( 
.A(n_3761),
.B(n_2512),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_3950),
.B(n_2514),
.Y(n_4327)
);

AOI22xp5_ASAP7_75t_L g4328 ( 
.A1(n_3950),
.A2(n_2521),
.B1(n_2522),
.B2(n_2520),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_SL g4329 ( 
.A(n_3761),
.B(n_2523),
.Y(n_4329)
);

NOR2xp33_ASAP7_75t_L g4330 ( 
.A(n_3780),
.B(n_2526),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_3950),
.B(n_2528),
.Y(n_4331)
);

NOR3xp33_ASAP7_75t_L g4332 ( 
.A(n_3806),
.B(n_2532),
.C(n_2530),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_3950),
.B(n_2533),
.Y(n_4333)
);

OR2x2_ASAP7_75t_L g4334 ( 
.A(n_3747),
.B(n_2534),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_3950),
.B(n_2536),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_3705),
.Y(n_4336)
);

AO221x1_ASAP7_75t_L g4337 ( 
.A1(n_3810),
.A2(n_2263),
.B1(n_2265),
.B2(n_2260),
.C(n_2256),
.Y(n_4337)
);

NAND2xp33_ASAP7_75t_L g4338 ( 
.A(n_3889),
.B(n_2539),
.Y(n_4338)
);

INVx2_ASAP7_75t_SL g4339 ( 
.A(n_3722),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_3950),
.B(n_2542),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_SL g4341 ( 
.A(n_3761),
.B(n_2545),
.Y(n_4341)
);

INVx2_ASAP7_75t_L g4342 ( 
.A(n_3709),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_3950),
.B(n_2546),
.Y(n_4343)
);

INVxp67_ASAP7_75t_SL g4344 ( 
.A(n_4000),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_3950),
.B(n_2547),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_3950),
.B(n_2548),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_3709),
.Y(n_4347)
);

AOI21xp5_ASAP7_75t_L g4348 ( 
.A1(n_4000),
.A2(n_2267),
.B(n_2266),
.Y(n_4348)
);

NOR2xp33_ASAP7_75t_SL g4349 ( 
.A(n_3728),
.B(n_2675),
.Y(n_4349)
);

NAND2xp33_ASAP7_75t_L g4350 ( 
.A(n_3889),
.B(n_2550),
.Y(n_4350)
);

INVx2_ASAP7_75t_SL g4351 ( 
.A(n_3722),
.Y(n_4351)
);

AOI22xp33_ASAP7_75t_L g4352 ( 
.A1(n_3950),
.A2(n_2971),
.B1(n_2967),
.B2(n_2273),
.Y(n_4352)
);

NOR2xp67_ASAP7_75t_L g4353 ( 
.A(n_3722),
.B(n_1806),
.Y(n_4353)
);

NOR2xp33_ASAP7_75t_L g4354 ( 
.A(n_3780),
.B(n_2554),
.Y(n_4354)
);

CKINVDCx5p33_ASAP7_75t_R g4355 ( 
.A(n_3728),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_3709),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_3709),
.Y(n_4357)
);

OAI221xp5_ASAP7_75t_L g4358 ( 
.A1(n_3950),
.A2(n_2286),
.B1(n_2289),
.B2(n_2274),
.C(n_2271),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_3714),
.B(n_2760),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_L g4360 ( 
.A(n_3950),
.B(n_2555),
.Y(n_4360)
);

OR2x6_ASAP7_75t_L g4361 ( 
.A(n_3777),
.B(n_2297),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_L g4362 ( 
.A(n_3950),
.B(n_2558),
.Y(n_4362)
);

INVxp67_ASAP7_75t_L g4363 ( 
.A(n_3754),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_3705),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_4007),
.B(n_2559),
.Y(n_4365)
);

AOI22xp33_ASAP7_75t_L g4366 ( 
.A1(n_4087),
.A2(n_2310),
.B1(n_2311),
.B2(n_2299),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4020),
.Y(n_4367)
);

BUFx3_ASAP7_75t_L g4368 ( 
.A(n_4078),
.Y(n_4368)
);

BUFx3_ASAP7_75t_L g4369 ( 
.A(n_4078),
.Y(n_4369)
);

HB1xp67_ASAP7_75t_L g4370 ( 
.A(n_4307),
.Y(n_4370)
);

INVxp33_ASAP7_75t_L g4371 ( 
.A(n_4093),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4006),
.Y(n_4372)
);

AOI22xp33_ASAP7_75t_L g4373 ( 
.A1(n_4063),
.A2(n_2317),
.B1(n_2319),
.B2(n_2315),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_4059),
.B(n_2560),
.Y(n_4374)
);

NAND2xp33_ASAP7_75t_SL g4375 ( 
.A(n_4247),
.B(n_4355),
.Y(n_4375)
);

BUFx6f_ASAP7_75t_L g4376 ( 
.A(n_4046),
.Y(n_4376)
);

AND2x6_ASAP7_75t_L g4377 ( 
.A(n_4024),
.B(n_2322),
.Y(n_4377)
);

AND2x4_ASAP7_75t_L g4378 ( 
.A(n_4025),
.B(n_2323),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4018),
.Y(n_4379)
);

INVx2_ASAP7_75t_L g4380 ( 
.A(n_4032),
.Y(n_4380)
);

NAND2xp33_ASAP7_75t_L g4381 ( 
.A(n_4250),
.B(n_2561),
.Y(n_4381)
);

INVx5_ASAP7_75t_L g4382 ( 
.A(n_4205),
.Y(n_4382)
);

BUFx3_ASAP7_75t_L g4383 ( 
.A(n_4205),
.Y(n_4383)
);

INVx4_ASAP7_75t_L g4384 ( 
.A(n_4046),
.Y(n_4384)
);

AND2x4_ASAP7_75t_L g4385 ( 
.A(n_4318),
.B(n_2325),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_L g4386 ( 
.A(n_4107),
.B(n_2562),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_4031),
.B(n_2564),
.Y(n_4387)
);

AOI22xp5_ASAP7_75t_L g4388 ( 
.A1(n_4158),
.A2(n_2566),
.B1(n_2568),
.B2(n_2565),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_4037),
.Y(n_4389)
);

A2O1A1Ixp33_ASAP7_75t_L g4390 ( 
.A1(n_4113),
.A2(n_2332),
.B(n_2335),
.C(n_2326),
.Y(n_4390)
);

BUFx6f_ASAP7_75t_L g4391 ( 
.A(n_4184),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4036),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4011),
.B(n_2760),
.Y(n_4393)
);

INVx3_ASAP7_75t_L g4394 ( 
.A(n_4289),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_4038),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_SL g4396 ( 
.A(n_4041),
.B(n_2569),
.Y(n_4396)
);

AO22x1_ASAP7_75t_L g4397 ( 
.A1(n_4090),
.A2(n_2571),
.B1(n_2573),
.B2(n_2570),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_SL g4398 ( 
.A(n_4008),
.B(n_2577),
.Y(n_4398)
);

AOI22xp33_ASAP7_75t_L g4399 ( 
.A1(n_4117),
.A2(n_2339),
.B1(n_2342),
.B2(n_2338),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_4305),
.B(n_4308),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_4309),
.B(n_2578),
.Y(n_4401)
);

AOI22xp5_ASAP7_75t_L g4402 ( 
.A1(n_4072),
.A2(n_2581),
.B1(n_2583),
.B2(n_2580),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_4313),
.B(n_4316),
.Y(n_4403)
);

NOR2xp33_ASAP7_75t_L g4404 ( 
.A(n_4014),
.B(n_2586),
.Y(n_4404)
);

AND2x4_ASAP7_75t_L g4405 ( 
.A(n_4249),
.B(n_2360),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_SL g4406 ( 
.A(n_4071),
.B(n_2587),
.Y(n_4406)
);

INVx3_ASAP7_75t_L g4407 ( 
.A(n_4289),
.Y(n_4407)
);

INVx3_ASAP7_75t_L g4408 ( 
.A(n_4183),
.Y(n_4408)
);

NOR2xp33_ASAP7_75t_R g4409 ( 
.A(n_4064),
.B(n_2588),
.Y(n_4409)
);

HB1xp67_ASAP7_75t_L g4410 ( 
.A(n_4028),
.Y(n_4410)
);

NAND2x1p5_ASAP7_75t_L g4411 ( 
.A(n_4030),
.B(n_2362),
.Y(n_4411)
);

INVx2_ASAP7_75t_L g4412 ( 
.A(n_4039),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_4057),
.Y(n_4413)
);

BUFx3_ASAP7_75t_L g4414 ( 
.A(n_4184),
.Y(n_4414)
);

OAI22xp5_ASAP7_75t_SL g4415 ( 
.A1(n_4016),
.A2(n_2590),
.B1(n_2591),
.B2(n_2589),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_L g4416 ( 
.A(n_4322),
.B(n_2593),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_4325),
.B(n_2595),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_L g4418 ( 
.A(n_4327),
.B(n_2596),
.Y(n_4418)
);

AND2x4_ASAP7_75t_L g4419 ( 
.A(n_4257),
.B(n_2364),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_SL g4420 ( 
.A(n_4085),
.B(n_4363),
.Y(n_4420)
);

INVx5_ASAP7_75t_L g4421 ( 
.A(n_4116),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4043),
.Y(n_4422)
);

AND2x4_ASAP7_75t_SL g4423 ( 
.A(n_4053),
.B(n_2824),
.Y(n_4423)
);

BUFx2_ASAP7_75t_L g4424 ( 
.A(n_4221),
.Y(n_4424)
);

AOI22xp33_ASAP7_75t_L g4425 ( 
.A1(n_4042),
.A2(n_2369),
.B1(n_2373),
.B2(n_2367),
.Y(n_4425)
);

OR2x2_ASAP7_75t_L g4426 ( 
.A(n_4334),
.B(n_2600),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_4331),
.B(n_2601),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_SL g4428 ( 
.A(n_4061),
.B(n_2602),
.Y(n_4428)
);

AND2x4_ASAP7_75t_L g4429 ( 
.A(n_4276),
.B(n_2374),
.Y(n_4429)
);

BUFx6f_ASAP7_75t_L g4430 ( 
.A(n_4251),
.Y(n_4430)
);

NAND2x1p5_ASAP7_75t_L g4431 ( 
.A(n_4030),
.B(n_2375),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_4333),
.B(n_4335),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_4058),
.Y(n_4433)
);

INVx2_ASAP7_75t_L g4434 ( 
.A(n_4060),
.Y(n_4434)
);

INVx2_ASAP7_75t_SL g4435 ( 
.A(n_4192),
.Y(n_4435)
);

INVx2_ASAP7_75t_L g4436 ( 
.A(n_4070),
.Y(n_4436)
);

NAND2xp5_ASAP7_75t_L g4437 ( 
.A(n_4340),
.B(n_2603),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4343),
.B(n_2609),
.Y(n_4438)
);

BUFx2_ASAP7_75t_L g4439 ( 
.A(n_4199),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_4074),
.Y(n_4440)
);

NOR2x1p5_ASAP7_75t_L g4441 ( 
.A(n_4232),
.B(n_2614),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_4345),
.B(n_2615),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_4346),
.B(n_2624),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_4360),
.B(n_2625),
.Y(n_4444)
);

AND2x4_ASAP7_75t_L g4445 ( 
.A(n_4030),
.B(n_2383),
.Y(n_4445)
);

NOR2x1_ASAP7_75t_R g4446 ( 
.A(n_4150),
.B(n_2626),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4362),
.B(n_2628),
.Y(n_4447)
);

INVx6_ASAP7_75t_L g4448 ( 
.A(n_4108),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_4027),
.B(n_2629),
.Y(n_4449)
);

AOI21xp5_ASAP7_75t_L g4450 ( 
.A1(n_4189),
.A2(n_2387),
.B(n_2386),
.Y(n_4450)
);

BUFx12f_ASAP7_75t_L g4451 ( 
.A(n_4081),
.Y(n_4451)
);

OAI22xp5_ASAP7_75t_L g4452 ( 
.A1(n_4344),
.A2(n_4220),
.B1(n_4010),
.B2(n_4013),
.Y(n_4452)
);

INVx2_ASAP7_75t_SL g4453 ( 
.A(n_4277),
.Y(n_4453)
);

INVx4_ASAP7_75t_L g4454 ( 
.A(n_4150),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_L g4455 ( 
.A(n_4009),
.B(n_2632),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4047),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4048),
.Y(n_4457)
);

BUFx8_ASAP7_75t_L g4458 ( 
.A(n_4021),
.Y(n_4458)
);

AND2x6_ASAP7_75t_SL g4459 ( 
.A(n_4175),
.B(n_2393),
.Y(n_4459)
);

CKINVDCx8_ASAP7_75t_R g4460 ( 
.A(n_4118),
.Y(n_4460)
);

HB1xp67_ASAP7_75t_L g4461 ( 
.A(n_4218),
.Y(n_4461)
);

AND2x2_ASAP7_75t_SL g4462 ( 
.A(n_4069),
.B(n_2395),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_L g4463 ( 
.A(n_4012),
.B(n_4019),
.Y(n_4463)
);

OAI21xp33_ASAP7_75t_SL g4464 ( 
.A1(n_4086),
.A2(n_2411),
.B(n_2404),
.Y(n_4464)
);

BUFx8_ASAP7_75t_L g4465 ( 
.A(n_4173),
.Y(n_4465)
);

AOI22xp33_ASAP7_75t_L g4466 ( 
.A1(n_4153),
.A2(n_2423),
.B1(n_2428),
.B2(n_2416),
.Y(n_4466)
);

INVx2_ASAP7_75t_SL g4467 ( 
.A(n_4279),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4067),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_4075),
.Y(n_4469)
);

INVx2_ASAP7_75t_SL g4470 ( 
.A(n_4079),
.Y(n_4470)
);

NOR3xp33_ASAP7_75t_SL g4471 ( 
.A(n_4015),
.B(n_2634),
.C(n_2633),
.Y(n_4471)
);

INVx2_ASAP7_75t_L g4472 ( 
.A(n_4096),
.Y(n_4472)
);

INVxp33_ASAP7_75t_SL g4473 ( 
.A(n_4170),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_4022),
.B(n_4045),
.Y(n_4474)
);

AND2x6_ASAP7_75t_SL g4475 ( 
.A(n_4303),
.B(n_2430),
.Y(n_4475)
);

INVx2_ASAP7_75t_L g4476 ( 
.A(n_4098),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4080),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4083),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4034),
.B(n_2636),
.Y(n_4479)
);

INVx2_ASAP7_75t_L g4480 ( 
.A(n_4100),
.Y(n_4480)
);

CKINVDCx5p33_ASAP7_75t_R g4481 ( 
.A(n_4261),
.Y(n_4481)
);

BUFx2_ASAP7_75t_L g4482 ( 
.A(n_4195),
.Y(n_4482)
);

HB1xp67_ASAP7_75t_L g4483 ( 
.A(n_4233),
.Y(n_4483)
);

BUFx12f_ASAP7_75t_SL g4484 ( 
.A(n_4361),
.Y(n_4484)
);

NOR2xp33_ASAP7_75t_L g4485 ( 
.A(n_4066),
.B(n_2638),
.Y(n_4485)
);

AOI21xp33_ASAP7_75t_L g4486 ( 
.A1(n_4147),
.A2(n_2642),
.B(n_2639),
.Y(n_4486)
);

AOI22xp5_ASAP7_75t_L g4487 ( 
.A1(n_4202),
.A2(n_2647),
.B1(n_2648),
.B2(n_2645),
.Y(n_4487)
);

NOR2x1p5_ASAP7_75t_L g4488 ( 
.A(n_4300),
.B(n_2651),
.Y(n_4488)
);

AND2x4_ASAP7_75t_L g4489 ( 
.A(n_4150),
.B(n_2438),
.Y(n_4489)
);

AND2x6_ASAP7_75t_L g4490 ( 
.A(n_4157),
.B(n_2439),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4091),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4092),
.Y(n_4492)
);

BUFx6f_ASAP7_75t_SL g4493 ( 
.A(n_4040),
.Y(n_4493)
);

BUFx6f_ASAP7_75t_L g4494 ( 
.A(n_4099),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_4210),
.B(n_2652),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4106),
.Y(n_4496)
);

AND2x4_ASAP7_75t_L g4497 ( 
.A(n_4255),
.B(n_2447),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4095),
.Y(n_4498)
);

AOI22xp33_ASAP7_75t_L g4499 ( 
.A1(n_4358),
.A2(n_2456),
.B1(n_2462),
.B2(n_2450),
.Y(n_4499)
);

INVx2_ASAP7_75t_L g4500 ( 
.A(n_4115),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4049),
.B(n_2654),
.Y(n_4501)
);

OR2x2_ASAP7_75t_L g4502 ( 
.A(n_4065),
.B(n_2657),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4122),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4130),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_L g4505 ( 
.A(n_4051),
.B(n_2658),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_L g4506 ( 
.A(n_4151),
.B(n_2660),
.Y(n_4506)
);

INVx2_ASAP7_75t_L g4507 ( 
.A(n_4124),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_SL g4508 ( 
.A(n_4219),
.B(n_2661),
.Y(n_4508)
);

BUFx3_ASAP7_75t_L g4509 ( 
.A(n_4134),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_4125),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_4132),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_4311),
.B(n_2665),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_4359),
.B(n_4330),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4354),
.B(n_4138),
.Y(n_4514)
);

INVx6_ASAP7_75t_L g4515 ( 
.A(n_4246),
.Y(n_4515)
);

NOR2xp33_ASAP7_75t_L g4516 ( 
.A(n_4029),
.B(n_2667),
.Y(n_4516)
);

INVxp67_ASAP7_75t_SL g4517 ( 
.A(n_4140),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4145),
.Y(n_4518)
);

AND2x2_ASAP7_75t_L g4519 ( 
.A(n_4129),
.B(n_2824),
.Y(n_4519)
);

AOI22xp33_ASAP7_75t_SL g4520 ( 
.A1(n_4176),
.A2(n_2669),
.B1(n_2673),
.B2(n_2668),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4143),
.B(n_2674),
.Y(n_4521)
);

BUFx3_ASAP7_75t_L g4522 ( 
.A(n_4141),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_4320),
.B(n_2676),
.Y(n_4523)
);

INVx2_ASAP7_75t_L g4524 ( 
.A(n_4127),
.Y(n_4524)
);

O2A1O1Ixp33_ASAP7_75t_L g4525 ( 
.A1(n_4319),
.A2(n_2469),
.B(n_2472),
.C(n_2468),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4324),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_4336),
.B(n_4364),
.Y(n_4527)
);

INVx4_ASAP7_75t_L g4528 ( 
.A(n_4266),
.Y(n_4528)
);

AOI22xp33_ASAP7_75t_L g4529 ( 
.A1(n_4044),
.A2(n_4104),
.B1(n_4329),
.B2(n_4326),
.Y(n_4529)
);

NOR2x1p5_ASAP7_75t_L g4530 ( 
.A(n_4299),
.B(n_2678),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_4211),
.B(n_2679),
.Y(n_4531)
);

INVx2_ASAP7_75t_SL g4532 ( 
.A(n_4312),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_SL g4533 ( 
.A(n_4146),
.B(n_4250),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4165),
.Y(n_4534)
);

INVx2_ASAP7_75t_SL g4535 ( 
.A(n_4339),
.Y(n_4535)
);

HB1xp67_ASAP7_75t_L g4536 ( 
.A(n_4272),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4177),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_4212),
.B(n_2683),
.Y(n_4538)
);

INVxp33_ASAP7_75t_L g4539 ( 
.A(n_4196),
.Y(n_4539)
);

INVx1_ASAP7_75t_SL g4540 ( 
.A(n_4290),
.Y(n_4540)
);

NOR2xp67_ASAP7_75t_L g4541 ( 
.A(n_4304),
.B(n_1808),
.Y(n_4541)
);

BUFx2_ASAP7_75t_L g4542 ( 
.A(n_4298),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4186),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4203),
.Y(n_4544)
);

INVx2_ASAP7_75t_L g4545 ( 
.A(n_4144),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_SL g4546 ( 
.A(n_4250),
.B(n_2684),
.Y(n_4546)
);

NOR2xp33_ASAP7_75t_L g4547 ( 
.A(n_4056),
.B(n_2685),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_SL g4548 ( 
.A(n_4250),
.B(n_2687),
.Y(n_4548)
);

NAND2xp33_ASAP7_75t_SL g4549 ( 
.A(n_4103),
.B(n_2688),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_4214),
.B(n_2690),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_L g4551 ( 
.A(n_4215),
.B(n_2691),
.Y(n_4551)
);

BUFx12f_ASAP7_75t_L g4552 ( 
.A(n_4351),
.Y(n_4552)
);

AOI21xp5_ASAP7_75t_L g4553 ( 
.A1(n_4163),
.A2(n_2474),
.B(n_2473),
.Y(n_4553)
);

AND2x4_ASAP7_75t_L g4554 ( 
.A(n_4253),
.B(n_2478),
.Y(n_4554)
);

AOI22xp5_ASAP7_75t_L g4555 ( 
.A1(n_4190),
.A2(n_2693),
.B1(n_2694),
.B2(n_2692),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_SL g4556 ( 
.A(n_4323),
.B(n_2695),
.Y(n_4556)
);

INVx2_ASAP7_75t_L g4557 ( 
.A(n_4149),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_4154),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4206),
.Y(n_4559)
);

NAND2xp33_ASAP7_75t_L g4560 ( 
.A(n_4119),
.B(n_4162),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4341),
.B(n_4033),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_4110),
.B(n_2698),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_4306),
.Y(n_4563)
);

INVx2_ASAP7_75t_SL g4564 ( 
.A(n_4283),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4204),
.Y(n_4565)
);

AOI21xp5_ASAP7_75t_L g4566 ( 
.A1(n_4155),
.A2(n_2487),
.B(n_2482),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4168),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_4321),
.Y(n_4568)
);

CKINVDCx5p33_ASAP7_75t_R g4569 ( 
.A(n_4361),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4342),
.Y(n_4570)
);

AOI22xp33_ASAP7_75t_L g4571 ( 
.A1(n_4315),
.A2(n_2498),
.B1(n_2502),
.B2(n_2497),
.Y(n_4571)
);

AOI22xp33_ASAP7_75t_L g4572 ( 
.A1(n_4315),
.A2(n_2507),
.B1(n_2509),
.B2(n_2504),
.Y(n_4572)
);

BUFx2_ASAP7_75t_L g4573 ( 
.A(n_4315),
.Y(n_4573)
);

INVx2_ASAP7_75t_SL g4574 ( 
.A(n_4294),
.Y(n_4574)
);

INVx4_ASAP7_75t_L g4575 ( 
.A(n_4282),
.Y(n_4575)
);

NAND2xp5_ASAP7_75t_L g4576 ( 
.A(n_4180),
.B(n_4188),
.Y(n_4576)
);

NOR2xp33_ASAP7_75t_L g4577 ( 
.A(n_4142),
.B(n_2699),
.Y(n_4577)
);

NAND2xp5_ASAP7_75t_L g4578 ( 
.A(n_4097),
.B(n_2701),
.Y(n_4578)
);

BUFx6f_ASAP7_75t_L g4579 ( 
.A(n_4258),
.Y(n_4579)
);

NOR2x1p5_ASAP7_75t_L g4580 ( 
.A(n_4301),
.B(n_2704),
.Y(n_4580)
);

BUFx6f_ASAP7_75t_L g4581 ( 
.A(n_4280),
.Y(n_4581)
);

AOI22xp5_ASAP7_75t_L g4582 ( 
.A1(n_4174),
.A2(n_2707),
.B1(n_2710),
.B2(n_2706),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4347),
.Y(n_4583)
);

INVx2_ASAP7_75t_L g4584 ( 
.A(n_4356),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4357),
.B(n_2711),
.Y(n_4585)
);

HB1xp67_ASAP7_75t_L g4586 ( 
.A(n_4239),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_SL g4587 ( 
.A(n_4228),
.B(n_4169),
.Y(n_4587)
);

INVx1_ASAP7_75t_SL g4588 ( 
.A(n_4193),
.Y(n_4588)
);

NAND2xp5_ASAP7_75t_L g4589 ( 
.A(n_4152),
.B(n_4310),
.Y(n_4589)
);

BUFx8_ASAP7_75t_SL g4590 ( 
.A(n_4094),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4245),
.Y(n_4591)
);

INVx2_ASAP7_75t_SL g4592 ( 
.A(n_4278),
.Y(n_4592)
);

AOI22xp5_ASAP7_75t_L g4593 ( 
.A1(n_4123),
.A2(n_2713),
.B1(n_2714),
.B2(n_2712),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4207),
.Y(n_4594)
);

AND2x4_ASAP7_75t_L g4595 ( 
.A(n_4240),
.B(n_2519),
.Y(n_4595)
);

INVxp67_ASAP7_75t_SL g4596 ( 
.A(n_4119),
.Y(n_4596)
);

AND2x2_ASAP7_75t_L g4597 ( 
.A(n_4159),
.B(n_2715),
.Y(n_4597)
);

OR2x2_ASAP7_75t_SL g4598 ( 
.A(n_4236),
.B(n_2524),
.Y(n_4598)
);

INVx2_ASAP7_75t_L g4599 ( 
.A(n_4224),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_4229),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_L g4601 ( 
.A(n_4348),
.B(n_2716),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_SL g4602 ( 
.A(n_4248),
.B(n_2718),
.Y(n_4602)
);

NOR2xp33_ASAP7_75t_R g4603 ( 
.A(n_4338),
.B(n_2720),
.Y(n_4603)
);

A2O1A1Ixp33_ASAP7_75t_SL g4604 ( 
.A1(n_4172),
.A2(n_2529),
.B(n_2531),
.C(n_2527),
.Y(n_4604)
);

NOR2x1_ASAP7_75t_L g4605 ( 
.A(n_4068),
.B(n_2535),
.Y(n_4605)
);

NAND2xp33_ASAP7_75t_SL g4606 ( 
.A(n_4148),
.B(n_2723),
.Y(n_4606)
);

NOR2xp33_ASAP7_75t_L g4607 ( 
.A(n_4054),
.B(n_2729),
.Y(n_4607)
);

AOI22xp33_ASAP7_75t_L g4608 ( 
.A1(n_4337),
.A2(n_2540),
.B1(n_2543),
.B2(n_2538),
.Y(n_4608)
);

OR2x6_ASAP7_75t_L g4609 ( 
.A(n_4291),
.B(n_4243),
.Y(n_4609)
);

HB1xp67_ASAP7_75t_L g4610 ( 
.A(n_4225),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_4254),
.B(n_4077),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4252),
.Y(n_4612)
);

AND2x4_ASAP7_75t_L g4613 ( 
.A(n_4260),
.B(n_2544),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_4082),
.B(n_2730),
.Y(n_4614)
);

INVx5_ASAP7_75t_L g4615 ( 
.A(n_4296),
.Y(n_4615)
);

HB1xp67_ASAP7_75t_L g4616 ( 
.A(n_4267),
.Y(n_4616)
);

NOR2xp33_ASAP7_75t_L g4617 ( 
.A(n_4035),
.B(n_2731),
.Y(n_4617)
);

AOI22xp5_ASAP7_75t_L g4618 ( 
.A1(n_4213),
.A2(n_2739),
.B1(n_2740),
.B2(n_2735),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4167),
.Y(n_4619)
);

AOI21xp5_ASAP7_75t_L g4620 ( 
.A1(n_4160),
.A2(n_2551),
.B(n_2549),
.Y(n_4620)
);

AND2x4_ASAP7_75t_L g4621 ( 
.A(n_4293),
.B(n_2552),
.Y(n_4621)
);

BUFx6f_ASAP7_75t_L g4622 ( 
.A(n_4296),
.Y(n_4622)
);

BUFx2_ASAP7_75t_L g4623 ( 
.A(n_4296),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_SL g4624 ( 
.A(n_4208),
.B(n_2741),
.Y(n_4624)
);

HB1xp67_ASAP7_75t_L g4625 ( 
.A(n_4262),
.Y(n_4625)
);

INVx5_ASAP7_75t_L g4626 ( 
.A(n_4265),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4084),
.B(n_2746),
.Y(n_4627)
);

NOR2xp33_ASAP7_75t_L g4628 ( 
.A(n_4073),
.B(n_2750),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4164),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4088),
.B(n_2751),
.Y(n_4630)
);

INVx2_ASAP7_75t_L g4631 ( 
.A(n_4105),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4101),
.B(n_2752),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4166),
.Y(n_4633)
);

NAND2xp5_ASAP7_75t_SL g4634 ( 
.A(n_4235),
.B(n_4349),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4178),
.Y(n_4635)
);

AND2x4_ASAP7_75t_SL g4636 ( 
.A(n_4287),
.B(n_4264),
.Y(n_4636)
);

HB1xp67_ASAP7_75t_L g4637 ( 
.A(n_4263),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4102),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4109),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_4111),
.B(n_2754),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4119),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_L g4642 ( 
.A(n_4121),
.B(n_2756),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4023),
.B(n_2758),
.Y(n_4643)
);

HB1xp67_ASAP7_75t_L g4644 ( 
.A(n_4268),
.Y(n_4644)
);

AOI22xp33_ASAP7_75t_L g4645 ( 
.A1(n_4026),
.A2(n_2582),
.B1(n_2584),
.B2(n_2576),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4126),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_L g4647 ( 
.A(n_4128),
.B(n_2762),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_SL g4648 ( 
.A(n_4131),
.B(n_2763),
.Y(n_4648)
);

BUFx6f_ASAP7_75t_L g4649 ( 
.A(n_4238),
.Y(n_4649)
);

INVx4_ASAP7_75t_L g4650 ( 
.A(n_4137),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4133),
.B(n_2767),
.Y(n_4651)
);

AND2x4_ASAP7_75t_L g4652 ( 
.A(n_4242),
.B(n_2585),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4135),
.Y(n_4653)
);

INVxp67_ASAP7_75t_L g4654 ( 
.A(n_4275),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4119),
.Y(n_4655)
);

AND3x1_ASAP7_75t_L g4656 ( 
.A(n_4017),
.B(n_2599),
.C(n_2598),
.Y(n_4656)
);

NOR2xp33_ASAP7_75t_L g4657 ( 
.A(n_4062),
.B(n_2768),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4181),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_SL g4659 ( 
.A(n_4513),
.B(n_4050),
.Y(n_4659)
);

NAND2xp5_ASAP7_75t_SL g4660 ( 
.A(n_4654),
.B(n_4055),
.Y(n_4660)
);

NAND2xp33_ASAP7_75t_SL g4661 ( 
.A(n_4454),
.B(n_4089),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_SL g4662 ( 
.A(n_4514),
.B(n_4611),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4474),
.B(n_4314),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_SL g4664 ( 
.A(n_4588),
.B(n_4269),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_SL g4665 ( 
.A(n_4400),
.B(n_4273),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_SL g4666 ( 
.A(n_4403),
.B(n_4332),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_SL g4667 ( 
.A(n_4432),
.B(n_4271),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_SL g4668 ( 
.A(n_4540),
.B(n_4274),
.Y(n_4668)
);

NAND2xp5_ASAP7_75t_SL g4669 ( 
.A(n_4463),
.B(n_4237),
.Y(n_4669)
);

NAND2xp33_ASAP7_75t_SL g4670 ( 
.A(n_4622),
.B(n_4230),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4638),
.B(n_4317),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4639),
.B(n_4646),
.Y(n_4672)
);

NAND2xp5_ASAP7_75t_SL g4673 ( 
.A(n_4371),
.B(n_4328),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_SL g4674 ( 
.A(n_4539),
.B(n_4353),
.Y(n_4674)
);

NAND2xp5_ASAP7_75t_SL g4675 ( 
.A(n_4587),
.B(n_4185),
.Y(n_4675)
);

NAND2xp33_ASAP7_75t_SL g4676 ( 
.A(n_4622),
.B(n_4259),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_SL g4677 ( 
.A(n_4653),
.B(n_4191),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_SL g4678 ( 
.A(n_4658),
.B(n_4200),
.Y(n_4678)
);

NAND2xp5_ASAP7_75t_SL g4679 ( 
.A(n_4615),
.B(n_4201),
.Y(n_4679)
);

NAND2xp5_ASAP7_75t_SL g4680 ( 
.A(n_4615),
.B(n_4281),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_4374),
.B(n_4352),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_SL g4682 ( 
.A(n_4629),
.B(n_4633),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_SL g4683 ( 
.A(n_4635),
.B(n_4285),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4365),
.B(n_4223),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_SL g4685 ( 
.A(n_4577),
.B(n_4286),
.Y(n_4685)
);

NAND2xp33_ASAP7_75t_SL g4686 ( 
.A(n_4471),
.B(n_4241),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_SL g4687 ( 
.A(n_4562),
.B(n_4288),
.Y(n_4687)
);

NAND2xp33_ASAP7_75t_SL g4688 ( 
.A(n_4573),
.B(n_4256),
.Y(n_4688)
);

NAND2xp33_ASAP7_75t_SL g4689 ( 
.A(n_4634),
.B(n_4623),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_SL g4690 ( 
.A(n_4430),
.B(n_4295),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_SL g4691 ( 
.A(n_4430),
.B(n_4234),
.Y(n_4691)
);

NAND2xp33_ASAP7_75t_SL g4692 ( 
.A(n_4376),
.B(n_4227),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4495),
.B(n_4226),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_SL g4694 ( 
.A(n_4561),
.B(n_4292),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_SL g4695 ( 
.A(n_4578),
.B(n_4302),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_SL g4696 ( 
.A(n_4404),
.B(n_4217),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_SL g4697 ( 
.A(n_4519),
.B(n_4161),
.Y(n_4697)
);

NAND2xp33_ASAP7_75t_SL g4698 ( 
.A(n_4376),
.B(n_4216),
.Y(n_4698)
);

NAND2xp33_ASAP7_75t_SL g4699 ( 
.A(n_4391),
.B(n_4171),
.Y(n_4699)
);

NAND2xp33_ASAP7_75t_L g4700 ( 
.A(n_4529),
.B(n_4179),
.Y(n_4700)
);

NAND2xp33_ASAP7_75t_SL g4701 ( 
.A(n_4391),
.B(n_4139),
.Y(n_4701)
);

AND2x4_ASAP7_75t_L g4702 ( 
.A(n_4609),
.B(n_4297),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_SL g4703 ( 
.A(n_4393),
.B(n_4197),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_SL g4704 ( 
.A(n_4386),
.B(n_4136),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_SL g4705 ( 
.A(n_4597),
.B(n_4156),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_SL g4706 ( 
.A(n_4547),
.B(n_4112),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_SL g4707 ( 
.A(n_4410),
.B(n_4120),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_SL g4708 ( 
.A(n_4370),
.B(n_4244),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4516),
.B(n_4076),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_SL g4710 ( 
.A(n_4649),
.B(n_4284),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4387),
.B(n_4182),
.Y(n_4711)
);

NAND2xp33_ASAP7_75t_SL g4712 ( 
.A(n_4603),
.B(n_4270),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_SL g4713 ( 
.A(n_4649),
.B(n_4222),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4643),
.B(n_4137),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4449),
.B(n_4187),
.Y(n_4715)
);

NAND2xp5_ASAP7_75t_SL g4716 ( 
.A(n_4581),
.B(n_4198),
.Y(n_4716)
);

NAND2xp33_ASAP7_75t_SL g4717 ( 
.A(n_4530),
.B(n_4194),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_SL g4718 ( 
.A(n_4581),
.B(n_4114),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4455),
.B(n_4350),
.Y(n_4719)
);

NAND2xp5_ASAP7_75t_SL g4720 ( 
.A(n_4626),
.B(n_4209),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_SL g4721 ( 
.A(n_4626),
.B(n_4052),
.Y(n_4721)
);

NAND2xp33_ASAP7_75t_SL g4722 ( 
.A(n_4580),
.B(n_2769),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_SL g4723 ( 
.A(n_4625),
.B(n_2770),
.Y(n_4723)
);

NAND2xp5_ASAP7_75t_SL g4724 ( 
.A(n_4637),
.B(n_2772),
.Y(n_4724)
);

AND2x2_ASAP7_75t_L g4725 ( 
.A(n_4462),
.B(n_2773),
.Y(n_4725)
);

NAND2xp5_ASAP7_75t_SL g4726 ( 
.A(n_4644),
.B(n_2775),
.Y(n_4726)
);

NAND2xp33_ASAP7_75t_SL g4727 ( 
.A(n_4494),
.B(n_2784),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4401),
.B(n_4231),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_SL g4729 ( 
.A(n_4657),
.B(n_2786),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_SL g4730 ( 
.A(n_4579),
.B(n_2787),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4416),
.B(n_2606),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_SL g4732 ( 
.A(n_4579),
.B(n_2788),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4485),
.B(n_2790),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_L g4734 ( 
.A(n_4417),
.B(n_2607),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_SL g4735 ( 
.A(n_4375),
.B(n_2791),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_L g4736 ( 
.A(n_4418),
.B(n_2612),
.Y(n_4736)
);

NAND2xp33_ASAP7_75t_SL g4737 ( 
.A(n_4494),
.B(n_2793),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_SL g4738 ( 
.A(n_4435),
.B(n_4512),
.Y(n_4738)
);

NAND2xp5_ASAP7_75t_SL g4739 ( 
.A(n_4527),
.B(n_2799),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4427),
.B(n_2613),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_SL g4741 ( 
.A(n_4439),
.B(n_2800),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_SL g4742 ( 
.A(n_4586),
.B(n_2803),
.Y(n_4742)
);

NAND2xp5_ASAP7_75t_L g4743 ( 
.A(n_4437),
.B(n_2616),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4628),
.B(n_2804),
.Y(n_4744)
);

AND2x2_ASAP7_75t_L g4745 ( 
.A(n_4613),
.B(n_2805),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4650),
.B(n_2808),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4438),
.B(n_2618),
.Y(n_4747)
);

NAND2xp33_ASAP7_75t_SL g4748 ( 
.A(n_4384),
.B(n_4542),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_SL g4749 ( 
.A(n_4517),
.B(n_2809),
.Y(n_4749)
);

OR2x2_ASAP7_75t_L g4750 ( 
.A(n_4426),
.B(n_2814),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4442),
.B(n_2619),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_SL g4752 ( 
.A(n_4497),
.B(n_2815),
.Y(n_4752)
);

NAND2xp5_ASAP7_75t_SL g4753 ( 
.A(n_4607),
.B(n_2816),
.Y(n_4753)
);

NAND2xp33_ASAP7_75t_SL g4754 ( 
.A(n_4372),
.B(n_2826),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_SL g4755 ( 
.A(n_4452),
.B(n_2827),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_4443),
.B(n_2620),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_SL g4757 ( 
.A(n_4616),
.B(n_2828),
.Y(n_4757)
);

OR2x2_ASAP7_75t_L g4758 ( 
.A(n_4502),
.B(n_2832),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_SL g4759 ( 
.A(n_4531),
.B(n_2834),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_SL g4760 ( 
.A(n_4538),
.B(n_2835),
.Y(n_4760)
);

NAND2xp33_ASAP7_75t_SL g4761 ( 
.A(n_4379),
.B(n_2837),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_SL g4762 ( 
.A(n_4550),
.B(n_2838),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_SL g4763 ( 
.A(n_4551),
.B(n_4479),
.Y(n_4763)
);

NAND2xp5_ASAP7_75t_SL g4764 ( 
.A(n_4501),
.B(n_2839),
.Y(n_4764)
);

NAND2xp33_ASAP7_75t_SL g4765 ( 
.A(n_4392),
.B(n_2844),
.Y(n_4765)
);

NAND2xp33_ASAP7_75t_SL g4766 ( 
.A(n_4422),
.B(n_2846),
.Y(n_4766)
);

NAND2xp33_ASAP7_75t_SL g4767 ( 
.A(n_4456),
.B(n_2847),
.Y(n_4767)
);

NAND2xp33_ASAP7_75t_SL g4768 ( 
.A(n_4457),
.B(n_2848),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_SL g4769 ( 
.A(n_4505),
.B(n_2850),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_SL g4770 ( 
.A(n_4444),
.B(n_2851),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_SL g4771 ( 
.A(n_4447),
.B(n_2853),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_SL g4772 ( 
.A(n_4610),
.B(n_2854),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4506),
.B(n_2622),
.Y(n_4773)
);

NAND2xp5_ASAP7_75t_L g4774 ( 
.A(n_4521),
.B(n_4614),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4627),
.B(n_2623),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_SL g4776 ( 
.A(n_4565),
.B(n_2857),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_SL g4777 ( 
.A(n_4617),
.B(n_2861),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_SL g4778 ( 
.A(n_4424),
.B(n_2863),
.Y(n_4778)
);

NAND2xp5_ASAP7_75t_SL g4779 ( 
.A(n_4630),
.B(n_2865),
.Y(n_4779)
);

NAND2xp33_ASAP7_75t_SL g4780 ( 
.A(n_4468),
.B(n_2866),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_SL g4781 ( 
.A(n_4632),
.B(n_2867),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_SL g4782 ( 
.A(n_4640),
.B(n_2868),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_SL g4783 ( 
.A(n_4642),
.B(n_2875),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4647),
.B(n_2631),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_SL g4785 ( 
.A(n_4651),
.B(n_2877),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4469),
.B(n_2643),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_SL g4787 ( 
.A(n_4567),
.B(n_2883),
.Y(n_4787)
);

XNOR2xp5_ASAP7_75t_SL g4788 ( 
.A(n_4481),
.B(n_4569),
.Y(n_4788)
);

AND2x2_ASAP7_75t_L g4789 ( 
.A(n_4429),
.B(n_2885),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_SL g4790 ( 
.A(n_4482),
.B(n_2890),
.Y(n_4790)
);

NAND2xp33_ASAP7_75t_SL g4791 ( 
.A(n_4477),
.B(n_2893),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_SL g4792 ( 
.A(n_4420),
.B(n_2894),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_SL g4793 ( 
.A(n_4396),
.B(n_2896),
.Y(n_4793)
);

NAND2xp33_ASAP7_75t_SL g4794 ( 
.A(n_4478),
.B(n_2898),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_SL g4795 ( 
.A(n_4394),
.B(n_2899),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_SL g4796 ( 
.A(n_4407),
.B(n_2901),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_SL g4797 ( 
.A(n_4491),
.B(n_2903),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_SL g4798 ( 
.A(n_4492),
.B(n_2908),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_SL g4799 ( 
.A(n_4498),
.B(n_2911),
.Y(n_4799)
);

NAND2xp33_ASAP7_75t_SL g4800 ( 
.A(n_4503),
.B(n_2912),
.Y(n_4800)
);

NAND2xp33_ASAP7_75t_SL g4801 ( 
.A(n_4504),
.B(n_2913),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_SL g4802 ( 
.A(n_4511),
.B(n_2914),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4518),
.B(n_2650),
.Y(n_4803)
);

OR2x2_ASAP7_75t_L g4804 ( 
.A(n_4523),
.B(n_2915),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_SL g4805 ( 
.A(n_4526),
.B(n_2918),
.Y(n_4805)
);

NAND2xp33_ASAP7_75t_SL g4806 ( 
.A(n_4534),
.B(n_2924),
.Y(n_4806)
);

NAND2xp5_ASAP7_75t_L g4807 ( 
.A(n_4537),
.B(n_2653),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_SL g4808 ( 
.A(n_4543),
.B(n_2925),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4544),
.B(n_2656),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_L g4810 ( 
.A(n_4559),
.B(n_2670),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_SL g4811 ( 
.A(n_4619),
.B(n_2926),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_SL g4812 ( 
.A(n_4589),
.B(n_2927),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_SL g4813 ( 
.A(n_4382),
.B(n_2930),
.Y(n_4813)
);

NAND2xp5_ASAP7_75t_SL g4814 ( 
.A(n_4382),
.B(n_2931),
.Y(n_4814)
);

AND2x4_ASAP7_75t_L g4815 ( 
.A(n_4609),
.B(n_2677),
.Y(n_4815)
);

NAND2xp33_ASAP7_75t_SL g4816 ( 
.A(n_4528),
.B(n_2933),
.Y(n_4816)
);

NAND2xp5_ASAP7_75t_SL g4817 ( 
.A(n_4636),
.B(n_2935),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_SL g4818 ( 
.A(n_4564),
.B(n_2938),
.Y(n_4818)
);

NAND2xp5_ASAP7_75t_SL g4819 ( 
.A(n_4574),
.B(n_2939),
.Y(n_4819)
);

NAND2xp5_ASAP7_75t_SL g4820 ( 
.A(n_4591),
.B(n_2942),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_SL g4821 ( 
.A(n_4599),
.B(n_2943),
.Y(n_4821)
);

AND2x4_ASAP7_75t_L g4822 ( 
.A(n_4414),
.B(n_2681),
.Y(n_4822)
);

NAND2xp33_ASAP7_75t_SL g4823 ( 
.A(n_4592),
.B(n_2944),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_SL g4824 ( 
.A(n_4600),
.B(n_2947),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_SL g4825 ( 
.A(n_4486),
.B(n_2948),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_SL g4826 ( 
.A(n_4536),
.B(n_2949),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4366),
.B(n_4377),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_L g4828 ( 
.A(n_4377),
.B(n_2697),
.Y(n_4828)
);

NAND2xp5_ASAP7_75t_SL g4829 ( 
.A(n_4520),
.B(n_2950),
.Y(n_4829)
);

NAND2xp5_ASAP7_75t_SL g4830 ( 
.A(n_4367),
.B(n_2951),
.Y(n_4830)
);

NAND2xp33_ASAP7_75t_SL g4831 ( 
.A(n_4408),
.B(n_2952),
.Y(n_4831)
);

NAND2xp5_ASAP7_75t_SL g4832 ( 
.A(n_4380),
.B(n_2955),
.Y(n_4832)
);

NAND2xp33_ASAP7_75t_SL g4833 ( 
.A(n_4533),
.B(n_2956),
.Y(n_4833)
);

NAND2xp33_ASAP7_75t_SL g4834 ( 
.A(n_4575),
.B(n_2957),
.Y(n_4834)
);

NAND2xp33_ASAP7_75t_SL g4835 ( 
.A(n_4532),
.B(n_2959),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_SL g4836 ( 
.A(n_4389),
.B(n_4395),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_SL g4837 ( 
.A(n_4412),
.B(n_2960),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_SL g4838 ( 
.A(n_4413),
.B(n_2961),
.Y(n_4838)
);

NAND2xp33_ASAP7_75t_SL g4839 ( 
.A(n_4535),
.B(n_2962),
.Y(n_4839)
);

AND2x4_ASAP7_75t_L g4840 ( 
.A(n_4368),
.B(n_2700),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_SL g4841 ( 
.A(n_4433),
.B(n_2964),
.Y(n_4841)
);

NAND2xp5_ASAP7_75t_SL g4842 ( 
.A(n_4434),
.B(n_2965),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4377),
.B(n_2705),
.Y(n_4843)
);

NAND2xp5_ASAP7_75t_SL g4844 ( 
.A(n_4436),
.B(n_4440),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_SL g4845 ( 
.A(n_4472),
.B(n_2966),
.Y(n_4845)
);

NAND2xp5_ASAP7_75t_SL g4846 ( 
.A(n_4476),
.B(n_2968),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_SL g4847 ( 
.A(n_4480),
.B(n_2970),
.Y(n_4847)
);

NAND2xp5_ASAP7_75t_SL g4848 ( 
.A(n_4496),
.B(n_2976),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_SL g4849 ( 
.A(n_4500),
.B(n_2978),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_SL g4850 ( 
.A(n_4507),
.B(n_2980),
.Y(n_4850)
);

NOR2xp33_ASAP7_75t_L g4851 ( 
.A(n_4515),
.B(n_2981),
.Y(n_4851)
);

NAND2xp5_ASAP7_75t_SL g4852 ( 
.A(n_4510),
.B(n_2982),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_SL g4853 ( 
.A(n_4524),
.B(n_2984),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_SL g4854 ( 
.A(n_4545),
.B(n_2985),
.Y(n_4854)
);

NAND2xp5_ASAP7_75t_L g4855 ( 
.A(n_4373),
.B(n_2721),
.Y(n_4855)
);

NAND2xp33_ASAP7_75t_SL g4856 ( 
.A(n_4470),
.B(n_2987),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4490),
.B(n_2725),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_L g4858 ( 
.A(n_4490),
.B(n_2728),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_SL g4859 ( 
.A(n_4557),
.B(n_2988),
.Y(n_4859)
);

NAND2xp33_ASAP7_75t_SL g4860 ( 
.A(n_4453),
.B(n_2990),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_SL g4861 ( 
.A(n_4558),
.B(n_2993),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_SL g4862 ( 
.A(n_4563),
.B(n_2994),
.Y(n_4862)
);

NAND2xp5_ASAP7_75t_L g4863 ( 
.A(n_4490),
.B(n_2732),
.Y(n_4863)
);

NAND2xp5_ASAP7_75t_SL g4864 ( 
.A(n_4568),
.B(n_2995),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_SL g4865 ( 
.A(n_4584),
.B(n_2998),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_SL g4866 ( 
.A(n_4399),
.B(n_2733),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_SL g4867 ( 
.A(n_4593),
.B(n_4656),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_SL g4868 ( 
.A(n_4570),
.B(n_2737),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_SL g4869 ( 
.A(n_4583),
.B(n_2738),
.Y(n_4869)
);

NAND2x1p5_ASAP7_75t_L g4870 ( 
.A(n_4641),
.B(n_2743),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_SL g4871 ( 
.A(n_4594),
.B(n_2744),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_SL g4872 ( 
.A(n_4378),
.B(n_2745),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_4585),
.B(n_2747),
.Y(n_4873)
);

NAND2xp33_ASAP7_75t_SL g4874 ( 
.A(n_4467),
.B(n_2753),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_SL g4875 ( 
.A(n_4576),
.B(n_2757),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_SL g4876 ( 
.A(n_4411),
.B(n_2759),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_SL g4877 ( 
.A(n_4431),
.B(n_2765),
.Y(n_4877)
);

NAND2xp33_ASAP7_75t_SL g4878 ( 
.A(n_4546),
.B(n_2766),
.Y(n_4878)
);

AND2x4_ASAP7_75t_L g4879 ( 
.A(n_4369),
.B(n_4383),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_SL g4880 ( 
.A(n_4409),
.B(n_2777),
.Y(n_4880)
);

NAND2x1p5_ASAP7_75t_L g4881 ( 
.A(n_4655),
.B(n_2778),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_L g4882 ( 
.A(n_4566),
.B(n_2779),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_SL g4883 ( 
.A(n_4473),
.B(n_2781),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_SL g4884 ( 
.A(n_4388),
.B(n_2782),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_SL g4885 ( 
.A(n_4428),
.B(n_2795),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_SL g4886 ( 
.A(n_4555),
.B(n_2797),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_SL g4887 ( 
.A(n_4487),
.B(n_2798),
.Y(n_4887)
);

AND2x2_ASAP7_75t_L g4888 ( 
.A(n_4595),
.B(n_2801),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_SL g4889 ( 
.A(n_4612),
.B(n_2806),
.Y(n_4889)
);

NAND2xp33_ASAP7_75t_SL g4890 ( 
.A(n_4548),
.B(n_2810),
.Y(n_4890)
);

NAND2xp5_ASAP7_75t_SL g4891 ( 
.A(n_4461),
.B(n_2813),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_SL g4892 ( 
.A(n_4483),
.B(n_2817),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_SL g4893 ( 
.A(n_4385),
.B(n_2822),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_SL g4894 ( 
.A(n_4405),
.B(n_2823),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_SL g4895 ( 
.A(n_4419),
.B(n_2825),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_SL g4896 ( 
.A(n_4445),
.B(n_2829),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_SL g4897 ( 
.A(n_4489),
.B(n_2831),
.Y(n_4897)
);

NAND2xp5_ASAP7_75t_SL g4898 ( 
.A(n_4652),
.B(n_2833),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_SL g4899 ( 
.A(n_4582),
.B(n_4648),
.Y(n_4899)
);

NAND2xp5_ASAP7_75t_SL g4900 ( 
.A(n_4549),
.B(n_2836),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_SL g4901 ( 
.A(n_4402),
.B(n_2840),
.Y(n_4901)
);

NAND2xp5_ASAP7_75t_SL g4902 ( 
.A(n_4618),
.B(n_2843),
.Y(n_4902)
);

NAND2xp5_ASAP7_75t_SL g4903 ( 
.A(n_4571),
.B(n_2856),
.Y(n_4903)
);

NAND2xp5_ASAP7_75t_SL g4904 ( 
.A(n_4572),
.B(n_2858),
.Y(n_4904)
);

NAND2xp5_ASAP7_75t_SL g4905 ( 
.A(n_4554),
.B(n_2859),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_SL g4906 ( 
.A(n_4606),
.B(n_2860),
.Y(n_4906)
);

AND2x2_ASAP7_75t_SL g4907 ( 
.A(n_4381),
.B(n_4560),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_SL g4908 ( 
.A(n_4601),
.B(n_2864),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_SL g4909 ( 
.A(n_4621),
.B(n_2869),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4425),
.B(n_2871),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_SL g4911 ( 
.A(n_4398),
.B(n_2873),
.Y(n_4911)
);

NAND2xp33_ASAP7_75t_SL g4912 ( 
.A(n_4493),
.B(n_2879),
.Y(n_4912)
);

NAND2xp5_ASAP7_75t_SL g4913 ( 
.A(n_4406),
.B(n_2882),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_SL g4914 ( 
.A(n_4415),
.B(n_2884),
.Y(n_4914)
);

NAND2xp5_ASAP7_75t_SL g4915 ( 
.A(n_4509),
.B(n_2889),
.Y(n_4915)
);

NAND2xp5_ASAP7_75t_SL g4916 ( 
.A(n_4522),
.B(n_2897),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_SL g4917 ( 
.A(n_4423),
.B(n_2900),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_SL g4918 ( 
.A(n_4508),
.B(n_2906),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_SL g4919 ( 
.A(n_4602),
.B(n_2909),
.Y(n_4919)
);

NAND2xp33_ASAP7_75t_SL g4920 ( 
.A(n_4488),
.B(n_2910),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_SL g4921 ( 
.A(n_4421),
.B(n_2920),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_SL g4922 ( 
.A(n_4421),
.B(n_2921),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_SL g4923 ( 
.A(n_4624),
.B(n_2922),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4390),
.B(n_2928),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_SL g4925 ( 
.A(n_4541),
.B(n_2941),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_SL g4926 ( 
.A(n_4556),
.B(n_2954),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_SL g4927 ( 
.A(n_4466),
.B(n_2958),
.Y(n_4927)
);

NAND2xp33_ASAP7_75t_SL g4928 ( 
.A(n_4441),
.B(n_2969),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4397),
.B(n_2973),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_L g4930 ( 
.A(n_4450),
.B(n_2975),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4620),
.B(n_2977),
.Y(n_4931)
);

NAND2xp5_ASAP7_75t_SL g4932 ( 
.A(n_4605),
.B(n_4460),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_SL g4933 ( 
.A(n_4608),
.B(n_4465),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_SL g4934 ( 
.A(n_4552),
.B(n_4553),
.Y(n_4934)
);

NAND2xp33_ASAP7_75t_SL g4935 ( 
.A(n_4499),
.B(n_2),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4464),
.B(n_2),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_SL g4937 ( 
.A(n_4525),
.B(n_3),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_SL g4938 ( 
.A(n_4596),
.B(n_3),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_SL g4939 ( 
.A(n_4645),
.B(n_5),
.Y(n_4939)
);

AND2x2_ASAP7_75t_L g4940 ( 
.A(n_4448),
.B(n_5),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_SL g4941 ( 
.A(n_4631),
.B(n_6),
.Y(n_4941)
);

NAND2xp5_ASAP7_75t_SL g4942 ( 
.A(n_4458),
.B(n_6),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_SL g4943 ( 
.A(n_4451),
.B(n_7),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_SL g4944 ( 
.A(n_4598),
.B(n_8),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_SL g4945 ( 
.A(n_4459),
.B(n_8),
.Y(n_4945)
);

NAND2xp5_ASAP7_75t_SL g4946 ( 
.A(n_4484),
.B(n_4590),
.Y(n_4946)
);

NAND2xp33_ASAP7_75t_SL g4947 ( 
.A(n_4446),
.B(n_9),
.Y(n_4947)
);

NAND2xp5_ASAP7_75t_SL g4948 ( 
.A(n_4475),
.B(n_9),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_SL g4949 ( 
.A(n_4604),
.B(n_10),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_SL g4950 ( 
.A(n_4513),
.B(n_11),
.Y(n_4950)
);

NAND2xp33_ASAP7_75t_SL g4951 ( 
.A(n_4454),
.B(n_11),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_SL g4952 ( 
.A(n_4513),
.B(n_12),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_SL g4953 ( 
.A(n_4513),
.B(n_12),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_SL g4954 ( 
.A(n_4513),
.B(n_13),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_SL g4955 ( 
.A(n_4513),
.B(n_13),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_SL g4956 ( 
.A(n_4513),
.B(n_15),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_SL g4957 ( 
.A(n_4513),
.B(n_16),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_L g4958 ( 
.A(n_4514),
.B(n_16),
.Y(n_4958)
);

INVxp67_ASAP7_75t_L g4959 ( 
.A(n_4851),
.Y(n_4959)
);

INVx2_ASAP7_75t_L g4960 ( 
.A(n_4836),
.Y(n_4960)
);

INVx3_ASAP7_75t_L g4961 ( 
.A(n_4879),
.Y(n_4961)
);

AOI22xp33_ASAP7_75t_L g4962 ( 
.A1(n_4700),
.A2(n_20),
.B1(n_17),
.B2(n_18),
.Y(n_4962)
);

INVx2_ASAP7_75t_L g4963 ( 
.A(n_4844),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4672),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4682),
.Y(n_4965)
);

AND2x2_ASAP7_75t_L g4966 ( 
.A(n_4714),
.B(n_17),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4786),
.Y(n_4967)
);

AND2x2_ASAP7_75t_L g4968 ( 
.A(n_4725),
.B(n_18),
.Y(n_4968)
);

AND3x1_ASAP7_75t_SL g4969 ( 
.A(n_4945),
.B(n_4942),
.C(n_4948),
.Y(n_4969)
);

AND2x2_ASAP7_75t_L g4970 ( 
.A(n_4744),
.B(n_20),
.Y(n_4970)
);

BUFx2_ASAP7_75t_L g4971 ( 
.A(n_4748),
.Y(n_4971)
);

CKINVDCx5p33_ASAP7_75t_R g4972 ( 
.A(n_4879),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_4662),
.B(n_21),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4870),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4803),
.Y(n_4975)
);

OAI22xp5_ASAP7_75t_SL g4976 ( 
.A1(n_4663),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4774),
.B(n_23),
.Y(n_4977)
);

INVx1_ASAP7_75t_L g4978 ( 
.A(n_4807),
.Y(n_4978)
);

NOR2xp33_ASAP7_75t_L g4979 ( 
.A(n_4665),
.B(n_1809),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4809),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4810),
.Y(n_4981)
);

NOR2xp67_ASAP7_75t_L g4982 ( 
.A(n_4873),
.B(n_1810),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_4693),
.B(n_25),
.Y(n_4983)
);

NAND2xp33_ASAP7_75t_L g4984 ( 
.A(n_4709),
.B(n_26),
.Y(n_4984)
);

BUFx3_ASAP7_75t_L g4985 ( 
.A(n_4822),
.Y(n_4985)
);

AND2x2_ASAP7_75t_L g4986 ( 
.A(n_4733),
.B(n_26),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4882),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4684),
.B(n_27),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4931),
.Y(n_4989)
);

A2O1A1Ixp33_ASAP7_75t_SL g4990 ( 
.A1(n_4936),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_4990)
);

AND2x4_ASAP7_75t_L g4991 ( 
.A(n_4702),
.B(n_4815),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4958),
.Y(n_4992)
);

AND2x4_ASAP7_75t_L g4993 ( 
.A(n_4702),
.B(n_4815),
.Y(n_4993)
);

BUFx6f_ASAP7_75t_L g4994 ( 
.A(n_4822),
.Y(n_4994)
);

INVx2_ASAP7_75t_L g4995 ( 
.A(n_4870),
.Y(n_4995)
);

INVx2_ASAP7_75t_L g4996 ( 
.A(n_4881),
.Y(n_4996)
);

CKINVDCx5p33_ASAP7_75t_R g4997 ( 
.A(n_4946),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4930),
.Y(n_4998)
);

AOI22xp33_ASAP7_75t_L g4999 ( 
.A1(n_4867),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_4999)
);

BUFx3_ASAP7_75t_L g5000 ( 
.A(n_4840),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_SL g5001 ( 
.A(n_4671),
.B(n_33),
.Y(n_5001)
);

HB1xp67_ASAP7_75t_L g5002 ( 
.A(n_4738),
.Y(n_5002)
);

AND2x2_ASAP7_75t_L g5003 ( 
.A(n_4888),
.B(n_4746),
.Y(n_5003)
);

NAND2x1p5_ASAP7_75t_L g5004 ( 
.A(n_4690),
.B(n_1814),
.Y(n_5004)
);

AND2x2_ASAP7_75t_L g5005 ( 
.A(n_4745),
.B(n_33),
.Y(n_5005)
);

AND2x2_ASAP7_75t_L g5006 ( 
.A(n_4713),
.B(n_34),
.Y(n_5006)
);

AND3x1_ASAP7_75t_SL g5007 ( 
.A(n_4944),
.B(n_35),
.C(n_36),
.Y(n_5007)
);

INVx3_ASAP7_75t_L g5008 ( 
.A(n_4840),
.Y(n_5008)
);

OR2x2_ASAP7_75t_L g5009 ( 
.A(n_4659),
.B(n_36),
.Y(n_5009)
);

AND2x2_ASAP7_75t_L g5010 ( 
.A(n_4940),
.B(n_37),
.Y(n_5010)
);

AOI22xp33_ASAP7_75t_L g5011 ( 
.A1(n_4935),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4677),
.Y(n_5012)
);

AO22x1_ASAP7_75t_L g5013 ( 
.A1(n_4827),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_5013)
);

CKINVDCx5p33_ASAP7_75t_R g5014 ( 
.A(n_4727),
.Y(n_5014)
);

AOI22xp5_ASAP7_75t_L g5015 ( 
.A1(n_4817),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4678),
.Y(n_5016)
);

INVx3_ASAP7_75t_L g5017 ( 
.A(n_4881),
.Y(n_5017)
);

BUFx2_ASAP7_75t_L g5018 ( 
.A(n_4692),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4924),
.Y(n_5019)
);

BUFx8_ASAP7_75t_L g5020 ( 
.A(n_4789),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4763),
.B(n_42),
.Y(n_5021)
);

BUFx2_ASAP7_75t_L g5022 ( 
.A(n_4698),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4683),
.Y(n_5023)
);

AOI22xp5_ASAP7_75t_L g5024 ( 
.A1(n_4753),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_5024)
);

NAND2xp5_ASAP7_75t_L g5025 ( 
.A(n_4667),
.B(n_46),
.Y(n_5025)
);

AND2x2_ASAP7_75t_L g5026 ( 
.A(n_4758),
.B(n_47),
.Y(n_5026)
);

NAND2xp5_ASAP7_75t_L g5027 ( 
.A(n_4696),
.B(n_47),
.Y(n_5027)
);

INVx2_ASAP7_75t_L g5028 ( 
.A(n_4875),
.Y(n_5028)
);

INVx4_ASAP7_75t_L g5029 ( 
.A(n_4907),
.Y(n_5029)
);

NOR2xp33_ASAP7_75t_R g5030 ( 
.A(n_4689),
.B(n_4712),
.Y(n_5030)
);

BUFx3_ASAP7_75t_L g5031 ( 
.A(n_4750),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_4728),
.B(n_48),
.Y(n_5032)
);

BUFx6f_ASAP7_75t_L g5033 ( 
.A(n_4710),
.Y(n_5033)
);

AND2x2_ASAP7_75t_L g5034 ( 
.A(n_4950),
.B(n_48),
.Y(n_5034)
);

NAND2xp5_ASAP7_75t_L g5035 ( 
.A(n_4685),
.B(n_49),
.Y(n_5035)
);

INVx3_ASAP7_75t_L g5036 ( 
.A(n_4804),
.Y(n_5036)
);

BUFx3_ASAP7_75t_L g5037 ( 
.A(n_4857),
.Y(n_5037)
);

NOR2xp33_ASAP7_75t_R g5038 ( 
.A(n_4701),
.B(n_1815),
.Y(n_5038)
);

AND2x2_ASAP7_75t_L g5039 ( 
.A(n_4952),
.B(n_49),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4681),
.B(n_50),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_L g5041 ( 
.A(n_4731),
.B(n_51),
.Y(n_5041)
);

BUFx3_ASAP7_75t_L g5042 ( 
.A(n_4858),
.Y(n_5042)
);

OAI21xp5_ASAP7_75t_L g5043 ( 
.A1(n_4666),
.A2(n_51),
.B(n_52),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4718),
.Y(n_5044)
);

BUFx3_ASAP7_75t_L g5045 ( 
.A(n_4863),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4868),
.Y(n_5046)
);

NOR2x1p5_ASAP7_75t_SL g5047 ( 
.A(n_4686),
.B(n_1816),
.Y(n_5047)
);

NAND2xp5_ASAP7_75t_L g5048 ( 
.A(n_4734),
.B(n_4736),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_L g5049 ( 
.A(n_4740),
.B(n_52),
.Y(n_5049)
);

A2O1A1Ixp33_ASAP7_75t_L g5050 ( 
.A1(n_4899),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_5050)
);

OAI22xp5_ASAP7_75t_SL g5051 ( 
.A1(n_4929),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_5051)
);

AND2x2_ASAP7_75t_L g5052 ( 
.A(n_4953),
.B(n_56),
.Y(n_5052)
);

INVx1_ASAP7_75t_SL g5053 ( 
.A(n_4708),
.Y(n_5053)
);

INVx2_ASAP7_75t_L g5054 ( 
.A(n_4869),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_4743),
.B(n_57),
.Y(n_5055)
);

AND2x2_ASAP7_75t_L g5056 ( 
.A(n_4954),
.B(n_58),
.Y(n_5056)
);

BUFx6f_ASAP7_75t_L g5057 ( 
.A(n_4932),
.Y(n_5057)
);

INVx3_ASAP7_75t_L g5058 ( 
.A(n_4711),
.Y(n_5058)
);

BUFx8_ASAP7_75t_L g5059 ( 
.A(n_4788),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_4871),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4889),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_4955),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4747),
.B(n_58),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4956),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_4751),
.B(n_59),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4957),
.Y(n_5066)
);

INVx3_ASAP7_75t_L g5067 ( 
.A(n_4715),
.Y(n_5067)
);

INVx2_ASAP7_75t_L g5068 ( 
.A(n_4775),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_4756),
.B(n_59),
.Y(n_5069)
);

NAND2x1p5_ASAP7_75t_L g5070 ( 
.A(n_4679),
.B(n_1817),
.Y(n_5070)
);

BUFx6f_ASAP7_75t_L g5071 ( 
.A(n_4915),
.Y(n_5071)
);

AND3x1_ASAP7_75t_SL g5072 ( 
.A(n_4947),
.B(n_60),
.C(n_61),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_4675),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_4938),
.Y(n_5074)
);

AND2x2_ASAP7_75t_L g5075 ( 
.A(n_4660),
.B(n_60),
.Y(n_5075)
);

CKINVDCx5p33_ASAP7_75t_R g5076 ( 
.A(n_4737),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_4773),
.B(n_61),
.Y(n_5077)
);

INVx2_ASAP7_75t_L g5078 ( 
.A(n_4784),
.Y(n_5078)
);

OR2x6_ASAP7_75t_L g5079 ( 
.A(n_4934),
.B(n_1820),
.Y(n_5079)
);

INVxp67_ASAP7_75t_SL g5080 ( 
.A(n_4668),
.Y(n_5080)
);

AND3x1_ASAP7_75t_SL g5081 ( 
.A(n_4943),
.B(n_62),
.C(n_63),
.Y(n_5081)
);

OAI22xp5_ASAP7_75t_L g5082 ( 
.A1(n_4673),
.A2(n_4664),
.B1(n_4777),
.B2(n_4703),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_4669),
.B(n_63),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4716),
.Y(n_5084)
);

INVx3_ASAP7_75t_SL g5085 ( 
.A(n_4790),
.Y(n_5085)
);

NAND2xp33_ASAP7_75t_SL g5086 ( 
.A(n_4706),
.B(n_64),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4941),
.Y(n_5087)
);

AND2x2_ASAP7_75t_L g5088 ( 
.A(n_4828),
.B(n_64),
.Y(n_5088)
);

AND2x2_ASAP7_75t_L g5089 ( 
.A(n_4843),
.B(n_65),
.Y(n_5089)
);

NAND2xp33_ASAP7_75t_L g5090 ( 
.A(n_4719),
.B(n_66),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_4694),
.Y(n_5091)
);

AND2x2_ASAP7_75t_L g5092 ( 
.A(n_4898),
.B(n_67),
.Y(n_5092)
);

INVx2_ASAP7_75t_L g5093 ( 
.A(n_4721),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_4687),
.B(n_67),
.Y(n_5094)
);

INVx2_ASAP7_75t_SL g5095 ( 
.A(n_4707),
.Y(n_5095)
);

AND2x4_ASAP7_75t_L g5096 ( 
.A(n_4680),
.B(n_4916),
.Y(n_5096)
);

BUFx2_ASAP7_75t_L g5097 ( 
.A(n_4699),
.Y(n_5097)
);

INVx2_ASAP7_75t_L g5098 ( 
.A(n_4821),
.Y(n_5098)
);

AOI22x1_ASAP7_75t_L g5099 ( 
.A1(n_4688),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_5099)
);

BUFx3_ASAP7_75t_L g5100 ( 
.A(n_4910),
.Y(n_5100)
);

INVx2_ASAP7_75t_L g5101 ( 
.A(n_4824),
.Y(n_5101)
);

NAND2xp5_ASAP7_75t_L g5102 ( 
.A(n_4704),
.B(n_68),
.Y(n_5102)
);

AND2x2_ASAP7_75t_L g5103 ( 
.A(n_4901),
.B(n_70),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_4695),
.B(n_71),
.Y(n_5104)
);

NAND2x1p5_ASAP7_75t_L g5105 ( 
.A(n_4691),
.B(n_1821),
.Y(n_5105)
);

CKINVDCx5p33_ASAP7_75t_R g5106 ( 
.A(n_4912),
.Y(n_5106)
);

NAND2xp5_ASAP7_75t_L g5107 ( 
.A(n_4729),
.B(n_71),
.Y(n_5107)
);

AND2x2_ASAP7_75t_L g5108 ( 
.A(n_4909),
.B(n_72),
.Y(n_5108)
);

INVxp67_ASAP7_75t_L g5109 ( 
.A(n_4826),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_4830),
.Y(n_5110)
);

O2A1O1Ixp33_ASAP7_75t_L g5111 ( 
.A1(n_4914),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_4832),
.Y(n_5112)
);

INVx2_ASAP7_75t_L g5113 ( 
.A(n_4837),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_4705),
.B(n_73),
.Y(n_5114)
);

INVx2_ASAP7_75t_L g5115 ( 
.A(n_4838),
.Y(n_5115)
);

INVx2_ASAP7_75t_L g5116 ( 
.A(n_4841),
.Y(n_5116)
);

HB1xp67_ASAP7_75t_L g5117 ( 
.A(n_4891),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_4842),
.Y(n_5118)
);

BUFx6f_ASAP7_75t_L g5119 ( 
.A(n_4730),
.Y(n_5119)
);

NOR2xp33_ASAP7_75t_R g5120 ( 
.A(n_4661),
.B(n_1824),
.Y(n_5120)
);

INVxp33_ASAP7_75t_SL g5121 ( 
.A(n_4917),
.Y(n_5121)
);

NAND2x1p5_ASAP7_75t_L g5122 ( 
.A(n_4732),
.B(n_1832),
.Y(n_5122)
);

OAI22xp5_ASAP7_75t_L g5123 ( 
.A1(n_4674),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_5123)
);

AND2x2_ASAP7_75t_L g5124 ( 
.A(n_4884),
.B(n_75),
.Y(n_5124)
);

AND2x2_ASAP7_75t_L g5125 ( 
.A(n_4887),
.B(n_76),
.Y(n_5125)
);

OAI22xp5_ASAP7_75t_SL g5126 ( 
.A1(n_4855),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_5126)
);

INVx3_ASAP7_75t_L g5127 ( 
.A(n_4676),
.Y(n_5127)
);

BUFx12f_ASAP7_75t_L g5128 ( 
.A(n_4928),
.Y(n_5128)
);

INVx2_ASAP7_75t_L g5129 ( 
.A(n_4845),
.Y(n_5129)
);

INVx3_ASAP7_75t_L g5130 ( 
.A(n_4670),
.Y(n_5130)
);

BUFx2_ASAP7_75t_SL g5131 ( 
.A(n_4892),
.Y(n_5131)
);

INVx1_ASAP7_75t_L g5132 ( 
.A(n_4846),
.Y(n_5132)
);

NAND2xp5_ASAP7_75t_L g5133 ( 
.A(n_4720),
.B(n_77),
.Y(n_5133)
);

AND2x2_ASAP7_75t_L g5134 ( 
.A(n_4886),
.B(n_79),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_L g5135 ( 
.A(n_4779),
.B(n_80),
.Y(n_5135)
);

BUFx2_ASAP7_75t_L g5136 ( 
.A(n_4823),
.Y(n_5136)
);

INVx1_ASAP7_75t_L g5137 ( 
.A(n_4847),
.Y(n_5137)
);

NAND2x1_ASAP7_75t_L g5138 ( 
.A(n_4812),
.B(n_1834),
.Y(n_5138)
);

NAND2x1p5_ASAP7_75t_L g5139 ( 
.A(n_4742),
.B(n_1835),
.Y(n_5139)
);

BUFx2_ASAP7_75t_L g5140 ( 
.A(n_4816),
.Y(n_5140)
);

CKINVDCx5p33_ASAP7_75t_R g5141 ( 
.A(n_4883),
.Y(n_5141)
);

AOI22xp5_ASAP7_75t_L g5142 ( 
.A1(n_4717),
.A2(n_84),
.B1(n_81),
.B2(n_83),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_4848),
.Y(n_5143)
);

INVx2_ASAP7_75t_L g5144 ( 
.A(n_4849),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_4850),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_4852),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_L g5147 ( 
.A(n_4781),
.B(n_81),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_4853),
.Y(n_5148)
);

BUFx3_ASAP7_75t_L g5149 ( 
.A(n_4778),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_4854),
.Y(n_5150)
);

AOI22xp5_ASAP7_75t_L g5151 ( 
.A1(n_4933),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_5151)
);

INVx2_ASAP7_75t_L g5152 ( 
.A(n_4859),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_4782),
.B(n_85),
.Y(n_5153)
);

NAND2xp5_ASAP7_75t_L g5154 ( 
.A(n_4783),
.B(n_86),
.Y(n_5154)
);

INVx2_ASAP7_75t_L g5155 ( 
.A(n_4861),
.Y(n_5155)
);

INVx3_ASAP7_75t_SL g5156 ( 
.A(n_4741),
.Y(n_5156)
);

OAI21xp5_ASAP7_75t_L g5157 ( 
.A1(n_4755),
.A2(n_86),
.B(n_87),
.Y(n_5157)
);

NAND2xp5_ASAP7_75t_L g5158 ( 
.A(n_4785),
.B(n_88),
.Y(n_5158)
);

AOI22xp33_ASAP7_75t_L g5159 ( 
.A1(n_4939),
.A2(n_92),
.B1(n_88),
.B2(n_89),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_4862),
.Y(n_5160)
);

OAI22xp5_ASAP7_75t_L g5161 ( 
.A1(n_4697),
.A2(n_93),
.B1(n_89),
.B2(n_92),
.Y(n_5161)
);

INVx2_ASAP7_75t_L g5162 ( 
.A(n_4864),
.Y(n_5162)
);

BUFx6f_ASAP7_75t_L g5163 ( 
.A(n_4795),
.Y(n_5163)
);

INVx8_ASAP7_75t_L g5164 ( 
.A(n_4856),
.Y(n_5164)
);

CKINVDCx20_ASAP7_75t_R g5165 ( 
.A(n_4834),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_4865),
.Y(n_5166)
);

NAND2xp5_ASAP7_75t_L g5167 ( 
.A(n_4759),
.B(n_93),
.Y(n_5167)
);

BUFx12f_ASAP7_75t_L g5168 ( 
.A(n_4920),
.Y(n_5168)
);

AND2x2_ASAP7_75t_L g5169 ( 
.A(n_4902),
.B(n_95),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_4760),
.B(n_95),
.Y(n_5170)
);

AOI22xp33_ASAP7_75t_L g5171 ( 
.A1(n_4829),
.A2(n_4825),
.B1(n_4937),
.B2(n_4906),
.Y(n_5171)
);

HB1xp67_ASAP7_75t_L g5172 ( 
.A(n_4772),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_4776),
.Y(n_5173)
);

BUFx8_ASAP7_75t_L g5174 ( 
.A(n_4921),
.Y(n_5174)
);

INVx1_ASAP7_75t_L g5175 ( 
.A(n_4787),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_4762),
.B(n_96),
.Y(n_5176)
);

AOI21xp5_ASAP7_75t_L g5177 ( 
.A1(n_4770),
.A2(n_1837),
.B(n_1836),
.Y(n_5177)
);

NAND2xp5_ASAP7_75t_L g5178 ( 
.A(n_4764),
.B(n_96),
.Y(n_5178)
);

INVx2_ASAP7_75t_L g5179 ( 
.A(n_4739),
.Y(n_5179)
);

AOI22xp5_ASAP7_75t_L g5180 ( 
.A1(n_4878),
.A2(n_100),
.B1(n_97),
.B2(n_99),
.Y(n_5180)
);

INVxp67_ASAP7_75t_L g5181 ( 
.A(n_4757),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_SL g5182 ( 
.A(n_4749),
.B(n_97),
.Y(n_5182)
);

CKINVDCx20_ASAP7_75t_R g5183 ( 
.A(n_4835),
.Y(n_5183)
);

INVx2_ASAP7_75t_L g5184 ( 
.A(n_4797),
.Y(n_5184)
);

NAND2xp5_ASAP7_75t_SL g5185 ( 
.A(n_4723),
.B(n_100),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_4908),
.Y(n_5186)
);

BUFx8_ASAP7_75t_L g5187 ( 
.A(n_4922),
.Y(n_5187)
);

BUFx12f_ASAP7_75t_L g5188 ( 
.A(n_4839),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_4925),
.Y(n_5189)
);

NOR2x1p5_ASAP7_75t_SL g5190 ( 
.A(n_4890),
.B(n_1838),
.Y(n_5190)
);

AND2x2_ASAP7_75t_SL g5191 ( 
.A(n_4951),
.B(n_101),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_4798),
.Y(n_5192)
);

BUFx2_ASAP7_75t_L g5193 ( 
.A(n_5022),
.Y(n_5193)
);

AO21x2_ASAP7_75t_L g5194 ( 
.A1(n_5030),
.A2(n_4949),
.B(n_4900),
.Y(n_5194)
);

INVx1_ASAP7_75t_SL g5195 ( 
.A(n_5031),
.Y(n_5195)
);

BUFx3_ASAP7_75t_L g5196 ( 
.A(n_4972),
.Y(n_5196)
);

BUFx10_ASAP7_75t_L g5197 ( 
.A(n_5106),
.Y(n_5197)
);

INVx2_ASAP7_75t_L g5198 ( 
.A(n_4960),
.Y(n_5198)
);

OAI21x1_ASAP7_75t_L g5199 ( 
.A1(n_5044),
.A2(n_4926),
.B(n_4923),
.Y(n_5199)
);

BUFx3_ASAP7_75t_L g5200 ( 
.A(n_4961),
.Y(n_5200)
);

OAI21x1_ASAP7_75t_L g5201 ( 
.A1(n_5084),
.A2(n_5091),
.B(n_5093),
.Y(n_5201)
);

AO21x2_ASAP7_75t_L g5202 ( 
.A1(n_5157),
.A2(n_4771),
.B(n_4735),
.Y(n_5202)
);

OAI21x1_ASAP7_75t_L g5203 ( 
.A1(n_5138),
.A2(n_4811),
.B(n_4769),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_4965),
.Y(n_5204)
);

AO21x2_ASAP7_75t_L g5205 ( 
.A1(n_5120),
.A2(n_4793),
.B(n_4885),
.Y(n_5205)
);

INVx1_ASAP7_75t_SL g5206 ( 
.A(n_5003),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_4963),
.Y(n_5207)
);

AND2x4_ASAP7_75t_L g5208 ( 
.A(n_4991),
.B(n_4796),
.Y(n_5208)
);

OAI21xp5_ASAP7_75t_L g5209 ( 
.A1(n_5082),
.A2(n_4880),
.B(n_4726),
.Y(n_5209)
);

BUFx6f_ASAP7_75t_L g5210 ( 
.A(n_4994),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_4964),
.Y(n_5211)
);

OAI21x1_ASAP7_75t_L g5212 ( 
.A1(n_5105),
.A2(n_4802),
.B(n_4799),
.Y(n_5212)
);

INVx2_ASAP7_75t_L g5213 ( 
.A(n_5012),
.Y(n_5213)
);

BUFx3_ASAP7_75t_L g5214 ( 
.A(n_4993),
.Y(n_5214)
);

INVx2_ASAP7_75t_SL g5215 ( 
.A(n_5000),
.Y(n_5215)
);

AO21x2_ASAP7_75t_L g5216 ( 
.A1(n_5043),
.A2(n_4808),
.B(n_4805),
.Y(n_5216)
);

BUFx12f_ASAP7_75t_L g5217 ( 
.A(n_5059),
.Y(n_5217)
);

OAI21x1_ASAP7_75t_L g5218 ( 
.A1(n_5177),
.A2(n_4820),
.B(n_4918),
.Y(n_5218)
);

AOI22x1_ASAP7_75t_L g5219 ( 
.A1(n_5097),
.A2(n_4722),
.B1(n_4874),
.B2(n_4833),
.Y(n_5219)
);

AO21x2_ASAP7_75t_L g5220 ( 
.A1(n_5040),
.A2(n_4792),
.B(n_4919),
.Y(n_5220)
);

INVx2_ASAP7_75t_SL g5221 ( 
.A(n_5057),
.Y(n_5221)
);

INVx2_ASAP7_75t_L g5222 ( 
.A(n_5016),
.Y(n_5222)
);

BUFx3_ASAP7_75t_L g5223 ( 
.A(n_5057),
.Y(n_5223)
);

BUFx3_ASAP7_75t_L g5224 ( 
.A(n_5020),
.Y(n_5224)
);

INVx3_ASAP7_75t_L g5225 ( 
.A(n_4994),
.Y(n_5225)
);

NAND2x1p5_ASAP7_75t_L g5226 ( 
.A(n_5127),
.B(n_4724),
.Y(n_5226)
);

INVx2_ASAP7_75t_SL g5227 ( 
.A(n_4985),
.Y(n_5227)
);

BUFx4f_ASAP7_75t_SL g5228 ( 
.A(n_5188),
.Y(n_5228)
);

BUFx6f_ASAP7_75t_L g5229 ( 
.A(n_5033),
.Y(n_5229)
);

INVx5_ASAP7_75t_L g5230 ( 
.A(n_5168),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_5023),
.Y(n_5231)
);

AND2x6_ASAP7_75t_L g5232 ( 
.A(n_5096),
.B(n_4860),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5073),
.Y(n_5233)
);

AOI22x1_ASAP7_75t_L g5234 ( 
.A1(n_5018),
.A2(n_4831),
.B1(n_4754),
.B2(n_4765),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_5002),
.Y(n_5235)
);

INVx2_ASAP7_75t_L g5236 ( 
.A(n_4967),
.Y(n_5236)
);

INVx3_ASAP7_75t_L g5237 ( 
.A(n_5033),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_5080),
.Y(n_5238)
);

INVx1_ASAP7_75t_SL g5239 ( 
.A(n_5053),
.Y(n_5239)
);

INVxp67_ASAP7_75t_SL g5240 ( 
.A(n_5058),
.Y(n_5240)
);

OR2x2_ASAP7_75t_L g5241 ( 
.A(n_5067),
.B(n_4894),
.Y(n_5241)
);

AO21x2_ASAP7_75t_L g5242 ( 
.A1(n_4990),
.A2(n_4913),
.B(n_4911),
.Y(n_5242)
);

AND2x2_ASAP7_75t_L g5243 ( 
.A(n_4966),
.B(n_4818),
.Y(n_5243)
);

NAND2xp5_ASAP7_75t_L g5244 ( 
.A(n_4992),
.B(n_4895),
.Y(n_5244)
);

INVx2_ASAP7_75t_SL g5245 ( 
.A(n_5119),
.Y(n_5245)
);

NOR2xp33_ASAP7_75t_L g5246 ( 
.A(n_4959),
.B(n_4752),
.Y(n_5246)
);

OAI21x1_ASAP7_75t_L g5247 ( 
.A1(n_5130),
.A2(n_4819),
.B(n_4903),
.Y(n_5247)
);

INVxp67_ASAP7_75t_SL g5248 ( 
.A(n_4975),
.Y(n_5248)
);

OAI21x1_ASAP7_75t_L g5249 ( 
.A1(n_5004),
.A2(n_4904),
.B(n_4866),
.Y(n_5249)
);

INVx2_ASAP7_75t_SL g5250 ( 
.A(n_5119),
.Y(n_5250)
);

INVx2_ASAP7_75t_L g5251 ( 
.A(n_4978),
.Y(n_5251)
);

OAI21x1_ASAP7_75t_L g5252 ( 
.A1(n_5099),
.A2(n_4814),
.B(n_4813),
.Y(n_5252)
);

NOR2xp33_ASAP7_75t_L g5253 ( 
.A(n_5121),
.B(n_4872),
.Y(n_5253)
);

AO21x2_ASAP7_75t_L g5254 ( 
.A1(n_5083),
.A2(n_4877),
.B(n_4876),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_4973),
.Y(n_5255)
);

OA21x2_ASAP7_75t_L g5256 ( 
.A1(n_5087),
.A2(n_4927),
.B(n_4905),
.Y(n_5256)
);

OAI21x1_ASAP7_75t_L g5257 ( 
.A1(n_5019),
.A2(n_5122),
.B(n_5070),
.Y(n_5257)
);

OAI21x1_ASAP7_75t_L g5258 ( 
.A1(n_4998),
.A2(n_4897),
.B(n_4896),
.Y(n_5258)
);

AO21x2_ASAP7_75t_L g5259 ( 
.A1(n_5025),
.A2(n_5094),
.B(n_5032),
.Y(n_5259)
);

INVx1_ASAP7_75t_SL g5260 ( 
.A(n_5036),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_5009),
.Y(n_5261)
);

OAI21x1_ASAP7_75t_L g5262 ( 
.A1(n_4987),
.A2(n_4893),
.B(n_4766),
.Y(n_5262)
);

OAI21x1_ASAP7_75t_L g5263 ( 
.A1(n_4989),
.A2(n_4767),
.B(n_4761),
.Y(n_5263)
);

AO21x1_ASAP7_75t_SL g5264 ( 
.A1(n_5062),
.A2(n_4780),
.B(n_4768),
.Y(n_5264)
);

OAI21xp5_ASAP7_75t_L g5265 ( 
.A1(n_5048),
.A2(n_4794),
.B(n_4791),
.Y(n_5265)
);

OAI21xp5_ASAP7_75t_L g5266 ( 
.A1(n_4984),
.A2(n_4801),
.B(n_4800),
.Y(n_5266)
);

INVx2_ASAP7_75t_SL g5267 ( 
.A(n_5163),
.Y(n_5267)
);

AO21x2_ASAP7_75t_L g5268 ( 
.A1(n_4988),
.A2(n_5021),
.B(n_5102),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_5064),
.Y(n_5269)
);

BUFx6f_ASAP7_75t_L g5270 ( 
.A(n_5163),
.Y(n_5270)
);

AOI22x1_ASAP7_75t_L g5271 ( 
.A1(n_4971),
.A2(n_4806),
.B1(n_104),
.B2(n_102),
.Y(n_5271)
);

OAI21x1_ASAP7_75t_L g5272 ( 
.A1(n_5139),
.A2(n_1840),
.B(n_1839),
.Y(n_5272)
);

AND2x2_ASAP7_75t_L g5273 ( 
.A(n_5075),
.B(n_1841),
.Y(n_5273)
);

AO21x2_ASAP7_75t_L g5274 ( 
.A1(n_5027),
.A2(n_103),
.B(n_104),
.Y(n_5274)
);

BUFx2_ASAP7_75t_SL g5275 ( 
.A(n_5008),
.Y(n_5275)
);

OAI21x1_ASAP7_75t_L g5276 ( 
.A1(n_4974),
.A2(n_1843),
.B(n_1842),
.Y(n_5276)
);

INVx3_ASAP7_75t_L g5277 ( 
.A(n_5071),
.Y(n_5277)
);

OAI21x1_ASAP7_75t_L g5278 ( 
.A1(n_4995),
.A2(n_1845),
.B(n_1844),
.Y(n_5278)
);

INVx6_ASAP7_75t_L g5279 ( 
.A(n_5174),
.Y(n_5279)
);

AND2x4_ASAP7_75t_L g5280 ( 
.A(n_4996),
.B(n_1846),
.Y(n_5280)
);

NAND2x1p5_ASAP7_75t_L g5281 ( 
.A(n_5017),
.B(n_5037),
.Y(n_5281)
);

INVx5_ASAP7_75t_SL g5282 ( 
.A(n_5071),
.Y(n_5282)
);

AO21x2_ASAP7_75t_L g5283 ( 
.A1(n_5035),
.A2(n_103),
.B(n_105),
.Y(n_5283)
);

INVx4_ASAP7_75t_L g5284 ( 
.A(n_5128),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_5066),
.Y(n_5285)
);

BUFx12f_ASAP7_75t_L g5286 ( 
.A(n_5014),
.Y(n_5286)
);

OR2x2_ASAP7_75t_L g5287 ( 
.A(n_4977),
.B(n_106),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_5104),
.Y(n_5288)
);

AO21x2_ASAP7_75t_L g5289 ( 
.A1(n_4983),
.A2(n_106),
.B(n_107),
.Y(n_5289)
);

BUFx2_ASAP7_75t_R g5290 ( 
.A(n_4997),
.Y(n_5290)
);

HB1xp67_ASAP7_75t_L g5291 ( 
.A(n_5095),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_5074),
.Y(n_5292)
);

INVx5_ASAP7_75t_L g5293 ( 
.A(n_5164),
.Y(n_5293)
);

NAND2xp5_ASAP7_75t_SL g5294 ( 
.A(n_5068),
.B(n_1848),
.Y(n_5294)
);

OAI21x1_ASAP7_75t_L g5295 ( 
.A1(n_5171),
.A2(n_1850),
.B(n_1849),
.Y(n_5295)
);

BUFx2_ASAP7_75t_L g5296 ( 
.A(n_5042),
.Y(n_5296)
);

INVx6_ASAP7_75t_L g5297 ( 
.A(n_5187),
.Y(n_5297)
);

AO21x2_ASAP7_75t_L g5298 ( 
.A1(n_5038),
.A2(n_108),
.B(n_109),
.Y(n_5298)
);

OAI21x1_ASAP7_75t_L g5299 ( 
.A1(n_5114),
.A2(n_1852),
.B(n_1851),
.Y(n_5299)
);

NAND2x1p5_ASAP7_75t_L g5300 ( 
.A(n_5045),
.B(n_1855),
.Y(n_5300)
);

BUFx3_ASAP7_75t_L g5301 ( 
.A(n_5149),
.Y(n_5301)
);

AO21x2_ASAP7_75t_L g5302 ( 
.A1(n_5090),
.A2(n_109),
.B(n_110),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_5133),
.Y(n_5303)
);

BUFx12f_ASAP7_75t_L g5304 ( 
.A(n_5076),
.Y(n_5304)
);

INVx2_ASAP7_75t_L g5305 ( 
.A(n_4980),
.Y(n_5305)
);

INVx4_ASAP7_75t_L g5306 ( 
.A(n_5164),
.Y(n_5306)
);

BUFx10_ASAP7_75t_L g5307 ( 
.A(n_5141),
.Y(n_5307)
);

AO21x2_ASAP7_75t_L g5308 ( 
.A1(n_5001),
.A2(n_110),
.B(n_111),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_4981),
.Y(n_5309)
);

AO21x2_ASAP7_75t_L g5310 ( 
.A1(n_5050),
.A2(n_111),
.B(n_112),
.Y(n_5310)
);

INVx1_ASAP7_75t_SL g5311 ( 
.A(n_5156),
.Y(n_5311)
);

BUFx6f_ASAP7_75t_L g5312 ( 
.A(n_5085),
.Y(n_5312)
);

BUFx3_ASAP7_75t_L g5313 ( 
.A(n_5183),
.Y(n_5313)
);

BUFx6f_ASAP7_75t_L g5314 ( 
.A(n_5005),
.Y(n_5314)
);

OAI22xp33_ASAP7_75t_L g5315 ( 
.A1(n_5151),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_5315)
);

BUFx6f_ASAP7_75t_L g5316 ( 
.A(n_5010),
.Y(n_5316)
);

OR3x4_ASAP7_75t_SL g5317 ( 
.A(n_4976),
.B(n_113),
.C(n_114),
.Y(n_5317)
);

BUFx6f_ASAP7_75t_L g5318 ( 
.A(n_5026),
.Y(n_5318)
);

BUFx2_ASAP7_75t_L g5319 ( 
.A(n_5172),
.Y(n_5319)
);

AO21x2_ASAP7_75t_L g5320 ( 
.A1(n_5107),
.A2(n_115),
.B(n_116),
.Y(n_5320)
);

BUFx3_ASAP7_75t_L g5321 ( 
.A(n_5165),
.Y(n_5321)
);

AO21x2_ASAP7_75t_L g5322 ( 
.A1(n_5041),
.A2(n_5055),
.B(n_5049),
.Y(n_5322)
);

NAND2x1p5_ASAP7_75t_L g5323 ( 
.A(n_5140),
.B(n_1856),
.Y(n_5323)
);

AND2x4_ASAP7_75t_L g5324 ( 
.A(n_5079),
.B(n_1859),
.Y(n_5324)
);

INVx2_ASAP7_75t_L g5325 ( 
.A(n_5078),
.Y(n_5325)
);

NOR2xp33_ASAP7_75t_L g5326 ( 
.A(n_5109),
.B(n_1860),
.Y(n_5326)
);

BUFx2_ASAP7_75t_SL g5327 ( 
.A(n_5117),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_5006),
.Y(n_5328)
);

INVx3_ASAP7_75t_L g5329 ( 
.A(n_5029),
.Y(n_5329)
);

AND2x4_ASAP7_75t_L g5330 ( 
.A(n_5079),
.B(n_1861),
.Y(n_5330)
);

INVx3_ASAP7_75t_L g5331 ( 
.A(n_5098),
.Y(n_5331)
);

OAI21xp5_ASAP7_75t_L g5332 ( 
.A1(n_4979),
.A2(n_115),
.B(n_116),
.Y(n_5332)
);

OAI21x1_ASAP7_75t_L g5333 ( 
.A1(n_5046),
.A2(n_1863),
.B(n_1862),
.Y(n_5333)
);

NAND2xp5_ASAP7_75t_L g5334 ( 
.A(n_5100),
.B(n_117),
.Y(n_5334)
);

BUFx3_ASAP7_75t_L g5335 ( 
.A(n_5136),
.Y(n_5335)
);

BUFx4f_ASAP7_75t_L g5336 ( 
.A(n_5192),
.Y(n_5336)
);

NOR2xp33_ASAP7_75t_L g5337 ( 
.A(n_5181),
.B(n_1865),
.Y(n_5337)
);

INVx2_ASAP7_75t_L g5338 ( 
.A(n_5054),
.Y(n_5338)
);

INVx2_ASAP7_75t_L g5339 ( 
.A(n_5028),
.Y(n_5339)
);

INVx6_ASAP7_75t_L g5340 ( 
.A(n_4970),
.Y(n_5340)
);

AO21x2_ASAP7_75t_L g5341 ( 
.A1(n_5063),
.A2(n_118),
.B(n_119),
.Y(n_5341)
);

INVx3_ASAP7_75t_L g5342 ( 
.A(n_5101),
.Y(n_5342)
);

AO21x1_ASAP7_75t_L g5343 ( 
.A1(n_5086),
.A2(n_119),
.B(n_120),
.Y(n_5343)
);

OA21x2_ASAP7_75t_L g5344 ( 
.A1(n_5135),
.A2(n_121),
.B(n_122),
.Y(n_5344)
);

AO21x2_ASAP7_75t_L g5345 ( 
.A1(n_5065),
.A2(n_123),
.B(n_124),
.Y(n_5345)
);

AO21x2_ASAP7_75t_L g5346 ( 
.A1(n_5069),
.A2(n_123),
.B(n_124),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5186),
.Y(n_5347)
);

OR3x4_ASAP7_75t_SL g5348 ( 
.A(n_4969),
.B(n_125),
.C(n_126),
.Y(n_5348)
);

INVx2_ASAP7_75t_SL g5349 ( 
.A(n_5113),
.Y(n_5349)
);

BUFx3_ASAP7_75t_L g5350 ( 
.A(n_5184),
.Y(n_5350)
);

INVx1_ASAP7_75t_SL g5351 ( 
.A(n_5131),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5110),
.Y(n_5352)
);

NOR2x1_ASAP7_75t_R g5353 ( 
.A(n_5185),
.B(n_1866),
.Y(n_5353)
);

BUFx2_ASAP7_75t_R g5354 ( 
.A(n_5182),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_5112),
.Y(n_5355)
);

INVx2_ASAP7_75t_L g5356 ( 
.A(n_5060),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_5204),
.Y(n_5357)
);

AOI22xp33_ASAP7_75t_SL g5358 ( 
.A1(n_5332),
.A2(n_5191),
.B1(n_5051),
.B2(n_5126),
.Y(n_5358)
);

AOI22xp33_ASAP7_75t_SL g5359 ( 
.A1(n_5271),
.A2(n_5161),
.B1(n_4968),
.B2(n_5123),
.Y(n_5359)
);

INVx2_ASAP7_75t_L g5360 ( 
.A(n_5213),
.Y(n_5360)
);

AOI22xp33_ASAP7_75t_L g5361 ( 
.A1(n_5343),
.A2(n_4962),
.B1(n_4999),
.B2(n_5011),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_5292),
.Y(n_5362)
);

OAI22xp5_ASAP7_75t_L g5363 ( 
.A1(n_5354),
.A2(n_5015),
.B1(n_5142),
.B2(n_5024),
.Y(n_5363)
);

CKINVDCx11_ASAP7_75t_R g5364 ( 
.A(n_5217),
.Y(n_5364)
);

BUFx3_ASAP7_75t_L g5365 ( 
.A(n_5196),
.Y(n_5365)
);

OAI22xp33_ASAP7_75t_L g5366 ( 
.A1(n_5209),
.A2(n_5180),
.B1(n_5077),
.B2(n_5153),
.Y(n_5366)
);

CKINVDCx11_ASAP7_75t_R g5367 ( 
.A(n_5307),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5248),
.Y(n_5368)
);

AOI22xp5_ASAP7_75t_L g5369 ( 
.A1(n_5266),
.A2(n_4982),
.B1(n_5072),
.B2(n_5103),
.Y(n_5369)
);

INVx1_ASAP7_75t_L g5370 ( 
.A(n_5233),
.Y(n_5370)
);

INVx6_ASAP7_75t_L g5371 ( 
.A(n_5293),
.Y(n_5371)
);

CKINVDCx5p33_ASAP7_75t_R g5372 ( 
.A(n_5286),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_L g5373 ( 
.A(n_5240),
.B(n_5088),
.Y(n_5373)
);

BUFx2_ASAP7_75t_SL g5374 ( 
.A(n_5293),
.Y(n_5374)
);

OAI22xp33_ASAP7_75t_L g5375 ( 
.A1(n_5336),
.A2(n_5154),
.B1(n_5158),
.B2(n_5147),
.Y(n_5375)
);

INVx1_ASAP7_75t_L g5376 ( 
.A(n_5231),
.Y(n_5376)
);

AOI22xp33_ASAP7_75t_SL g5377 ( 
.A1(n_5298),
.A2(n_5169),
.B1(n_5125),
.B2(n_5134),
.Y(n_5377)
);

INVx6_ASAP7_75t_L g5378 ( 
.A(n_5306),
.Y(n_5378)
);

OAI22xp5_ASAP7_75t_L g5379 ( 
.A1(n_5351),
.A2(n_5159),
.B1(n_5170),
.B2(n_5167),
.Y(n_5379)
);

BUFx3_ASAP7_75t_L g5380 ( 
.A(n_5270),
.Y(n_5380)
);

BUFx10_ASAP7_75t_L g5381 ( 
.A(n_5279),
.Y(n_5381)
);

BUFx8_ASAP7_75t_SL g5382 ( 
.A(n_5304),
.Y(n_5382)
);

CKINVDCx11_ASAP7_75t_R g5383 ( 
.A(n_5197),
.Y(n_5383)
);

INVx2_ASAP7_75t_L g5384 ( 
.A(n_5222),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_5269),
.Y(n_5385)
);

AOI22xp33_ASAP7_75t_L g5386 ( 
.A1(n_5315),
.A2(n_5124),
.B1(n_5179),
.B2(n_4986),
.Y(n_5386)
);

AOI22xp33_ASAP7_75t_L g5387 ( 
.A1(n_5302),
.A2(n_5089),
.B1(n_5175),
.B2(n_5173),
.Y(n_5387)
);

INVx3_ASAP7_75t_L g5388 ( 
.A(n_5229),
.Y(n_5388)
);

OAI22xp33_ASAP7_75t_L g5389 ( 
.A1(n_5317),
.A2(n_5178),
.B1(n_5176),
.B2(n_5189),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_5238),
.B(n_5034),
.Y(n_5390)
);

AOI22xp5_ASAP7_75t_L g5391 ( 
.A1(n_5205),
.A2(n_5081),
.B1(n_5007),
.B2(n_5118),
.Y(n_5391)
);

INVx6_ASAP7_75t_L g5392 ( 
.A(n_5230),
.Y(n_5392)
);

INVx6_ASAP7_75t_L g5393 ( 
.A(n_5230),
.Y(n_5393)
);

INVx1_ASAP7_75t_L g5394 ( 
.A(n_5285),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_5347),
.Y(n_5395)
);

AOI22xp33_ASAP7_75t_L g5396 ( 
.A1(n_5202),
.A2(n_5137),
.B1(n_5143),
.B2(n_5132),
.Y(n_5396)
);

BUFx12f_ASAP7_75t_L g5397 ( 
.A(n_5312),
.Y(n_5397)
);

AOI22xp33_ASAP7_75t_SL g5398 ( 
.A1(n_5310),
.A2(n_5039),
.B1(n_5056),
.B2(n_5052),
.Y(n_5398)
);

BUFx12f_ASAP7_75t_L g5399 ( 
.A(n_5210),
.Y(n_5399)
);

INVx2_ASAP7_75t_L g5400 ( 
.A(n_5211),
.Y(n_5400)
);

BUFx6f_ASAP7_75t_L g5401 ( 
.A(n_5223),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5352),
.Y(n_5402)
);

OAI22xp5_ASAP7_75t_L g5403 ( 
.A1(n_5193),
.A2(n_5061),
.B1(n_5146),
.B2(n_5145),
.Y(n_5403)
);

OAI22xp33_ASAP7_75t_L g5404 ( 
.A1(n_5311),
.A2(n_5150),
.B1(n_5160),
.B2(n_5148),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5355),
.Y(n_5405)
);

AOI22xp33_ASAP7_75t_SL g5406 ( 
.A1(n_5265),
.A2(n_5092),
.B1(n_5108),
.B2(n_5166),
.Y(n_5406)
);

INVx2_ASAP7_75t_L g5407 ( 
.A(n_5356),
.Y(n_5407)
);

INVx3_ASAP7_75t_L g5408 ( 
.A(n_5301),
.Y(n_5408)
);

BUFx2_ASAP7_75t_L g5409 ( 
.A(n_5335),
.Y(n_5409)
);

AOI22xp33_ASAP7_75t_SL g5410 ( 
.A1(n_5324),
.A2(n_5115),
.B1(n_5129),
.B2(n_5116),
.Y(n_5410)
);

CKINVDCx11_ASAP7_75t_R g5411 ( 
.A(n_5224),
.Y(n_5411)
);

OAI22xp5_ASAP7_75t_L g5412 ( 
.A1(n_5226),
.A2(n_5152),
.B1(n_5155),
.B2(n_5144),
.Y(n_5412)
);

INVx2_ASAP7_75t_SL g5413 ( 
.A(n_5277),
.Y(n_5413)
);

INVx2_ASAP7_75t_L g5414 ( 
.A(n_5236),
.Y(n_5414)
);

AOI22xp33_ASAP7_75t_L g5415 ( 
.A1(n_5242),
.A2(n_5162),
.B1(n_5013),
.B2(n_5111),
.Y(n_5415)
);

OAI21xp5_ASAP7_75t_SL g5416 ( 
.A1(n_5330),
.A2(n_5047),
.B(n_5190),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_5235),
.Y(n_5417)
);

AOI22xp33_ASAP7_75t_L g5418 ( 
.A1(n_5219),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_5418)
);

AOI22xp33_ASAP7_75t_L g5419 ( 
.A1(n_5216),
.A2(n_130),
.B1(n_127),
.B2(n_129),
.Y(n_5419)
);

INVx2_ASAP7_75t_L g5420 ( 
.A(n_5251),
.Y(n_5420)
);

INVx2_ASAP7_75t_L g5421 ( 
.A(n_5305),
.Y(n_5421)
);

INVxp67_ASAP7_75t_SL g5422 ( 
.A(n_5201),
.Y(n_5422)
);

HB1xp67_ASAP7_75t_L g5423 ( 
.A(n_5319),
.Y(n_5423)
);

INVx2_ASAP7_75t_L g5424 ( 
.A(n_5309),
.Y(n_5424)
);

INVx1_ASAP7_75t_SL g5425 ( 
.A(n_5195),
.Y(n_5425)
);

INVx1_ASAP7_75t_L g5426 ( 
.A(n_5198),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_5325),
.Y(n_5427)
);

AOI22xp33_ASAP7_75t_L g5428 ( 
.A1(n_5234),
.A2(n_5194),
.B1(n_5259),
.B2(n_5268),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_5207),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_5261),
.Y(n_5430)
);

CKINVDCx6p67_ASAP7_75t_R g5431 ( 
.A(n_5313),
.Y(n_5431)
);

INVxp67_ASAP7_75t_L g5432 ( 
.A(n_5296),
.Y(n_5432)
);

BUFx2_ASAP7_75t_SL g5433 ( 
.A(n_5215),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_5339),
.Y(n_5434)
);

INVx4_ASAP7_75t_L g5435 ( 
.A(n_5316),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_5338),
.Y(n_5436)
);

INVx1_ASAP7_75t_L g5437 ( 
.A(n_5327),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_5331),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5255),
.Y(n_5439)
);

INVx2_ASAP7_75t_L g5440 ( 
.A(n_5342),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_5288),
.Y(n_5441)
);

OAI22xp5_ASAP7_75t_L g5442 ( 
.A1(n_5239),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_5442)
);

OAI22xp5_ASAP7_75t_L g5443 ( 
.A1(n_5253),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_5443)
);

AOI22xp33_ASAP7_75t_L g5444 ( 
.A1(n_5246),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_5444)
);

INVx11_ASAP7_75t_L g5445 ( 
.A(n_5232),
.Y(n_5445)
);

INVx2_ASAP7_75t_L g5446 ( 
.A(n_5349),
.Y(n_5446)
);

OAI22xp33_ASAP7_75t_L g5447 ( 
.A1(n_5348),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_5447)
);

AND2x2_ASAP7_75t_L g5448 ( 
.A(n_5243),
.B(n_136),
.Y(n_5448)
);

BUFx4f_ASAP7_75t_SL g5449 ( 
.A(n_5321),
.Y(n_5449)
);

AOI22xp5_ASAP7_75t_L g5450 ( 
.A1(n_5232),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_5450)
);

INVx3_ASAP7_75t_L g5451 ( 
.A(n_5214),
.Y(n_5451)
);

OAI22xp33_ASAP7_75t_L g5452 ( 
.A1(n_5323),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_5452)
);

BUFx8_ASAP7_75t_L g5453 ( 
.A(n_5318),
.Y(n_5453)
);

BUFx2_ASAP7_75t_L g5454 ( 
.A(n_5281),
.Y(n_5454)
);

OAI22x1_ASAP7_75t_L g5455 ( 
.A1(n_5303),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_5455)
);

AOI22xp33_ASAP7_75t_SL g5456 ( 
.A1(n_5341),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_5456)
);

INVx1_ASAP7_75t_SL g5457 ( 
.A(n_5260),
.Y(n_5457)
);

INVx2_ASAP7_75t_L g5458 ( 
.A(n_5350),
.Y(n_5458)
);

BUFx3_ASAP7_75t_L g5459 ( 
.A(n_5267),
.Y(n_5459)
);

OAI22xp33_ASAP7_75t_L g5460 ( 
.A1(n_5329),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_5460)
);

OR2x2_ASAP7_75t_L g5461 ( 
.A(n_5328),
.B(n_145),
.Y(n_5461)
);

AOI22xp33_ASAP7_75t_L g5462 ( 
.A1(n_5322),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_5462)
);

OAI22xp5_ASAP7_75t_L g5463 ( 
.A1(n_5340),
.A2(n_150),
.B1(n_147),
.B2(n_149),
.Y(n_5463)
);

BUFx6f_ASAP7_75t_L g5464 ( 
.A(n_5200),
.Y(n_5464)
);

CKINVDCx14_ASAP7_75t_R g5465 ( 
.A(n_5297),
.Y(n_5465)
);

CKINVDCx5p33_ASAP7_75t_R g5466 ( 
.A(n_5290),
.Y(n_5466)
);

CKINVDCx11_ASAP7_75t_R g5467 ( 
.A(n_5314),
.Y(n_5467)
);

INVx6_ASAP7_75t_L g5468 ( 
.A(n_5284),
.Y(n_5468)
);

AOI22xp33_ASAP7_75t_L g5469 ( 
.A1(n_5220),
.A2(n_153),
.B1(n_149),
.B2(n_151),
.Y(n_5469)
);

AOI22xp33_ASAP7_75t_SL g5470 ( 
.A1(n_5345),
.A2(n_154),
.B1(n_151),
.B2(n_153),
.Y(n_5470)
);

AOI22xp33_ASAP7_75t_L g5471 ( 
.A1(n_5346),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_5291),
.Y(n_5472)
);

INVx2_ASAP7_75t_L g5473 ( 
.A(n_5237),
.Y(n_5473)
);

AOI22xp33_ASAP7_75t_SL g5474 ( 
.A1(n_5289),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_5474)
);

BUFx10_ASAP7_75t_L g5475 ( 
.A(n_5326),
.Y(n_5475)
);

OAI21xp33_ASAP7_75t_L g5476 ( 
.A1(n_5334),
.A2(n_158),
.B(n_161),
.Y(n_5476)
);

CKINVDCx20_ASAP7_75t_R g5477 ( 
.A(n_5228),
.Y(n_5477)
);

AOI22xp33_ASAP7_75t_L g5478 ( 
.A1(n_5320),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_5478)
);

HB1xp67_ASAP7_75t_L g5479 ( 
.A(n_5206),
.Y(n_5479)
);

AOI22xp5_ASAP7_75t_L g5480 ( 
.A1(n_5208),
.A2(n_167),
.B1(n_164),
.B2(n_165),
.Y(n_5480)
);

INVx2_ASAP7_75t_L g5481 ( 
.A(n_5241),
.Y(n_5481)
);

OR2x2_ASAP7_75t_SL g5482 ( 
.A(n_5344),
.B(n_165),
.Y(n_5482)
);

BUFx3_ASAP7_75t_L g5483 ( 
.A(n_5245),
.Y(n_5483)
);

CKINVDCx20_ASAP7_75t_R g5484 ( 
.A(n_5282),
.Y(n_5484)
);

AOI22xp33_ASAP7_75t_L g5485 ( 
.A1(n_5337),
.A2(n_170),
.B1(n_167),
.B2(n_168),
.Y(n_5485)
);

AOI22xp33_ASAP7_75t_SL g5486 ( 
.A1(n_5274),
.A2(n_171),
.B1(n_168),
.B2(n_170),
.Y(n_5486)
);

INVx2_ASAP7_75t_SL g5487 ( 
.A(n_5250),
.Y(n_5487)
);

AOI22xp33_ASAP7_75t_L g5488 ( 
.A1(n_5308),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_5488)
);

BUFx6f_ASAP7_75t_L g5489 ( 
.A(n_5221),
.Y(n_5489)
);

INVxp67_ASAP7_75t_SL g5490 ( 
.A(n_5263),
.Y(n_5490)
);

INVxp67_ASAP7_75t_SL g5491 ( 
.A(n_5262),
.Y(n_5491)
);

CKINVDCx20_ASAP7_75t_R g5492 ( 
.A(n_5227),
.Y(n_5492)
);

INVx2_ASAP7_75t_SL g5493 ( 
.A(n_5225),
.Y(n_5493)
);

OAI22xp33_ASAP7_75t_L g5494 ( 
.A1(n_5287),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_5494)
);

HB1xp67_ASAP7_75t_L g5495 ( 
.A(n_5283),
.Y(n_5495)
);

AO22x1_ASAP7_75t_L g5496 ( 
.A1(n_5244),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_5496)
);

CKINVDCx20_ASAP7_75t_R g5497 ( 
.A(n_5273),
.Y(n_5497)
);

AOI22xp5_ASAP7_75t_L g5498 ( 
.A1(n_5254),
.A2(n_178),
.B1(n_175),
.B2(n_176),
.Y(n_5498)
);

OAI22xp33_ASAP7_75t_L g5499 ( 
.A1(n_5300),
.A2(n_181),
.B1(n_178),
.B2(n_180),
.Y(n_5499)
);

INVx3_ASAP7_75t_L g5500 ( 
.A(n_5280),
.Y(n_5500)
);

INVx2_ASAP7_75t_L g5501 ( 
.A(n_5257),
.Y(n_5501)
);

BUFx10_ASAP7_75t_L g5502 ( 
.A(n_5264),
.Y(n_5502)
);

INVx3_ASAP7_75t_L g5503 ( 
.A(n_5247),
.Y(n_5503)
);

BUFx3_ASAP7_75t_L g5504 ( 
.A(n_5276),
.Y(n_5504)
);

OAI221xp5_ASAP7_75t_L g5505 ( 
.A1(n_5358),
.A2(n_5294),
.B1(n_5275),
.B2(n_5256),
.C(n_5353),
.Y(n_5505)
);

NAND2xp5_ASAP7_75t_L g5506 ( 
.A(n_5481),
.B(n_5199),
.Y(n_5506)
);

AND2x4_ASAP7_75t_L g5507 ( 
.A(n_5423),
.B(n_5278),
.Y(n_5507)
);

AOI21xp5_ASAP7_75t_L g5508 ( 
.A1(n_5366),
.A2(n_5203),
.B(n_5218),
.Y(n_5508)
);

BUFx2_ASAP7_75t_L g5509 ( 
.A(n_5409),
.Y(n_5509)
);

AND2x2_ASAP7_75t_L g5510 ( 
.A(n_5479),
.B(n_5295),
.Y(n_5510)
);

AOI22xp5_ASAP7_75t_L g5511 ( 
.A1(n_5363),
.A2(n_5252),
.B1(n_5212),
.B2(n_5258),
.Y(n_5511)
);

OA21x2_ASAP7_75t_L g5512 ( 
.A1(n_5428),
.A2(n_5299),
.B(n_5333),
.Y(n_5512)
);

NAND2xp5_ASAP7_75t_L g5513 ( 
.A(n_5439),
.B(n_5272),
.Y(n_5513)
);

NAND2xp5_ASAP7_75t_SL g5514 ( 
.A(n_5404),
.B(n_5249),
.Y(n_5514)
);

AOI22xp33_ASAP7_75t_SL g5515 ( 
.A1(n_5475),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_5515)
);

INVx2_ASAP7_75t_L g5516 ( 
.A(n_5400),
.Y(n_5516)
);

AOI21xp5_ASAP7_75t_L g5517 ( 
.A1(n_5375),
.A2(n_182),
.B(n_183),
.Y(n_5517)
);

OAI221xp5_ASAP7_75t_L g5518 ( 
.A1(n_5406),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.C(n_187),
.Y(n_5518)
);

OA21x2_ASAP7_75t_L g5519 ( 
.A1(n_5396),
.A2(n_184),
.B(n_185),
.Y(n_5519)
);

OAI22xp5_ASAP7_75t_L g5520 ( 
.A1(n_5361),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_5357),
.Y(n_5521)
);

INVx2_ASAP7_75t_L g5522 ( 
.A(n_5424),
.Y(n_5522)
);

BUFx2_ASAP7_75t_L g5523 ( 
.A(n_5437),
.Y(n_5523)
);

AO31x2_ASAP7_75t_L g5524 ( 
.A1(n_5501),
.A2(n_191),
.A3(n_189),
.B(n_190),
.Y(n_5524)
);

AOI21xp5_ASAP7_75t_L g5525 ( 
.A1(n_5490),
.A2(n_191),
.B(n_192),
.Y(n_5525)
);

BUFx6f_ASAP7_75t_SL g5526 ( 
.A(n_5381),
.Y(n_5526)
);

OAI22xp5_ASAP7_75t_L g5527 ( 
.A1(n_5447),
.A2(n_195),
.B1(n_192),
.B2(n_194),
.Y(n_5527)
);

OAI211xp5_ASAP7_75t_SL g5528 ( 
.A1(n_5391),
.A2(n_197),
.B(n_194),
.C(n_196),
.Y(n_5528)
);

OAI21xp5_ASAP7_75t_L g5529 ( 
.A1(n_5369),
.A2(n_197),
.B(n_198),
.Y(n_5529)
);

AOI21x1_ASAP7_75t_L g5530 ( 
.A1(n_5496),
.A2(n_198),
.B(n_199),
.Y(n_5530)
);

AND2x4_ASAP7_75t_L g5531 ( 
.A(n_5472),
.B(n_1867),
.Y(n_5531)
);

AOI22xp33_ASAP7_75t_L g5532 ( 
.A1(n_5359),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_5532)
);

AOI21x1_ASAP7_75t_L g5533 ( 
.A1(n_5495),
.A2(n_200),
.B(n_202),
.Y(n_5533)
);

INVx2_ASAP7_75t_L g5534 ( 
.A(n_5441),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_5362),
.Y(n_5535)
);

NAND2xp5_ASAP7_75t_L g5536 ( 
.A(n_5430),
.B(n_5417),
.Y(n_5536)
);

HB1xp67_ASAP7_75t_L g5537 ( 
.A(n_5368),
.Y(n_5537)
);

AOI21xp5_ASAP7_75t_L g5538 ( 
.A1(n_5416),
.A2(n_203),
.B(n_204),
.Y(n_5538)
);

OAI21xp5_ASAP7_75t_L g5539 ( 
.A1(n_5498),
.A2(n_204),
.B(n_205),
.Y(n_5539)
);

NAND2xp5_ASAP7_75t_L g5540 ( 
.A(n_5360),
.B(n_205),
.Y(n_5540)
);

BUFx3_ASAP7_75t_L g5541 ( 
.A(n_5484),
.Y(n_5541)
);

OAI21xp33_ASAP7_75t_L g5542 ( 
.A1(n_5476),
.A2(n_206),
.B(n_207),
.Y(n_5542)
);

OAI21x1_ASAP7_75t_L g5543 ( 
.A1(n_5503),
.A2(n_1869),
.B(n_1868),
.Y(n_5543)
);

OAI21xp33_ASAP7_75t_L g5544 ( 
.A1(n_5456),
.A2(n_206),
.B(n_207),
.Y(n_5544)
);

AOI22xp33_ASAP7_75t_L g5545 ( 
.A1(n_5389),
.A2(n_211),
.B1(n_208),
.B2(n_210),
.Y(n_5545)
);

AOI21xp5_ASAP7_75t_L g5546 ( 
.A1(n_5491),
.A2(n_210),
.B(n_211),
.Y(n_5546)
);

AND2x2_ASAP7_75t_L g5547 ( 
.A(n_5432),
.B(n_212),
.Y(n_5547)
);

OAI22xp5_ASAP7_75t_SL g5548 ( 
.A1(n_5465),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_5548)
);

AOI21xp5_ASAP7_75t_L g5549 ( 
.A1(n_5412),
.A2(n_213),
.B(n_214),
.Y(n_5549)
);

AO21x2_ASAP7_75t_L g5550 ( 
.A1(n_5422),
.A2(n_216),
.B(n_217),
.Y(n_5550)
);

NAND2xp5_ASAP7_75t_L g5551 ( 
.A(n_5384),
.B(n_216),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5370),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5376),
.Y(n_5553)
);

OAI221xp5_ASAP7_75t_L g5554 ( 
.A1(n_5377),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.C(n_220),
.Y(n_5554)
);

OA21x2_ASAP7_75t_L g5555 ( 
.A1(n_5387),
.A2(n_5394),
.B(n_5385),
.Y(n_5555)
);

A2O1A1Ixp33_ASAP7_75t_L g5556 ( 
.A1(n_5450),
.A2(n_221),
.B(n_218),
.C(n_220),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_5395),
.Y(n_5557)
);

AOI22xp33_ASAP7_75t_L g5558 ( 
.A1(n_5398),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_5558)
);

NAND2x1p5_ASAP7_75t_L g5559 ( 
.A(n_5454),
.B(n_5408),
.Y(n_5559)
);

OAI21xp5_ASAP7_75t_L g5560 ( 
.A1(n_5415),
.A2(n_224),
.B(n_225),
.Y(n_5560)
);

OAI22xp5_ASAP7_75t_L g5561 ( 
.A1(n_5418),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_5561)
);

INVx1_ASAP7_75t_L g5562 ( 
.A(n_5402),
.Y(n_5562)
);

AOI21xp5_ASAP7_75t_L g5563 ( 
.A1(n_5379),
.A2(n_226),
.B(n_228),
.Y(n_5563)
);

INVx2_ASAP7_75t_SL g5564 ( 
.A(n_5464),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_5405),
.Y(n_5565)
);

NAND2xp5_ASAP7_75t_L g5566 ( 
.A(n_5407),
.B(n_229),
.Y(n_5566)
);

OA21x2_ASAP7_75t_L g5567 ( 
.A1(n_5390),
.A2(n_5373),
.B(n_5426),
.Y(n_5567)
);

NAND2xp5_ASAP7_75t_L g5568 ( 
.A(n_5414),
.B(n_229),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_5420),
.Y(n_5569)
);

OAI22xp5_ASAP7_75t_L g5570 ( 
.A1(n_5485),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_5421),
.Y(n_5571)
);

INVx2_ASAP7_75t_L g5572 ( 
.A(n_5429),
.Y(n_5572)
);

CKINVDCx11_ASAP7_75t_R g5573 ( 
.A(n_5364),
.Y(n_5573)
);

OA21x2_ASAP7_75t_L g5574 ( 
.A1(n_5434),
.A2(n_231),
.B(n_232),
.Y(n_5574)
);

NAND2xp5_ASAP7_75t_L g5575 ( 
.A(n_5436),
.B(n_233),
.Y(n_5575)
);

AO31x2_ASAP7_75t_L g5576 ( 
.A1(n_5403),
.A2(n_235),
.A3(n_233),
.B(n_234),
.Y(n_5576)
);

OR2x2_ASAP7_75t_L g5577 ( 
.A(n_5457),
.B(n_235),
.Y(n_5577)
);

OA21x2_ASAP7_75t_L g5578 ( 
.A1(n_5419),
.A2(n_236),
.B(n_237),
.Y(n_5578)
);

HB1xp67_ASAP7_75t_L g5579 ( 
.A(n_5446),
.Y(n_5579)
);

OR2x2_ASAP7_75t_L g5580 ( 
.A(n_5458),
.B(n_237),
.Y(n_5580)
);

BUFx12f_ASAP7_75t_L g5581 ( 
.A(n_5411),
.Y(n_5581)
);

OAI22xp5_ASAP7_75t_L g5582 ( 
.A1(n_5386),
.A2(n_241),
.B1(n_238),
.B2(n_240),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5427),
.Y(n_5583)
);

AOI22xp33_ASAP7_75t_SL g5584 ( 
.A1(n_5443),
.A2(n_242),
.B1(n_238),
.B2(n_240),
.Y(n_5584)
);

AND2x2_ASAP7_75t_L g5585 ( 
.A(n_5425),
.B(n_242),
.Y(n_5585)
);

OA21x2_ASAP7_75t_L g5586 ( 
.A1(n_5469),
.A2(n_243),
.B(n_244),
.Y(n_5586)
);

OAI21x1_ASAP7_75t_L g5587 ( 
.A1(n_5438),
.A2(n_1872),
.B(n_1871),
.Y(n_5587)
);

INVx1_ASAP7_75t_L g5588 ( 
.A(n_5440),
.Y(n_5588)
);

OR2x2_ASAP7_75t_L g5589 ( 
.A(n_5461),
.B(n_243),
.Y(n_5589)
);

INVx2_ASAP7_75t_L g5590 ( 
.A(n_5473),
.Y(n_5590)
);

INVx2_ASAP7_75t_L g5591 ( 
.A(n_5504),
.Y(n_5591)
);

NAND2xp5_ASAP7_75t_L g5592 ( 
.A(n_5448),
.B(n_5451),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_5482),
.Y(n_5593)
);

AOI21xp5_ASAP7_75t_L g5594 ( 
.A1(n_5452),
.A2(n_244),
.B(n_245),
.Y(n_5594)
);

A2O1A1Ixp33_ASAP7_75t_L g5595 ( 
.A1(n_5480),
.A2(n_248),
.B(n_246),
.C(n_247),
.Y(n_5595)
);

AOI21xp5_ASAP7_75t_L g5596 ( 
.A1(n_5499),
.A2(n_247),
.B(n_248),
.Y(n_5596)
);

AOI21xp5_ASAP7_75t_L g5597 ( 
.A1(n_5410),
.A2(n_249),
.B(n_250),
.Y(n_5597)
);

INVx1_ASAP7_75t_SL g5598 ( 
.A(n_5433),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5459),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_5374),
.Y(n_5600)
);

NAND2xp5_ASAP7_75t_L g5601 ( 
.A(n_5413),
.B(n_250),
.Y(n_5601)
);

O2A1O1Ixp33_ASAP7_75t_L g5602 ( 
.A1(n_5442),
.A2(n_253),
.B(n_251),
.C(n_252),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_5371),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_5371),
.Y(n_5604)
);

CKINVDCx20_ASAP7_75t_R g5605 ( 
.A(n_5477),
.Y(n_5605)
);

OR2x2_ASAP7_75t_L g5606 ( 
.A(n_5431),
.B(n_251),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_5483),
.Y(n_5607)
);

HB1xp67_ASAP7_75t_L g5608 ( 
.A(n_5487),
.Y(n_5608)
);

AND2x4_ASAP7_75t_L g5609 ( 
.A(n_5500),
.B(n_1876),
.Y(n_5609)
);

AO31x2_ASAP7_75t_L g5610 ( 
.A1(n_5455),
.A2(n_255),
.A3(n_253),
.B(n_254),
.Y(n_5610)
);

INVx4_ASAP7_75t_L g5611 ( 
.A(n_5449),
.Y(n_5611)
);

INVx2_ASAP7_75t_L g5612 ( 
.A(n_5493),
.Y(n_5612)
);

NAND2xp5_ASAP7_75t_L g5613 ( 
.A(n_5478),
.B(n_254),
.Y(n_5613)
);

NAND2xp5_ASAP7_75t_L g5614 ( 
.A(n_5470),
.B(n_255),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_5392),
.Y(n_5615)
);

AOI22xp33_ASAP7_75t_L g5616 ( 
.A1(n_5444),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_5616)
);

BUFx2_ASAP7_75t_L g5617 ( 
.A(n_5392),
.Y(n_5617)
);

BUFx10_ASAP7_75t_L g5618 ( 
.A(n_5372),
.Y(n_5618)
);

INVx2_ASAP7_75t_L g5619 ( 
.A(n_5393),
.Y(n_5619)
);

OAI21x1_ASAP7_75t_L g5620 ( 
.A1(n_5471),
.A2(n_1879),
.B(n_1878),
.Y(n_5620)
);

INVx1_ASAP7_75t_L g5621 ( 
.A(n_5393),
.Y(n_5621)
);

AOI22xp33_ASAP7_75t_L g5622 ( 
.A1(n_5474),
.A2(n_261),
.B1(n_257),
.B2(n_260),
.Y(n_5622)
);

AOI22xp33_ASAP7_75t_L g5623 ( 
.A1(n_5486),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5502),
.Y(n_5624)
);

INVx1_ASAP7_75t_L g5625 ( 
.A(n_5464),
.Y(n_5625)
);

AOI21xp5_ASAP7_75t_L g5626 ( 
.A1(n_5462),
.A2(n_266),
.B(n_267),
.Y(n_5626)
);

OAI21xp5_ASAP7_75t_L g5627 ( 
.A1(n_5488),
.A2(n_267),
.B(n_268),
.Y(n_5627)
);

NAND2xp5_ASAP7_75t_L g5628 ( 
.A(n_5494),
.B(n_268),
.Y(n_5628)
);

NAND2xp5_ASAP7_75t_L g5629 ( 
.A(n_5489),
.B(n_269),
.Y(n_5629)
);

AOI21xp5_ASAP7_75t_L g5630 ( 
.A1(n_5460),
.A2(n_269),
.B(n_270),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_5489),
.Y(n_5631)
);

OA21x2_ASAP7_75t_L g5632 ( 
.A1(n_5463),
.A2(n_270),
.B(n_271),
.Y(n_5632)
);

AOI21xp5_ASAP7_75t_L g5633 ( 
.A1(n_5497),
.A2(n_271),
.B(n_273),
.Y(n_5633)
);

INVx2_ASAP7_75t_L g5634 ( 
.A(n_5401),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_5401),
.Y(n_5635)
);

OA21x2_ASAP7_75t_L g5636 ( 
.A1(n_5466),
.A2(n_274),
.B(n_275),
.Y(n_5636)
);

INVx1_ASAP7_75t_L g5637 ( 
.A(n_5492),
.Y(n_5637)
);

INVx4_ASAP7_75t_SL g5638 ( 
.A(n_5468),
.Y(n_5638)
);

AOI221xp5_ASAP7_75t_L g5639 ( 
.A1(n_5388),
.A2(n_5435),
.B1(n_5380),
.B2(n_5365),
.C(n_277),
.Y(n_5639)
);

AOI22xp33_ASAP7_75t_L g5640 ( 
.A1(n_5397),
.A2(n_277),
.B1(n_274),
.B2(n_276),
.Y(n_5640)
);

AND2x2_ASAP7_75t_L g5641 ( 
.A(n_5467),
.B(n_276),
.Y(n_5641)
);

OA21x2_ASAP7_75t_L g5642 ( 
.A1(n_5445),
.A2(n_278),
.B(n_279),
.Y(n_5642)
);

OAI21xp5_ASAP7_75t_L g5643 ( 
.A1(n_5367),
.A2(n_280),
.B(n_281),
.Y(n_5643)
);

INVx1_ASAP7_75t_L g5644 ( 
.A(n_5378),
.Y(n_5644)
);

INVx4_ASAP7_75t_L g5645 ( 
.A(n_5399),
.Y(n_5645)
);

NAND2xp5_ASAP7_75t_SL g5646 ( 
.A(n_5453),
.B(n_1880),
.Y(n_5646)
);

INVx2_ASAP7_75t_L g5647 ( 
.A(n_5378),
.Y(n_5647)
);

AOI21x1_ASAP7_75t_L g5648 ( 
.A1(n_5383),
.A2(n_282),
.B(n_283),
.Y(n_5648)
);

CKINVDCx20_ASAP7_75t_R g5649 ( 
.A(n_5382),
.Y(n_5649)
);

BUFx2_ASAP7_75t_L g5650 ( 
.A(n_5468),
.Y(n_5650)
);

NAND2xp5_ASAP7_75t_SL g5651 ( 
.A(n_5404),
.B(n_1881),
.Y(n_5651)
);

OAI22xp5_ASAP7_75t_L g5652 ( 
.A1(n_5358),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_5652)
);

AOI21xp5_ASAP7_75t_L g5653 ( 
.A1(n_5366),
.A2(n_285),
.B(n_286),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_5357),
.Y(n_5654)
);

OAI21x1_ASAP7_75t_L g5655 ( 
.A1(n_5503),
.A2(n_1883),
.B(n_1882),
.Y(n_5655)
);

BUFx3_ASAP7_75t_L g5656 ( 
.A(n_5484),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_5357),
.Y(n_5657)
);

AND3x2_ASAP7_75t_L g5658 ( 
.A(n_5495),
.B(n_286),
.C(n_287),
.Y(n_5658)
);

AND2x2_ASAP7_75t_L g5659 ( 
.A(n_5423),
.B(n_287),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_5357),
.Y(n_5660)
);

OAI21x1_ASAP7_75t_L g5661 ( 
.A1(n_5503),
.A2(n_1885),
.B(n_1884),
.Y(n_5661)
);

AOI22xp33_ASAP7_75t_L g5662 ( 
.A1(n_5358),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_5662)
);

A2O1A1Ixp33_ASAP7_75t_L g5663 ( 
.A1(n_5358),
.A2(n_290),
.B(n_288),
.C(n_289),
.Y(n_5663)
);

NAND2xp5_ASAP7_75t_L g5664 ( 
.A(n_5481),
.B(n_291),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5357),
.Y(n_5665)
);

AOI21xp5_ASAP7_75t_L g5666 ( 
.A1(n_5366),
.A2(n_292),
.B(n_293),
.Y(n_5666)
);

OAI21x1_ASAP7_75t_L g5667 ( 
.A1(n_5503),
.A2(n_1891),
.B(n_1886),
.Y(n_5667)
);

OAI22xp5_ASAP7_75t_L g5668 ( 
.A1(n_5545),
.A2(n_5529),
.B1(n_5554),
.B2(n_5518),
.Y(n_5668)
);

AOI22xp5_ASAP7_75t_L g5669 ( 
.A1(n_5528),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_5669)
);

AND2x2_ASAP7_75t_L g5670 ( 
.A(n_5509),
.B(n_5523),
.Y(n_5670)
);

AOI22xp5_ASAP7_75t_L g5671 ( 
.A1(n_5520),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_5671)
);

A2O1A1Ixp33_ASAP7_75t_L g5672 ( 
.A1(n_5653),
.A2(n_5666),
.B(n_5563),
.C(n_5517),
.Y(n_5672)
);

AOI21xp33_ASAP7_75t_L g5673 ( 
.A1(n_5511),
.A2(n_295),
.B(n_296),
.Y(n_5673)
);

AOI22xp33_ASAP7_75t_L g5674 ( 
.A1(n_5560),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_5674)
);

AOI21xp5_ASAP7_75t_L g5675 ( 
.A1(n_5508),
.A2(n_1893),
.B(n_1892),
.Y(n_5675)
);

INVx5_ASAP7_75t_SL g5676 ( 
.A(n_5573),
.Y(n_5676)
);

AOI21xp33_ASAP7_75t_L g5677 ( 
.A1(n_5514),
.A2(n_298),
.B(n_299),
.Y(n_5677)
);

AND2x4_ASAP7_75t_L g5678 ( 
.A(n_5507),
.B(n_300),
.Y(n_5678)
);

INVx3_ASAP7_75t_L g5679 ( 
.A(n_5619),
.Y(n_5679)
);

OAI221xp5_ASAP7_75t_L g5680 ( 
.A1(n_5539),
.A2(n_304),
.B1(n_300),
.B2(n_303),
.C(n_305),
.Y(n_5680)
);

OAI211xp5_ASAP7_75t_SL g5681 ( 
.A1(n_5663),
.A2(n_5639),
.B(n_5643),
.C(n_5662),
.Y(n_5681)
);

BUFx6f_ASAP7_75t_L g5682 ( 
.A(n_5581),
.Y(n_5682)
);

OAI22xp5_ASAP7_75t_L g5683 ( 
.A1(n_5556),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_5683)
);

AOI22xp5_ASAP7_75t_L g5684 ( 
.A1(n_5527),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_5684)
);

BUFx6f_ASAP7_75t_L g5685 ( 
.A(n_5541),
.Y(n_5685)
);

AOI221xp5_ASAP7_75t_L g5686 ( 
.A1(n_5652),
.A2(n_5602),
.B1(n_5548),
.B2(n_5544),
.C(n_5542),
.Y(n_5686)
);

NOR2xp33_ASAP7_75t_L g5687 ( 
.A(n_5650),
.B(n_307),
.Y(n_5687)
);

OAI21x1_ASAP7_75t_SL g5688 ( 
.A1(n_5530),
.A2(n_5648),
.B(n_5636),
.Y(n_5688)
);

OR2x2_ASAP7_75t_L g5689 ( 
.A(n_5537),
.B(n_308),
.Y(n_5689)
);

INVx1_ASAP7_75t_L g5690 ( 
.A(n_5521),
.Y(n_5690)
);

OAI221xp5_ASAP7_75t_L g5691 ( 
.A1(n_5532),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.C(n_313),
.Y(n_5691)
);

INVx2_ASAP7_75t_L g5692 ( 
.A(n_5535),
.Y(n_5692)
);

AOI22xp33_ASAP7_75t_L g5693 ( 
.A1(n_5593),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_5693)
);

AOI22xp33_ASAP7_75t_L g5694 ( 
.A1(n_5538),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_5552),
.Y(n_5695)
);

INVx2_ASAP7_75t_L g5696 ( 
.A(n_5553),
.Y(n_5696)
);

AOI22xp33_ASAP7_75t_L g5697 ( 
.A1(n_5651),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_5557),
.Y(n_5698)
);

OA21x2_ASAP7_75t_L g5699 ( 
.A1(n_5506),
.A2(n_316),
.B(n_317),
.Y(n_5699)
);

AOI22xp33_ASAP7_75t_L g5700 ( 
.A1(n_5627),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_5700)
);

AOI22xp33_ASAP7_75t_L g5701 ( 
.A1(n_5626),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_5701)
);

OA21x2_ASAP7_75t_L g5702 ( 
.A1(n_5600),
.A2(n_322),
.B(n_324),
.Y(n_5702)
);

AOI22xp33_ASAP7_75t_L g5703 ( 
.A1(n_5570),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_5703)
);

AOI221xp5_ASAP7_75t_L g5704 ( 
.A1(n_5628),
.A2(n_328),
.B1(n_325),
.B2(n_327),
.C(n_329),
.Y(n_5704)
);

INVx1_ASAP7_75t_L g5705 ( 
.A(n_5562),
.Y(n_5705)
);

BUFx6f_ASAP7_75t_L g5706 ( 
.A(n_5656),
.Y(n_5706)
);

INVx2_ASAP7_75t_L g5707 ( 
.A(n_5565),
.Y(n_5707)
);

AOI22xp33_ASAP7_75t_L g5708 ( 
.A1(n_5561),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_5708)
);

AOI22xp33_ASAP7_75t_L g5709 ( 
.A1(n_5582),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_5709)
);

AND2x4_ASAP7_75t_L g5710 ( 
.A(n_5603),
.B(n_331),
.Y(n_5710)
);

AND2x2_ASAP7_75t_L g5711 ( 
.A(n_5579),
.B(n_334),
.Y(n_5711)
);

AOI22xp33_ASAP7_75t_L g5712 ( 
.A1(n_5578),
.A2(n_338),
.B1(n_335),
.B2(n_337),
.Y(n_5712)
);

AOI222xp33_ASAP7_75t_L g5713 ( 
.A1(n_5613),
.A2(n_338),
.B1(n_340),
.B2(n_335),
.C1(n_337),
.C2(n_339),
.Y(n_5713)
);

AOI22xp33_ASAP7_75t_L g5714 ( 
.A1(n_5594),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_5714)
);

AOI22xp33_ASAP7_75t_SL g5715 ( 
.A1(n_5505),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.Y(n_5715)
);

AOI22xp33_ASAP7_75t_L g5716 ( 
.A1(n_5596),
.A2(n_345),
.B1(n_342),
.B2(n_343),
.Y(n_5716)
);

OAI22xp5_ASAP7_75t_L g5717 ( 
.A1(n_5595),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_5717)
);

AOI22xp33_ASAP7_75t_L g5718 ( 
.A1(n_5558),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_5718)
);

OAI221xp5_ASAP7_75t_L g5719 ( 
.A1(n_5515),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.C(n_351),
.Y(n_5719)
);

OAI221xp5_ASAP7_75t_L g5720 ( 
.A1(n_5633),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.C(n_352),
.Y(n_5720)
);

OAI211xp5_ASAP7_75t_SL g5721 ( 
.A1(n_5640),
.A2(n_354),
.B(n_352),
.C(n_353),
.Y(n_5721)
);

OAI221xp5_ASAP7_75t_L g5722 ( 
.A1(n_5584),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.C(n_356),
.Y(n_5722)
);

OAI22xp5_ASAP7_75t_SL g5723 ( 
.A1(n_5649),
.A2(n_358),
.B1(n_355),
.B2(n_357),
.Y(n_5723)
);

AOI221xp5_ASAP7_75t_L g5724 ( 
.A1(n_5614),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.C(n_360),
.Y(n_5724)
);

AND2x4_ASAP7_75t_L g5725 ( 
.A(n_5604),
.B(n_360),
.Y(n_5725)
);

AOI22xp33_ASAP7_75t_SL g5726 ( 
.A1(n_5586),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_5726)
);

BUFx2_ASAP7_75t_L g5727 ( 
.A(n_5559),
.Y(n_5727)
);

AOI22xp33_ASAP7_75t_L g5728 ( 
.A1(n_5630),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.Y(n_5728)
);

AOI22xp33_ASAP7_75t_L g5729 ( 
.A1(n_5632),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_5729)
);

INVx2_ASAP7_75t_L g5730 ( 
.A(n_5654),
.Y(n_5730)
);

OAI21x1_ASAP7_75t_L g5731 ( 
.A1(n_5513),
.A2(n_366),
.B(n_367),
.Y(n_5731)
);

AOI22xp33_ASAP7_75t_L g5732 ( 
.A1(n_5622),
.A2(n_5623),
.B1(n_5616),
.B2(n_5549),
.Y(n_5732)
);

AND2x2_ASAP7_75t_L g5733 ( 
.A(n_5617),
.B(n_367),
.Y(n_5733)
);

AOI22xp33_ASAP7_75t_L g5734 ( 
.A1(n_5525),
.A2(n_5546),
.B1(n_5597),
.B2(n_5510),
.Y(n_5734)
);

AOI22xp33_ASAP7_75t_L g5735 ( 
.A1(n_5550),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.Y(n_5735)
);

INVx3_ASAP7_75t_L g5736 ( 
.A(n_5647),
.Y(n_5736)
);

INVx2_ASAP7_75t_L g5737 ( 
.A(n_5657),
.Y(n_5737)
);

INVx1_ASAP7_75t_L g5738 ( 
.A(n_5660),
.Y(n_5738)
);

OR2x2_ASAP7_75t_L g5739 ( 
.A(n_5567),
.B(n_5536),
.Y(n_5739)
);

BUFx4f_ASAP7_75t_SL g5740 ( 
.A(n_5605),
.Y(n_5740)
);

AOI22xp33_ASAP7_75t_L g5741 ( 
.A1(n_5519),
.A2(n_372),
.B1(n_369),
.B2(n_370),
.Y(n_5741)
);

AOI221xp5_ASAP7_75t_SL g5742 ( 
.A1(n_5664),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.C(n_376),
.Y(n_5742)
);

OAI22xp5_ASAP7_75t_L g5743 ( 
.A1(n_5598),
.A2(n_377),
.B1(n_373),
.B2(n_376),
.Y(n_5743)
);

INVx2_ASAP7_75t_L g5744 ( 
.A(n_5665),
.Y(n_5744)
);

INVx1_ASAP7_75t_L g5745 ( 
.A(n_5534),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5572),
.Y(n_5746)
);

AOI22xp33_ASAP7_75t_L g5747 ( 
.A1(n_5620),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_5747)
);

AOI22xp33_ASAP7_75t_SL g5748 ( 
.A1(n_5642),
.A2(n_381),
.B1(n_378),
.B2(n_380),
.Y(n_5748)
);

OAI221xp5_ASAP7_75t_L g5749 ( 
.A1(n_5606),
.A2(n_5621),
.B1(n_5615),
.B2(n_5580),
.C(n_5592),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_5516),
.Y(n_5750)
);

NOR2x1_ASAP7_75t_R g5751 ( 
.A(n_5611),
.B(n_380),
.Y(n_5751)
);

INVx1_ASAP7_75t_SL g5752 ( 
.A(n_5644),
.Y(n_5752)
);

OAI21x1_ASAP7_75t_L g5753 ( 
.A1(n_5512),
.A2(n_381),
.B(n_382),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_5522),
.Y(n_5754)
);

AOI22xp33_ASAP7_75t_L g5755 ( 
.A1(n_5591),
.A2(n_5658),
.B1(n_5641),
.B2(n_5555),
.Y(n_5755)
);

AOI22xp33_ASAP7_75t_SL g5756 ( 
.A1(n_5574),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5569),
.Y(n_5757)
);

AND2x2_ASAP7_75t_L g5758 ( 
.A(n_5624),
.B(n_383),
.Y(n_5758)
);

OAI22xp5_ASAP7_75t_L g5759 ( 
.A1(n_5607),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_5759)
);

AND2x4_ASAP7_75t_L g5760 ( 
.A(n_5608),
.B(n_385),
.Y(n_5760)
);

CKINVDCx20_ASAP7_75t_R g5761 ( 
.A(n_5618),
.Y(n_5761)
);

AOI22xp33_ASAP7_75t_SL g5762 ( 
.A1(n_5659),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_5762)
);

A2O1A1Ixp33_ASAP7_75t_L g5763 ( 
.A1(n_5646),
.A2(n_5577),
.B(n_5655),
.C(n_5543),
.Y(n_5763)
);

HB1xp67_ASAP7_75t_L g5764 ( 
.A(n_5590),
.Y(n_5764)
);

OAI22xp5_ASAP7_75t_SL g5765 ( 
.A1(n_5645),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_5765)
);

AOI22xp33_ASAP7_75t_SL g5766 ( 
.A1(n_5531),
.A2(n_392),
.B1(n_389),
.B2(n_391),
.Y(n_5766)
);

CKINVDCx5p33_ASAP7_75t_R g5767 ( 
.A(n_5526),
.Y(n_5767)
);

INVx3_ASAP7_75t_L g5768 ( 
.A(n_5634),
.Y(n_5768)
);

BUFx3_ASAP7_75t_L g5769 ( 
.A(n_5564),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_5571),
.Y(n_5770)
);

AOI221xp5_ASAP7_75t_L g5771 ( 
.A1(n_5575),
.A2(n_5601),
.B1(n_5566),
.B2(n_5568),
.C(n_5551),
.Y(n_5771)
);

AOI22xp33_ASAP7_75t_L g5772 ( 
.A1(n_5599),
.A2(n_397),
.B1(n_393),
.B2(n_395),
.Y(n_5772)
);

AOI22xp33_ASAP7_75t_L g5773 ( 
.A1(n_5609),
.A2(n_399),
.B1(n_395),
.B2(n_398),
.Y(n_5773)
);

AOI22xp33_ASAP7_75t_L g5774 ( 
.A1(n_5625),
.A2(n_402),
.B1(n_399),
.B2(n_400),
.Y(n_5774)
);

AND2x2_ASAP7_75t_L g5775 ( 
.A(n_5588),
.B(n_400),
.Y(n_5775)
);

BUFx2_ASAP7_75t_L g5776 ( 
.A(n_5612),
.Y(n_5776)
);

AOI22xp33_ASAP7_75t_L g5777 ( 
.A1(n_5637),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_5777)
);

OR2x6_ASAP7_75t_L g5778 ( 
.A(n_5635),
.B(n_404),
.Y(n_5778)
);

AOI22xp33_ASAP7_75t_L g5779 ( 
.A1(n_5585),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_5779)
);

AOI22xp5_ASAP7_75t_L g5780 ( 
.A1(n_5631),
.A2(n_410),
.B1(n_406),
.B2(n_407),
.Y(n_5780)
);

AO31x2_ASAP7_75t_L g5781 ( 
.A1(n_5583),
.A2(n_413),
.A3(n_411),
.B(n_412),
.Y(n_5781)
);

INVx4_ASAP7_75t_L g5782 ( 
.A(n_5638),
.Y(n_5782)
);

BUFx6f_ASAP7_75t_L g5783 ( 
.A(n_5629),
.Y(n_5783)
);

OAI221xp5_ASAP7_75t_L g5784 ( 
.A1(n_5540),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.C(n_414),
.Y(n_5784)
);

OA21x2_ASAP7_75t_L g5785 ( 
.A1(n_5533),
.A2(n_415),
.B(n_416),
.Y(n_5785)
);

OAI21x1_ASAP7_75t_L g5786 ( 
.A1(n_5661),
.A2(n_416),
.B(n_417),
.Y(n_5786)
);

AND2x2_ASAP7_75t_SL g5787 ( 
.A(n_5589),
.B(n_419),
.Y(n_5787)
);

AND2x2_ASAP7_75t_L g5788 ( 
.A(n_5638),
.B(n_419),
.Y(n_5788)
);

OAI221xp5_ASAP7_75t_L g5789 ( 
.A1(n_5547),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.C(n_423),
.Y(n_5789)
);

AOI21xp33_ASAP7_75t_L g5790 ( 
.A1(n_5587),
.A2(n_420),
.B(n_421),
.Y(n_5790)
);

NOR2xp33_ASAP7_75t_L g5791 ( 
.A(n_5667),
.B(n_422),
.Y(n_5791)
);

OAI21x1_ASAP7_75t_L g5792 ( 
.A1(n_5524),
.A2(n_424),
.B(n_425),
.Y(n_5792)
);

OAI211xp5_ASAP7_75t_L g5793 ( 
.A1(n_5576),
.A2(n_426),
.B(n_424),
.C(n_425),
.Y(n_5793)
);

AND2x4_ASAP7_75t_L g5794 ( 
.A(n_5524),
.B(n_426),
.Y(n_5794)
);

AOI22xp33_ASAP7_75t_L g5795 ( 
.A1(n_5576),
.A2(n_430),
.B1(n_427),
.B2(n_428),
.Y(n_5795)
);

AOI221xp5_ASAP7_75t_L g5796 ( 
.A1(n_5610),
.A2(n_430),
.B1(n_427),
.B2(n_428),
.C(n_431),
.Y(n_5796)
);

INVx2_ASAP7_75t_L g5797 ( 
.A(n_5610),
.Y(n_5797)
);

HB1xp67_ASAP7_75t_L g5798 ( 
.A(n_5567),
.Y(n_5798)
);

OAI221xp5_ASAP7_75t_L g5799 ( 
.A1(n_5529),
.A2(n_434),
.B1(n_431),
.B2(n_433),
.C(n_435),
.Y(n_5799)
);

AND2x6_ASAP7_75t_L g5800 ( 
.A(n_5593),
.B(n_433),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5523),
.Y(n_5801)
);

AOI221xp5_ASAP7_75t_L g5802 ( 
.A1(n_5652),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.C(n_439),
.Y(n_5802)
);

INVxp67_ASAP7_75t_L g5803 ( 
.A(n_5579),
.Y(n_5803)
);

AOI22xp33_ASAP7_75t_L g5804 ( 
.A1(n_5529),
.A2(n_439),
.B1(n_436),
.B2(n_437),
.Y(n_5804)
);

AND2x2_ASAP7_75t_L g5805 ( 
.A(n_5509),
.B(n_441),
.Y(n_5805)
);

OR2x2_ASAP7_75t_L g5806 ( 
.A(n_5537),
.B(n_442),
.Y(n_5806)
);

OAI221xp5_ASAP7_75t_L g5807 ( 
.A1(n_5529),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.C(n_446),
.Y(n_5807)
);

OAI22xp5_ASAP7_75t_L g5808 ( 
.A1(n_5545),
.A2(n_448),
.B1(n_444),
.B2(n_447),
.Y(n_5808)
);

AOI22xp33_ASAP7_75t_L g5809 ( 
.A1(n_5529),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_5809)
);

AND2x4_ASAP7_75t_L g5810 ( 
.A(n_5507),
.B(n_449),
.Y(n_5810)
);

OAI33xp33_ASAP7_75t_L g5811 ( 
.A1(n_5652),
.A2(n_452),
.A3(n_454),
.B1(n_450),
.B2(n_451),
.B3(n_453),
.Y(n_5811)
);

INVx2_ASAP7_75t_L g5812 ( 
.A(n_5523),
.Y(n_5812)
);

BUFx2_ASAP7_75t_L g5813 ( 
.A(n_5559),
.Y(n_5813)
);

AOI31xp33_ASAP7_75t_SL g5814 ( 
.A1(n_5639),
.A2(n_453),
.A3(n_451),
.B(n_452),
.Y(n_5814)
);

AND2x2_ASAP7_75t_L g5815 ( 
.A(n_5509),
.B(n_455),
.Y(n_5815)
);

AOI21xp5_ASAP7_75t_L g5816 ( 
.A1(n_5508),
.A2(n_1895),
.B(n_1894),
.Y(n_5816)
);

OA21x2_ASAP7_75t_L g5817 ( 
.A1(n_5593),
.A2(n_456),
.B(n_457),
.Y(n_5817)
);

INVx1_ASAP7_75t_L g5818 ( 
.A(n_5521),
.Y(n_5818)
);

AOI22xp5_ASAP7_75t_L g5819 ( 
.A1(n_5528),
.A2(n_459),
.B1(n_457),
.B2(n_458),
.Y(n_5819)
);

AND2x2_ASAP7_75t_L g5820 ( 
.A(n_5509),
.B(n_458),
.Y(n_5820)
);

AOI21xp5_ASAP7_75t_L g5821 ( 
.A1(n_5508),
.A2(n_1898),
.B(n_1896),
.Y(n_5821)
);

AOI22xp33_ASAP7_75t_L g5822 ( 
.A1(n_5529),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_5822)
);

CKINVDCx20_ASAP7_75t_R g5823 ( 
.A(n_5605),
.Y(n_5823)
);

AOI221xp5_ASAP7_75t_L g5824 ( 
.A1(n_5652),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.C(n_465),
.Y(n_5824)
);

AOI21xp5_ASAP7_75t_L g5825 ( 
.A1(n_5508),
.A2(n_1902),
.B(n_1900),
.Y(n_5825)
);

INVx6_ASAP7_75t_L g5826 ( 
.A(n_5581),
.Y(n_5826)
);

OAI21x1_ASAP7_75t_L g5827 ( 
.A1(n_5508),
.A2(n_463),
.B(n_466),
.Y(n_5827)
);

NOR2xp33_ASAP7_75t_L g5828 ( 
.A(n_5650),
.B(n_467),
.Y(n_5828)
);

HB1xp67_ASAP7_75t_SL g5829 ( 
.A(n_5541),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5521),
.Y(n_5830)
);

AOI222xp33_ASAP7_75t_L g5831 ( 
.A1(n_5539),
.A2(n_471),
.B1(n_474),
.B2(n_467),
.C1(n_469),
.C2(n_472),
.Y(n_5831)
);

AOI221xp5_ASAP7_75t_L g5832 ( 
.A1(n_5652),
.A2(n_472),
.B1(n_469),
.B2(n_471),
.C(n_474),
.Y(n_5832)
);

AOI22xp5_ASAP7_75t_L g5833 ( 
.A1(n_5528),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.Y(n_5833)
);

AOI22xp33_ASAP7_75t_L g5834 ( 
.A1(n_5529),
.A2(n_480),
.B1(n_476),
.B2(n_479),
.Y(n_5834)
);

NAND2xp5_ASAP7_75t_L g5835 ( 
.A(n_5567),
.B(n_480),
.Y(n_5835)
);

BUFx6f_ASAP7_75t_L g5836 ( 
.A(n_5573),
.Y(n_5836)
);

AOI22xp33_ASAP7_75t_L g5837 ( 
.A1(n_5529),
.A2(n_484),
.B1(n_481),
.B2(n_483),
.Y(n_5837)
);

OAI21xp33_ASAP7_75t_SL g5838 ( 
.A1(n_5593),
.A2(n_481),
.B(n_484),
.Y(n_5838)
);

OAI22xp5_ASAP7_75t_L g5839 ( 
.A1(n_5545),
.A2(n_488),
.B1(n_485),
.B2(n_486),
.Y(n_5839)
);

OAI22xp5_ASAP7_75t_L g5840 ( 
.A1(n_5545),
.A2(n_489),
.B1(n_485),
.B2(n_486),
.Y(n_5840)
);

OAI22xp33_ASAP7_75t_SL g5841 ( 
.A1(n_5593),
.A2(n_493),
.B1(n_490),
.B2(n_491),
.Y(n_5841)
);

AOI22xp33_ASAP7_75t_L g5842 ( 
.A1(n_5529),
.A2(n_495),
.B1(n_491),
.B2(n_494),
.Y(n_5842)
);

AOI22xp33_ASAP7_75t_L g5843 ( 
.A1(n_5529),
.A2(n_497),
.B1(n_494),
.B2(n_496),
.Y(n_5843)
);

AOI22xp33_ASAP7_75t_L g5844 ( 
.A1(n_5529),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.Y(n_5844)
);

INVx2_ASAP7_75t_L g5845 ( 
.A(n_5523),
.Y(n_5845)
);

AOI22xp33_ASAP7_75t_L g5846 ( 
.A1(n_5529),
.A2(n_501),
.B1(n_498),
.B2(n_500),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_5521),
.Y(n_5847)
);

OAI22xp5_ASAP7_75t_L g5848 ( 
.A1(n_5545),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.Y(n_5848)
);

OAI22xp5_ASAP7_75t_L g5849 ( 
.A1(n_5545),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.Y(n_5849)
);

AOI221xp5_ASAP7_75t_SL g5850 ( 
.A1(n_5723),
.A2(n_509),
.B1(n_507),
.B2(n_508),
.C(n_511),
.Y(n_5850)
);

AND2x2_ASAP7_75t_L g5851 ( 
.A(n_5727),
.B(n_5813),
.Y(n_5851)
);

INVx2_ASAP7_75t_L g5852 ( 
.A(n_5692),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_5690),
.Y(n_5853)
);

INVx3_ASAP7_75t_L g5854 ( 
.A(n_5782),
.Y(n_5854)
);

INVx1_ASAP7_75t_L g5855 ( 
.A(n_5695),
.Y(n_5855)
);

AND2x2_ASAP7_75t_L g5856 ( 
.A(n_5670),
.B(n_509),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_5698),
.Y(n_5857)
);

AND2x2_ASAP7_75t_L g5858 ( 
.A(n_5801),
.B(n_511),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5705),
.Y(n_5859)
);

INVx2_ASAP7_75t_L g5860 ( 
.A(n_5696),
.Y(n_5860)
);

AOI21x1_ASAP7_75t_L g5861 ( 
.A1(n_5835),
.A2(n_512),
.B(n_513),
.Y(n_5861)
);

INVx1_ASAP7_75t_L g5862 ( 
.A(n_5738),
.Y(n_5862)
);

AOI222xp33_ASAP7_75t_L g5863 ( 
.A1(n_5686),
.A2(n_515),
.B1(n_517),
.B2(n_513),
.C1(n_514),
.C2(n_516),
.Y(n_5863)
);

BUFx2_ASAP7_75t_SL g5864 ( 
.A(n_5836),
.Y(n_5864)
);

AND2x2_ASAP7_75t_L g5865 ( 
.A(n_5812),
.B(n_514),
.Y(n_5865)
);

AOI211xp5_ASAP7_75t_L g5866 ( 
.A1(n_5814),
.A2(n_517),
.B(n_515),
.C(n_516),
.Y(n_5866)
);

NAND2xp5_ASAP7_75t_L g5867 ( 
.A(n_5803),
.B(n_518),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5818),
.Y(n_5868)
);

INVx1_ASAP7_75t_L g5869 ( 
.A(n_5830),
.Y(n_5869)
);

OR2x2_ASAP7_75t_L g5870 ( 
.A(n_5739),
.B(n_518),
.Y(n_5870)
);

AND2x2_ASAP7_75t_L g5871 ( 
.A(n_5845),
.B(n_519),
.Y(n_5871)
);

INVx2_ASAP7_75t_L g5872 ( 
.A(n_5707),
.Y(n_5872)
);

OR2x2_ASAP7_75t_L g5873 ( 
.A(n_5764),
.B(n_519),
.Y(n_5873)
);

AND2x2_ASAP7_75t_L g5874 ( 
.A(n_5679),
.B(n_520),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5847),
.Y(n_5875)
);

NOR2xp33_ASAP7_75t_L g5876 ( 
.A(n_5826),
.B(n_5836),
.Y(n_5876)
);

AND2x2_ASAP7_75t_L g5877 ( 
.A(n_5776),
.B(n_5736),
.Y(n_5877)
);

INVx2_ASAP7_75t_L g5878 ( 
.A(n_5730),
.Y(n_5878)
);

BUFx3_ASAP7_75t_L g5879 ( 
.A(n_5682),
.Y(n_5879)
);

AND2x2_ASAP7_75t_L g5880 ( 
.A(n_5752),
.B(n_520),
.Y(n_5880)
);

INVx1_ASAP7_75t_L g5881 ( 
.A(n_5737),
.Y(n_5881)
);

NAND2xp5_ASAP7_75t_L g5882 ( 
.A(n_5771),
.B(n_521),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_5744),
.Y(n_5883)
);

INVx2_ASAP7_75t_L g5884 ( 
.A(n_5757),
.Y(n_5884)
);

INVxp67_ASAP7_75t_L g5885 ( 
.A(n_5817),
.Y(n_5885)
);

AND2x4_ASAP7_75t_SL g5886 ( 
.A(n_5761),
.B(n_521),
.Y(n_5886)
);

INVx2_ASAP7_75t_L g5887 ( 
.A(n_5770),
.Y(n_5887)
);

INVx2_ASAP7_75t_L g5888 ( 
.A(n_5746),
.Y(n_5888)
);

NAND2xp5_ASAP7_75t_L g5889 ( 
.A(n_5750),
.B(n_5754),
.Y(n_5889)
);

INVx1_ASAP7_75t_L g5890 ( 
.A(n_5745),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_5798),
.Y(n_5891)
);

BUFx2_ASAP7_75t_L g5892 ( 
.A(n_5678),
.Y(n_5892)
);

INVxp67_ASAP7_75t_L g5893 ( 
.A(n_5749),
.Y(n_5893)
);

AND2x4_ASAP7_75t_L g5894 ( 
.A(n_5768),
.B(n_5769),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5797),
.Y(n_5895)
);

AND2x4_ASAP7_75t_L g5896 ( 
.A(n_5810),
.B(n_5783),
.Y(n_5896)
);

AND2x4_ASAP7_75t_L g5897 ( 
.A(n_5783),
.B(n_522),
.Y(n_5897)
);

BUFx2_ASAP7_75t_L g5898 ( 
.A(n_5826),
.Y(n_5898)
);

INVx5_ASAP7_75t_L g5899 ( 
.A(n_5676),
.Y(n_5899)
);

AO21x2_ASAP7_75t_L g5900 ( 
.A1(n_5688),
.A2(n_522),
.B(n_523),
.Y(n_5900)
);

AND2x2_ASAP7_75t_L g5901 ( 
.A(n_5676),
.B(n_5805),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5689),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5806),
.Y(n_5903)
);

AND2x2_ASAP7_75t_L g5904 ( 
.A(n_5815),
.B(n_524),
.Y(n_5904)
);

AND2x4_ASAP7_75t_L g5905 ( 
.A(n_5794),
.B(n_524),
.Y(n_5905)
);

BUFx2_ASAP7_75t_L g5906 ( 
.A(n_5800),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_5699),
.Y(n_5907)
);

AOI22xp33_ASAP7_75t_L g5908 ( 
.A1(n_5681),
.A2(n_528),
.B1(n_525),
.B2(n_527),
.Y(n_5908)
);

NAND2xp5_ASAP7_75t_L g5909 ( 
.A(n_5755),
.B(n_525),
.Y(n_5909)
);

INVx1_ASAP7_75t_L g5910 ( 
.A(n_5775),
.Y(n_5910)
);

AND2x4_ASAP7_75t_L g5911 ( 
.A(n_5763),
.B(n_528),
.Y(n_5911)
);

INVx3_ASAP7_75t_L g5912 ( 
.A(n_5682),
.Y(n_5912)
);

AND2x2_ASAP7_75t_L g5913 ( 
.A(n_5820),
.B(n_529),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_5753),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5711),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5702),
.Y(n_5916)
);

INVx4_ASAP7_75t_L g5917 ( 
.A(n_5767),
.Y(n_5917)
);

INVx1_ASAP7_75t_L g5918 ( 
.A(n_5781),
.Y(n_5918)
);

BUFx2_ASAP7_75t_L g5919 ( 
.A(n_5800),
.Y(n_5919)
);

INVx1_ASAP7_75t_L g5920 ( 
.A(n_5781),
.Y(n_5920)
);

AND2x2_ASAP7_75t_L g5921 ( 
.A(n_5733),
.B(n_529),
.Y(n_5921)
);

AND2x2_ASAP7_75t_L g5922 ( 
.A(n_5685),
.B(n_530),
.Y(n_5922)
);

AND2x4_ASAP7_75t_SL g5923 ( 
.A(n_5823),
.B(n_5685),
.Y(n_5923)
);

INVx2_ASAP7_75t_L g5924 ( 
.A(n_5792),
.Y(n_5924)
);

BUFx3_ASAP7_75t_L g5925 ( 
.A(n_5740),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5785),
.Y(n_5926)
);

NOR2xp33_ASAP7_75t_L g5927 ( 
.A(n_5829),
.B(n_530),
.Y(n_5927)
);

INVx2_ASAP7_75t_L g5928 ( 
.A(n_5731),
.Y(n_5928)
);

BUFx4f_ASAP7_75t_SL g5929 ( 
.A(n_5706),
.Y(n_5929)
);

INVx1_ASAP7_75t_L g5930 ( 
.A(n_5827),
.Y(n_5930)
);

NAND2xp5_ASAP7_75t_L g5931 ( 
.A(n_5734),
.B(n_531),
.Y(n_5931)
);

AND2x2_ASAP7_75t_L g5932 ( 
.A(n_5706),
.B(n_531),
.Y(n_5932)
);

AND2x2_ASAP7_75t_L g5933 ( 
.A(n_5758),
.B(n_532),
.Y(n_5933)
);

NAND3xp33_ASAP7_75t_L g5934 ( 
.A(n_5672),
.B(n_532),
.C(n_533),
.Y(n_5934)
);

HB1xp67_ASAP7_75t_L g5935 ( 
.A(n_5778),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5760),
.Y(n_5936)
);

INVx4_ASAP7_75t_L g5937 ( 
.A(n_5710),
.Y(n_5937)
);

AND2x2_ASAP7_75t_L g5938 ( 
.A(n_5787),
.B(n_533),
.Y(n_5938)
);

OR2x2_ASAP7_75t_L g5939 ( 
.A(n_5778),
.B(n_534),
.Y(n_5939)
);

INVx2_ASAP7_75t_L g5940 ( 
.A(n_5725),
.Y(n_5940)
);

NOR2x1_ASAP7_75t_L g5941 ( 
.A(n_5793),
.B(n_534),
.Y(n_5941)
);

OR2x2_ASAP7_75t_L g5942 ( 
.A(n_5687),
.B(n_535),
.Y(n_5942)
);

AND2x2_ASAP7_75t_L g5943 ( 
.A(n_5788),
.B(n_536),
.Y(n_5943)
);

INVx1_ASAP7_75t_L g5944 ( 
.A(n_5800),
.Y(n_5944)
);

AND2x2_ASAP7_75t_L g5945 ( 
.A(n_5828),
.B(n_536),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_5791),
.B(n_537),
.Y(n_5946)
);

OA21x2_ASAP7_75t_L g5947 ( 
.A1(n_5673),
.A2(n_537),
.B(n_538),
.Y(n_5947)
);

AND2x2_ASAP7_75t_L g5948 ( 
.A(n_5786),
.B(n_538),
.Y(n_5948)
);

INVx1_ASAP7_75t_L g5949 ( 
.A(n_5838),
.Y(n_5949)
);

HB1xp67_ASAP7_75t_L g5950 ( 
.A(n_5841),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5756),
.Y(n_5951)
);

NAND2xp5_ASAP7_75t_L g5952 ( 
.A(n_5742),
.B(n_539),
.Y(n_5952)
);

AND2x2_ASAP7_75t_L g5953 ( 
.A(n_5748),
.B(n_540),
.Y(n_5953)
);

BUFx3_ASAP7_75t_L g5954 ( 
.A(n_5765),
.Y(n_5954)
);

NAND2xp5_ASAP7_75t_L g5955 ( 
.A(n_5795),
.B(n_540),
.Y(n_5955)
);

INVx5_ASAP7_75t_L g5956 ( 
.A(n_5751),
.Y(n_5956)
);

INVx2_ASAP7_75t_L g5957 ( 
.A(n_5784),
.Y(n_5957)
);

AND2x2_ASAP7_75t_L g5958 ( 
.A(n_5741),
.B(n_541),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5780),
.Y(n_5959)
);

INVx2_ASAP7_75t_L g5960 ( 
.A(n_5789),
.Y(n_5960)
);

AND2x4_ASAP7_75t_L g5961 ( 
.A(n_5675),
.B(n_541),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5729),
.Y(n_5962)
);

NOR2x1_ASAP7_75t_SL g5963 ( 
.A(n_5743),
.B(n_542),
.Y(n_5963)
);

AND2x2_ASAP7_75t_L g5964 ( 
.A(n_5726),
.B(n_5790),
.Y(n_5964)
);

AND2x2_ASAP7_75t_L g5965 ( 
.A(n_5712),
.B(n_542),
.Y(n_5965)
);

NAND2xp5_ASAP7_75t_L g5966 ( 
.A(n_5677),
.B(n_543),
.Y(n_5966)
);

OR2x2_ASAP7_75t_L g5967 ( 
.A(n_5668),
.B(n_544),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5796),
.Y(n_5968)
);

AND2x2_ASAP7_75t_L g5969 ( 
.A(n_5747),
.B(n_544),
.Y(n_5969)
);

AND2x4_ASAP7_75t_SL g5970 ( 
.A(n_5779),
.B(n_545),
.Y(n_5970)
);

INVx2_ASAP7_75t_L g5971 ( 
.A(n_5720),
.Y(n_5971)
);

INVx2_ASAP7_75t_SL g5972 ( 
.A(n_5759),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5713),
.Y(n_5973)
);

AND2x4_ASAP7_75t_L g5974 ( 
.A(n_5816),
.B(n_546),
.Y(n_5974)
);

BUFx3_ASAP7_75t_L g5975 ( 
.A(n_5684),
.Y(n_5975)
);

AOI21xp5_ASAP7_75t_L g5976 ( 
.A1(n_5821),
.A2(n_546),
.B(n_547),
.Y(n_5976)
);

INVx2_ASAP7_75t_L g5977 ( 
.A(n_5680),
.Y(n_5977)
);

OR2x2_ASAP7_75t_L g5978 ( 
.A(n_5735),
.B(n_547),
.Y(n_5978)
);

INVx2_ASAP7_75t_L g5979 ( 
.A(n_5799),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5669),
.Y(n_5980)
);

AO21x2_ASAP7_75t_L g5981 ( 
.A1(n_5825),
.A2(n_548),
.B(n_549),
.Y(n_5981)
);

OR2x2_ASAP7_75t_L g5982 ( 
.A(n_5693),
.B(n_549),
.Y(n_5982)
);

AND2x4_ASAP7_75t_L g5983 ( 
.A(n_5819),
.B(n_550),
.Y(n_5983)
);

OAI321xp33_ASAP7_75t_L g5984 ( 
.A1(n_5807),
.A2(n_552),
.A3(n_554),
.B1(n_550),
.B2(n_551),
.C(n_553),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_5833),
.Y(n_5985)
);

INVx5_ASAP7_75t_L g5986 ( 
.A(n_5762),
.Y(n_5986)
);

OR2x2_ASAP7_75t_L g5987 ( 
.A(n_5732),
.B(n_551),
.Y(n_5987)
);

INVx2_ASAP7_75t_L g5988 ( 
.A(n_5719),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5683),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5717),
.Y(n_5990)
);

INVx1_ASAP7_75t_L g5991 ( 
.A(n_5831),
.Y(n_5991)
);

HB1xp67_ASAP7_75t_L g5992 ( 
.A(n_5704),
.Y(n_5992)
);

INVx3_ASAP7_75t_L g5993 ( 
.A(n_5766),
.Y(n_5993)
);

INVx1_ASAP7_75t_L g5994 ( 
.A(n_5724),
.Y(n_5994)
);

INVx2_ASAP7_75t_L g5995 ( 
.A(n_5671),
.Y(n_5995)
);

NAND2xp5_ASAP7_75t_L g5996 ( 
.A(n_5715),
.B(n_552),
.Y(n_5996)
);

BUFx3_ASAP7_75t_L g5997 ( 
.A(n_5722),
.Y(n_5997)
);

AND2x2_ASAP7_75t_L g5998 ( 
.A(n_5694),
.B(n_553),
.Y(n_5998)
);

INVxp67_ASAP7_75t_L g5999 ( 
.A(n_5811),
.Y(n_5999)
);

BUFx3_ASAP7_75t_L g6000 ( 
.A(n_5691),
.Y(n_6000)
);

INVx2_ASAP7_75t_L g6001 ( 
.A(n_5808),
.Y(n_6001)
);

AND2x2_ASAP7_75t_L g6002 ( 
.A(n_5773),
.B(n_555),
.Y(n_6002)
);

INVx2_ASAP7_75t_L g6003 ( 
.A(n_5839),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5728),
.Y(n_6004)
);

NAND2xp5_ASAP7_75t_L g6005 ( 
.A(n_5674),
.B(n_556),
.Y(n_6005)
);

INVx1_ASAP7_75t_L g6006 ( 
.A(n_5840),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5848),
.Y(n_6007)
);

INVx5_ASAP7_75t_L g6008 ( 
.A(n_5802),
.Y(n_6008)
);

HB1xp67_ASAP7_75t_L g6009 ( 
.A(n_5849),
.Y(n_6009)
);

AND2x2_ASAP7_75t_L g6010 ( 
.A(n_5714),
.B(n_556),
.Y(n_6010)
);

OR2x6_ASAP7_75t_L g6011 ( 
.A(n_5804),
.B(n_557),
.Y(n_6011)
);

AND2x2_ASAP7_75t_L g6012 ( 
.A(n_5716),
.B(n_557),
.Y(n_6012)
);

INVx1_ASAP7_75t_L g6013 ( 
.A(n_5774),
.Y(n_6013)
);

NAND2xp5_ASAP7_75t_L g6014 ( 
.A(n_5809),
.B(n_558),
.Y(n_6014)
);

NOR4xp25_ASAP7_75t_SL g6015 ( 
.A(n_5721),
.B(n_562),
.C(n_559),
.D(n_561),
.Y(n_6015)
);

INVxp67_ASAP7_75t_SL g6016 ( 
.A(n_5701),
.Y(n_6016)
);

INVxp67_ASAP7_75t_L g6017 ( 
.A(n_5824),
.Y(n_6017)
);

AND2x2_ASAP7_75t_L g6018 ( 
.A(n_5772),
.B(n_561),
.Y(n_6018)
);

AND2x2_ASAP7_75t_L g6019 ( 
.A(n_5697),
.B(n_562),
.Y(n_6019)
);

INVx2_ASAP7_75t_L g6020 ( 
.A(n_5832),
.Y(n_6020)
);

OAI222xp33_ASAP7_75t_L g6021 ( 
.A1(n_5822),
.A2(n_567),
.B1(n_569),
.B2(n_563),
.C1(n_566),
.C2(n_568),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_5700),
.Y(n_6022)
);

BUFx3_ASAP7_75t_L g6023 ( 
.A(n_5777),
.Y(n_6023)
);

INVx2_ASAP7_75t_SL g6024 ( 
.A(n_5834),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5837),
.Y(n_6025)
);

INVx1_ASAP7_75t_L g6026 ( 
.A(n_5842),
.Y(n_6026)
);

HB1xp67_ASAP7_75t_L g6027 ( 
.A(n_5843),
.Y(n_6027)
);

AND2x2_ASAP7_75t_L g6028 ( 
.A(n_5844),
.B(n_563),
.Y(n_6028)
);

OR2x2_ASAP7_75t_L g6029 ( 
.A(n_5846),
.B(n_567),
.Y(n_6029)
);

INVx2_ASAP7_75t_L g6030 ( 
.A(n_5708),
.Y(n_6030)
);

AND2x2_ASAP7_75t_L g6031 ( 
.A(n_5703),
.B(n_568),
.Y(n_6031)
);

INVx1_ASAP7_75t_L g6032 ( 
.A(n_5709),
.Y(n_6032)
);

INVx2_ASAP7_75t_L g6033 ( 
.A(n_5718),
.Y(n_6033)
);

INVx1_ASAP7_75t_L g6034 ( 
.A(n_5690),
.Y(n_6034)
);

AND2x2_ASAP7_75t_L g6035 ( 
.A(n_5727),
.B(n_570),
.Y(n_6035)
);

INVx2_ASAP7_75t_L g6036 ( 
.A(n_5692),
.Y(n_6036)
);

NAND2xp5_ASAP7_75t_L g6037 ( 
.A(n_5803),
.B(n_571),
.Y(n_6037)
);

AND2x2_ASAP7_75t_L g6038 ( 
.A(n_5727),
.B(n_571),
.Y(n_6038)
);

AND2x2_ASAP7_75t_L g6039 ( 
.A(n_5727),
.B(n_573),
.Y(n_6039)
);

AND2x2_ASAP7_75t_L g6040 ( 
.A(n_5727),
.B(n_573),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5690),
.Y(n_6041)
);

AND2x2_ASAP7_75t_L g6042 ( 
.A(n_5727),
.B(n_574),
.Y(n_6042)
);

CKINVDCx6p67_ASAP7_75t_R g6043 ( 
.A(n_5836),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5690),
.Y(n_6044)
);

AND2x2_ASAP7_75t_L g6045 ( 
.A(n_5727),
.B(n_574),
.Y(n_6045)
);

AND2x2_ASAP7_75t_L g6046 ( 
.A(n_5727),
.B(n_575),
.Y(n_6046)
);

INVx2_ASAP7_75t_L g6047 ( 
.A(n_5692),
.Y(n_6047)
);

INVx1_ASAP7_75t_L g6048 ( 
.A(n_5690),
.Y(n_6048)
);

NAND2xp5_ASAP7_75t_L g6049 ( 
.A(n_5803),
.B(n_575),
.Y(n_6049)
);

INVx2_ASAP7_75t_L g6050 ( 
.A(n_5692),
.Y(n_6050)
);

INVx1_ASAP7_75t_L g6051 ( 
.A(n_5690),
.Y(n_6051)
);

AND2x2_ASAP7_75t_L g6052 ( 
.A(n_5727),
.B(n_576),
.Y(n_6052)
);

AOI22xp33_ASAP7_75t_L g6053 ( 
.A1(n_5681),
.A2(n_579),
.B1(n_576),
.B2(n_577),
.Y(n_6053)
);

AOI21xp5_ASAP7_75t_L g6054 ( 
.A1(n_5934),
.A2(n_577),
.B(n_579),
.Y(n_6054)
);

AO31x2_ASAP7_75t_L g6055 ( 
.A1(n_5916),
.A2(n_582),
.A3(n_580),
.B(n_581),
.Y(n_6055)
);

AOI211xp5_ASAP7_75t_L g6056 ( 
.A1(n_5992),
.A2(n_583),
.B(n_580),
.C(n_581),
.Y(n_6056)
);

NAND2xp5_ASAP7_75t_L g6057 ( 
.A(n_5893),
.B(n_583),
.Y(n_6057)
);

HB1xp67_ASAP7_75t_L g6058 ( 
.A(n_5891),
.Y(n_6058)
);

OAI22xp5_ASAP7_75t_L g6059 ( 
.A1(n_5986),
.A2(n_586),
.B1(n_584),
.B2(n_585),
.Y(n_6059)
);

INVx2_ASAP7_75t_L g6060 ( 
.A(n_5851),
.Y(n_6060)
);

AND2x4_ASAP7_75t_L g6061 ( 
.A(n_5898),
.B(n_584),
.Y(n_6061)
);

BUFx2_ASAP7_75t_L g6062 ( 
.A(n_5906),
.Y(n_6062)
);

BUFx3_ASAP7_75t_L g6063 ( 
.A(n_5899),
.Y(n_6063)
);

NAND4xp25_ASAP7_75t_L g6064 ( 
.A(n_5866),
.B(n_588),
.C(n_585),
.D(n_587),
.Y(n_6064)
);

INVx2_ASAP7_75t_L g6065 ( 
.A(n_5944),
.Y(n_6065)
);

AOI22xp33_ASAP7_75t_L g6066 ( 
.A1(n_6008),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_6066)
);

INVx1_ASAP7_75t_L g6067 ( 
.A(n_5853),
.Y(n_6067)
);

INVx2_ASAP7_75t_L g6068 ( 
.A(n_5852),
.Y(n_6068)
);

INVx1_ASAP7_75t_L g6069 ( 
.A(n_5855),
.Y(n_6069)
);

AOI21xp33_ASAP7_75t_L g6070 ( 
.A1(n_5991),
.A2(n_589),
.B(n_590),
.Y(n_6070)
);

AOI221xp5_ASAP7_75t_L g6071 ( 
.A1(n_6017),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.C(n_593),
.Y(n_6071)
);

AOI22xp33_ASAP7_75t_SL g6072 ( 
.A1(n_5986),
.A2(n_594),
.B1(n_591),
.B2(n_593),
.Y(n_6072)
);

HB1xp67_ASAP7_75t_L g6073 ( 
.A(n_5907),
.Y(n_6073)
);

AND2x2_ASAP7_75t_L g6074 ( 
.A(n_5877),
.B(n_595),
.Y(n_6074)
);

NAND2xp5_ASAP7_75t_L g6075 ( 
.A(n_5928),
.B(n_595),
.Y(n_6075)
);

NOR3xp33_ASAP7_75t_L g6076 ( 
.A(n_5973),
.B(n_596),
.C(n_597),
.Y(n_6076)
);

INVx1_ASAP7_75t_L g6077 ( 
.A(n_5857),
.Y(n_6077)
);

INVx2_ASAP7_75t_SL g6078 ( 
.A(n_5899),
.Y(n_6078)
);

AND2x2_ASAP7_75t_L g6079 ( 
.A(n_5919),
.B(n_596),
.Y(n_6079)
);

INVx2_ASAP7_75t_L g6080 ( 
.A(n_5860),
.Y(n_6080)
);

AOI22xp33_ASAP7_75t_L g6081 ( 
.A1(n_6008),
.A2(n_600),
.B1(n_597),
.B2(n_599),
.Y(n_6081)
);

OA21x2_ASAP7_75t_L g6082 ( 
.A1(n_5885),
.A2(n_599),
.B(n_601),
.Y(n_6082)
);

NOR2xp33_ASAP7_75t_L g6083 ( 
.A(n_6043),
.B(n_601),
.Y(n_6083)
);

INVx2_ASAP7_75t_L g6084 ( 
.A(n_5872),
.Y(n_6084)
);

NOR2xp33_ASAP7_75t_L g6085 ( 
.A(n_5876),
.B(n_602),
.Y(n_6085)
);

NAND2xp5_ASAP7_75t_L g6086 ( 
.A(n_5870),
.B(n_602),
.Y(n_6086)
);

INVx2_ASAP7_75t_L g6087 ( 
.A(n_5878),
.Y(n_6087)
);

AOI22xp33_ASAP7_75t_L g6088 ( 
.A1(n_6000),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.Y(n_6088)
);

OAI21x1_ASAP7_75t_L g6089 ( 
.A1(n_5895),
.A2(n_5924),
.B(n_5914),
.Y(n_6089)
);

INVx2_ASAP7_75t_L g6090 ( 
.A(n_6036),
.Y(n_6090)
);

OAI21x1_ASAP7_75t_L g6091 ( 
.A1(n_5918),
.A2(n_5920),
.B(n_5926),
.Y(n_6091)
);

AND2x2_ASAP7_75t_L g6092 ( 
.A(n_5894),
.B(n_604),
.Y(n_6092)
);

AOI21xp33_ASAP7_75t_L g6093 ( 
.A1(n_6016),
.A2(n_605),
.B(n_606),
.Y(n_6093)
);

NAND4xp25_ASAP7_75t_L g6094 ( 
.A(n_5863),
.B(n_612),
.C(n_607),
.D(n_609),
.Y(n_6094)
);

OAI211xp5_ASAP7_75t_L g6095 ( 
.A1(n_5950),
.A2(n_612),
.B(n_607),
.C(n_609),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_5859),
.Y(n_6096)
);

AOI22xp33_ASAP7_75t_L g6097 ( 
.A1(n_5997),
.A2(n_616),
.B1(n_614),
.B2(n_615),
.Y(n_6097)
);

AOI21xp5_ASAP7_75t_L g6098 ( 
.A1(n_5941),
.A2(n_617),
.B(n_618),
.Y(n_6098)
);

INVx1_ASAP7_75t_L g6099 ( 
.A(n_5862),
.Y(n_6099)
);

OAI21xp33_ASAP7_75t_L g6100 ( 
.A1(n_5908),
.A2(n_617),
.B(n_619),
.Y(n_6100)
);

OAI22xp33_ASAP7_75t_L g6101 ( 
.A1(n_5968),
.A2(n_623),
.B1(n_620),
.B2(n_621),
.Y(n_6101)
);

INVx2_ASAP7_75t_L g6102 ( 
.A(n_6047),
.Y(n_6102)
);

AND2x4_ASAP7_75t_L g6103 ( 
.A(n_5854),
.B(n_620),
.Y(n_6103)
);

HB1xp67_ASAP7_75t_L g6104 ( 
.A(n_5930),
.Y(n_6104)
);

OAI22xp5_ASAP7_75t_L g6105 ( 
.A1(n_5990),
.A2(n_5985),
.B1(n_5980),
.B2(n_5999),
.Y(n_6105)
);

AND2x2_ASAP7_75t_L g6106 ( 
.A(n_5935),
.B(n_621),
.Y(n_6106)
);

INVx2_ASAP7_75t_SL g6107 ( 
.A(n_5879),
.Y(n_6107)
);

NOR2xp33_ASAP7_75t_L g6108 ( 
.A(n_5917),
.B(n_624),
.Y(n_6108)
);

OAI21x1_ASAP7_75t_L g6109 ( 
.A1(n_5888),
.A2(n_625),
.B(n_626),
.Y(n_6109)
);

INVx2_ASAP7_75t_L g6110 ( 
.A(n_6050),
.Y(n_6110)
);

OR2x2_ASAP7_75t_L g6111 ( 
.A(n_5902),
.B(n_625),
.Y(n_6111)
);

INVxp67_ASAP7_75t_R g6112 ( 
.A(n_5901),
.Y(n_6112)
);

AOI21xp5_ASAP7_75t_L g6113 ( 
.A1(n_5931),
.A2(n_626),
.B(n_627),
.Y(n_6113)
);

HB1xp67_ASAP7_75t_L g6114 ( 
.A(n_5949),
.Y(n_6114)
);

INVx1_ASAP7_75t_L g6115 ( 
.A(n_5868),
.Y(n_6115)
);

A2O1A1Ixp33_ASAP7_75t_L g6116 ( 
.A1(n_5911),
.A2(n_630),
.B(n_628),
.C(n_629),
.Y(n_6116)
);

INVx2_ASAP7_75t_L g6117 ( 
.A(n_5884),
.Y(n_6117)
);

AOI22xp33_ASAP7_75t_SL g6118 ( 
.A1(n_6027),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.Y(n_6118)
);

INVx2_ASAP7_75t_L g6119 ( 
.A(n_5887),
.Y(n_6119)
);

OAI22xp33_ASAP7_75t_L g6120 ( 
.A1(n_5957),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.Y(n_6120)
);

AO21x2_ASAP7_75t_L g6121 ( 
.A1(n_5909),
.A2(n_634),
.B(n_635),
.Y(n_6121)
);

INVx2_ASAP7_75t_L g6122 ( 
.A(n_5881),
.Y(n_6122)
);

NOR2xp33_ASAP7_75t_R g6123 ( 
.A(n_5956),
.B(n_636),
.Y(n_6123)
);

AOI221xp5_ASAP7_75t_L g6124 ( 
.A1(n_5994),
.A2(n_639),
.B1(n_635),
.B2(n_638),
.C(n_640),
.Y(n_6124)
);

INVx2_ASAP7_75t_L g6125 ( 
.A(n_5883),
.Y(n_6125)
);

NOR2xp33_ASAP7_75t_SL g6126 ( 
.A(n_5956),
.B(n_638),
.Y(n_6126)
);

INVx1_ASAP7_75t_L g6127 ( 
.A(n_5869),
.Y(n_6127)
);

HB1xp67_ASAP7_75t_L g6128 ( 
.A(n_5890),
.Y(n_6128)
);

OR2x2_ASAP7_75t_L g6129 ( 
.A(n_5903),
.B(n_5915),
.Y(n_6129)
);

BUFx5_ASAP7_75t_L g6130 ( 
.A(n_5897),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_5875),
.Y(n_6131)
);

INVx2_ASAP7_75t_L g6132 ( 
.A(n_6034),
.Y(n_6132)
);

AND2x2_ASAP7_75t_L g6133 ( 
.A(n_5892),
.B(n_639),
.Y(n_6133)
);

AND2x2_ASAP7_75t_L g6134 ( 
.A(n_5910),
.B(n_641),
.Y(n_6134)
);

AND4x1_ASAP7_75t_L g6135 ( 
.A(n_6053),
.B(n_645),
.C(n_641),
.D(n_642),
.Y(n_6135)
);

INVx1_ASAP7_75t_L g6136 ( 
.A(n_6041),
.Y(n_6136)
);

AND2x4_ASAP7_75t_L g6137 ( 
.A(n_5896),
.B(n_642),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_6044),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_6048),
.Y(n_6139)
);

AOI21xp5_ASAP7_75t_L g6140 ( 
.A1(n_5984),
.A2(n_645),
.B(n_646),
.Y(n_6140)
);

AO31x2_ASAP7_75t_L g6141 ( 
.A1(n_5882),
.A2(n_648),
.A3(n_646),
.B(n_647),
.Y(n_6141)
);

AND2x2_ASAP7_75t_L g6142 ( 
.A(n_5936),
.B(n_647),
.Y(n_6142)
);

INVxp67_ASAP7_75t_L g6143 ( 
.A(n_5971),
.Y(n_6143)
);

A2O1A1Ixp33_ASAP7_75t_L g6144 ( 
.A1(n_5977),
.A2(n_650),
.B(n_648),
.C(n_649),
.Y(n_6144)
);

AOI221x1_ASAP7_75t_SL g6145 ( 
.A1(n_5951),
.A2(n_651),
.B1(n_649),
.B2(n_650),
.C(n_652),
.Y(n_6145)
);

OR2x2_ASAP7_75t_L g6146 ( 
.A(n_5889),
.B(n_652),
.Y(n_6146)
);

OR2x2_ASAP7_75t_L g6147 ( 
.A(n_5873),
.B(n_653),
.Y(n_6147)
);

AOI22xp33_ASAP7_75t_L g6148 ( 
.A1(n_5979),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.Y(n_6148)
);

INVx2_ASAP7_75t_L g6149 ( 
.A(n_6051),
.Y(n_6149)
);

OA21x2_ASAP7_75t_L g6150 ( 
.A1(n_5867),
.A2(n_6049),
.B(n_6037),
.Y(n_6150)
);

AOI22xp33_ASAP7_75t_L g6151 ( 
.A1(n_6023),
.A2(n_656),
.B1(n_654),
.B2(n_655),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_5861),
.Y(n_6152)
);

OAI211xp5_ASAP7_75t_L g6153 ( 
.A1(n_5850),
.A2(n_658),
.B(n_656),
.C(n_657),
.Y(n_6153)
);

INVx2_ASAP7_75t_L g6154 ( 
.A(n_5940),
.Y(n_6154)
);

AOI21xp5_ASAP7_75t_L g6155 ( 
.A1(n_5952),
.A2(n_657),
.B(n_658),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_5858),
.Y(n_6156)
);

INVx1_ASAP7_75t_L g6157 ( 
.A(n_5865),
.Y(n_6157)
);

INVx2_ASAP7_75t_L g6158 ( 
.A(n_5905),
.Y(n_6158)
);

INVx2_ASAP7_75t_L g6159 ( 
.A(n_5937),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_5871),
.Y(n_6160)
);

AOI21xp5_ASAP7_75t_L g6161 ( 
.A1(n_5976),
.A2(n_659),
.B(n_660),
.Y(n_6161)
);

OA21x2_ASAP7_75t_L g6162 ( 
.A1(n_6035),
.A2(n_659),
.B(n_660),
.Y(n_6162)
);

INVx2_ASAP7_75t_L g6163 ( 
.A(n_5874),
.Y(n_6163)
);

INVx1_ASAP7_75t_L g6164 ( 
.A(n_5900),
.Y(n_6164)
);

INVx1_ASAP7_75t_L g6165 ( 
.A(n_5880),
.Y(n_6165)
);

INVxp67_ASAP7_75t_L g6166 ( 
.A(n_6009),
.Y(n_6166)
);

INVx1_ASAP7_75t_L g6167 ( 
.A(n_5948),
.Y(n_6167)
);

OAI21x1_ASAP7_75t_L g6168 ( 
.A1(n_6038),
.A2(n_661),
.B(n_662),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_6052),
.Y(n_6169)
);

AO21x2_ASAP7_75t_L g6170 ( 
.A1(n_6039),
.A2(n_661),
.B(n_664),
.Y(n_6170)
);

NAND3xp33_ASAP7_75t_L g6171 ( 
.A(n_6020),
.B(n_665),
.C(n_666),
.Y(n_6171)
);

INVx1_ASAP7_75t_L g6172 ( 
.A(n_6040),
.Y(n_6172)
);

AO21x2_ASAP7_75t_L g6173 ( 
.A1(n_6042),
.A2(n_667),
.B(n_668),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_6045),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_6046),
.Y(n_6175)
);

OAI22xp33_ASAP7_75t_L g6176 ( 
.A1(n_5993),
.A2(n_669),
.B1(n_667),
.B2(n_668),
.Y(n_6176)
);

INVx1_ASAP7_75t_SL g6177 ( 
.A(n_5864),
.Y(n_6177)
);

OR2x2_ASAP7_75t_L g6178 ( 
.A(n_5995),
.B(n_5989),
.Y(n_6178)
);

NAND2xp5_ASAP7_75t_L g6179 ( 
.A(n_5959),
.B(n_671),
.Y(n_6179)
);

INVx4_ASAP7_75t_SL g6180 ( 
.A(n_5929),
.Y(n_6180)
);

NAND2xp5_ASAP7_75t_L g6181 ( 
.A(n_5960),
.B(n_671),
.Y(n_6181)
);

OA21x2_ASAP7_75t_L g6182 ( 
.A1(n_5856),
.A2(n_672),
.B(n_673),
.Y(n_6182)
);

OA21x2_ASAP7_75t_L g6183 ( 
.A1(n_6006),
.A2(n_673),
.B(n_674),
.Y(n_6183)
);

BUFx6f_ASAP7_75t_L g6184 ( 
.A(n_5912),
.Y(n_6184)
);

INVx1_ASAP7_75t_L g6185 ( 
.A(n_6007),
.Y(n_6185)
);

INVx2_ASAP7_75t_L g6186 ( 
.A(n_5972),
.Y(n_6186)
);

OA21x2_ASAP7_75t_L g6187 ( 
.A1(n_5962),
.A2(n_674),
.B(n_675),
.Y(n_6187)
);

INVx1_ASAP7_75t_L g6188 ( 
.A(n_6001),
.Y(n_6188)
);

AOI21xp5_ASAP7_75t_L g6189 ( 
.A1(n_5955),
.A2(n_675),
.B(n_677),
.Y(n_6189)
);

OAI22xp33_ASAP7_75t_L g6190 ( 
.A1(n_5954),
.A2(n_680),
.B1(n_678),
.B2(n_679),
.Y(n_6190)
);

OAI211xp5_ASAP7_75t_L g6191 ( 
.A1(n_5996),
.A2(n_680),
.B(n_678),
.C(n_679),
.Y(n_6191)
);

A2O1A1Ixp33_ASAP7_75t_L g6192 ( 
.A1(n_5988),
.A2(n_683),
.B(n_681),
.C(n_682),
.Y(n_6192)
);

AND2x4_ASAP7_75t_L g6193 ( 
.A(n_5923),
.B(n_681),
.Y(n_6193)
);

INVx2_ASAP7_75t_L g6194 ( 
.A(n_5975),
.Y(n_6194)
);

INVxp67_ASAP7_75t_SL g6195 ( 
.A(n_5927),
.Y(n_6195)
);

OA21x2_ASAP7_75t_L g6196 ( 
.A1(n_6003),
.A2(n_683),
.B(n_684),
.Y(n_6196)
);

INVx1_ASAP7_75t_L g6197 ( 
.A(n_6004),
.Y(n_6197)
);

NAND2xp5_ASAP7_75t_L g6198 ( 
.A(n_5946),
.B(n_684),
.Y(n_6198)
);

AND2x4_ASAP7_75t_L g6199 ( 
.A(n_5925),
.B(n_685),
.Y(n_6199)
);

OR2x2_ASAP7_75t_L g6200 ( 
.A(n_6030),
.B(n_686),
.Y(n_6200)
);

INVx1_ASAP7_75t_L g6201 ( 
.A(n_6032),
.Y(n_6201)
);

INVx1_ASAP7_75t_L g6202 ( 
.A(n_6025),
.Y(n_6202)
);

AOI22xp33_ASAP7_75t_L g6203 ( 
.A1(n_5983),
.A2(n_6024),
.B1(n_5964),
.B2(n_6022),
.Y(n_6203)
);

NAND2xp5_ASAP7_75t_SL g6204 ( 
.A(n_5961),
.B(n_687),
.Y(n_6204)
);

INVx4_ASAP7_75t_SL g6205 ( 
.A(n_5938),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_6026),
.Y(n_6206)
);

OA21x2_ASAP7_75t_L g6207 ( 
.A1(n_5967),
.A2(n_687),
.B(n_689),
.Y(n_6207)
);

OAI21xp5_ASAP7_75t_L g6208 ( 
.A1(n_5987),
.A2(n_689),
.B(n_690),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_6033),
.Y(n_6209)
);

AOI211xp5_ASAP7_75t_L g6210 ( 
.A1(n_6021),
.A2(n_693),
.B(n_691),
.C(n_692),
.Y(n_6210)
);

INVx1_ASAP7_75t_L g6211 ( 
.A(n_6013),
.Y(n_6211)
);

OR2x2_ASAP7_75t_L g6212 ( 
.A(n_5942),
.B(n_692),
.Y(n_6212)
);

HB1xp67_ASAP7_75t_L g6213 ( 
.A(n_5939),
.Y(n_6213)
);

NAND2xp5_ASAP7_75t_L g6214 ( 
.A(n_5904),
.B(n_5913),
.Y(n_6214)
);

OA21x2_ASAP7_75t_L g6215 ( 
.A1(n_5943),
.A2(n_693),
.B(n_694),
.Y(n_6215)
);

OAI21x1_ASAP7_75t_L g6216 ( 
.A1(n_5921),
.A2(n_695),
.B(n_696),
.Y(n_6216)
);

AND2x2_ASAP7_75t_L g6217 ( 
.A(n_5933),
.B(n_695),
.Y(n_6217)
);

OAI22xp5_ASAP7_75t_L g6218 ( 
.A1(n_6011),
.A2(n_699),
.B1(n_697),
.B2(n_698),
.Y(n_6218)
);

OAI21xp5_ASAP7_75t_L g6219 ( 
.A1(n_5966),
.A2(n_697),
.B(n_699),
.Y(n_6219)
);

AND2x2_ASAP7_75t_L g6220 ( 
.A(n_5922),
.B(n_700),
.Y(n_6220)
);

INVx1_ASAP7_75t_L g6221 ( 
.A(n_5947),
.Y(n_6221)
);

INVx1_ASAP7_75t_L g6222 ( 
.A(n_5932),
.Y(n_6222)
);

INVx2_ASAP7_75t_L g6223 ( 
.A(n_5981),
.Y(n_6223)
);

NOR2xp33_ASAP7_75t_L g6224 ( 
.A(n_5945),
.B(n_700),
.Y(n_6224)
);

INVx1_ASAP7_75t_L g6225 ( 
.A(n_5963),
.Y(n_6225)
);

AOI21xp5_ASAP7_75t_L g6226 ( 
.A1(n_6005),
.A2(n_701),
.B(n_702),
.Y(n_6226)
);

OR2x2_ASAP7_75t_L g6227 ( 
.A(n_5978),
.B(n_704),
.Y(n_6227)
);

NOR2xp33_ASAP7_75t_L g6228 ( 
.A(n_5886),
.B(n_704),
.Y(n_6228)
);

NAND2xp5_ASAP7_75t_L g6229 ( 
.A(n_5953),
.B(n_705),
.Y(n_6229)
);

INVx2_ASAP7_75t_L g6230 ( 
.A(n_5974),
.Y(n_6230)
);

OAI22xp33_ASAP7_75t_L g6231 ( 
.A1(n_6011),
.A2(n_707),
.B1(n_705),
.B2(n_706),
.Y(n_6231)
);

INVx1_ASAP7_75t_L g6232 ( 
.A(n_6029),
.Y(n_6232)
);

AND2x2_ASAP7_75t_L g6233 ( 
.A(n_6002),
.B(n_706),
.Y(n_6233)
);

NAND4xp25_ASAP7_75t_L g6234 ( 
.A(n_6014),
.B(n_710),
.C(n_708),
.D(n_709),
.Y(n_6234)
);

INVx1_ASAP7_75t_L g6235 ( 
.A(n_5958),
.Y(n_6235)
);

NOR2x1_ASAP7_75t_L g6236 ( 
.A(n_5982),
.B(n_708),
.Y(n_6236)
);

AND2x2_ASAP7_75t_L g6237 ( 
.A(n_5965),
.B(n_709),
.Y(n_6237)
);

HB1xp67_ASAP7_75t_L g6238 ( 
.A(n_5969),
.Y(n_6238)
);

INVxp67_ASAP7_75t_L g6239 ( 
.A(n_6019),
.Y(n_6239)
);

BUFx6f_ASAP7_75t_L g6240 ( 
.A(n_6031),
.Y(n_6240)
);

AND2x2_ASAP7_75t_L g6241 ( 
.A(n_5970),
.B(n_711),
.Y(n_6241)
);

INVxp67_ASAP7_75t_SL g6242 ( 
.A(n_6018),
.Y(n_6242)
);

HB1xp67_ASAP7_75t_L g6243 ( 
.A(n_5998),
.Y(n_6243)
);

AO21x2_ASAP7_75t_L g6244 ( 
.A1(n_6028),
.A2(n_712),
.B(n_713),
.Y(n_6244)
);

BUFx2_ASAP7_75t_L g6245 ( 
.A(n_6010),
.Y(n_6245)
);

AND2x4_ASAP7_75t_SL g6246 ( 
.A(n_6012),
.B(n_712),
.Y(n_6246)
);

OAI21xp5_ASAP7_75t_L g6247 ( 
.A1(n_6015),
.A2(n_713),
.B(n_714),
.Y(n_6247)
);

OA21x2_ASAP7_75t_L g6248 ( 
.A1(n_5885),
.A2(n_715),
.B(n_716),
.Y(n_6248)
);

OA21x2_ASAP7_75t_L g6249 ( 
.A1(n_5885),
.A2(n_715),
.B(n_716),
.Y(n_6249)
);

INVx1_ASAP7_75t_L g6250 ( 
.A(n_5853),
.Y(n_6250)
);

INVx2_ASAP7_75t_L g6251 ( 
.A(n_5851),
.Y(n_6251)
);

INVxp67_ASAP7_75t_L g6252 ( 
.A(n_5935),
.Y(n_6252)
);

HB1xp67_ASAP7_75t_L g6253 ( 
.A(n_5891),
.Y(n_6253)
);

INVx2_ASAP7_75t_SL g6254 ( 
.A(n_5899),
.Y(n_6254)
);

INVx2_ASAP7_75t_L g6255 ( 
.A(n_5851),
.Y(n_6255)
);

OAI22xp5_ASAP7_75t_L g6256 ( 
.A1(n_5986),
.A2(n_719),
.B1(n_717),
.B2(n_718),
.Y(n_6256)
);

INVx3_ASAP7_75t_L g6257 ( 
.A(n_5879),
.Y(n_6257)
);

OR2x2_ASAP7_75t_L g6258 ( 
.A(n_5907),
.B(n_717),
.Y(n_6258)
);

AOI22xp33_ASAP7_75t_L g6259 ( 
.A1(n_6008),
.A2(n_721),
.B1(n_718),
.B2(n_720),
.Y(n_6259)
);

INVx1_ASAP7_75t_L g6260 ( 
.A(n_5853),
.Y(n_6260)
);

INVx2_ASAP7_75t_L g6261 ( 
.A(n_5851),
.Y(n_6261)
);

AO21x2_ASAP7_75t_L g6262 ( 
.A1(n_5891),
.A2(n_720),
.B(n_721),
.Y(n_6262)
);

INVx2_ASAP7_75t_L g6263 ( 
.A(n_5851),
.Y(n_6263)
);

INVx1_ASAP7_75t_L g6264 ( 
.A(n_5853),
.Y(n_6264)
);

AND2x2_ASAP7_75t_L g6265 ( 
.A(n_5851),
.B(n_722),
.Y(n_6265)
);

INVx3_ASAP7_75t_L g6266 ( 
.A(n_5879),
.Y(n_6266)
);

OAI22xp5_ASAP7_75t_L g6267 ( 
.A1(n_5986),
.A2(n_725),
.B1(n_723),
.B2(n_724),
.Y(n_6267)
);

AOI22xp33_ASAP7_75t_L g6268 ( 
.A1(n_6008),
.A2(n_726),
.B1(n_723),
.B2(n_725),
.Y(n_6268)
);

AND2x2_ASAP7_75t_L g6269 ( 
.A(n_5851),
.B(n_726),
.Y(n_6269)
);

NAND2xp5_ASAP7_75t_L g6270 ( 
.A(n_5893),
.B(n_728),
.Y(n_6270)
);

OAI21xp5_ASAP7_75t_SL g6271 ( 
.A1(n_5934),
.A2(n_728),
.B(n_729),
.Y(n_6271)
);

HB1xp67_ASAP7_75t_L g6272 ( 
.A(n_5891),
.Y(n_6272)
);

AOI22xp33_ASAP7_75t_L g6273 ( 
.A1(n_6008),
.A2(n_731),
.B1(n_729),
.B2(n_730),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_5853),
.Y(n_6274)
);

INVx2_ASAP7_75t_L g6275 ( 
.A(n_5851),
.Y(n_6275)
);

AND2x2_ASAP7_75t_L g6276 ( 
.A(n_5851),
.B(n_730),
.Y(n_6276)
);

AOI22xp5_ASAP7_75t_L g6277 ( 
.A1(n_6008),
.A2(n_733),
.B1(n_731),
.B2(n_732),
.Y(n_6277)
);

AO31x2_ASAP7_75t_L g6278 ( 
.A1(n_5916),
.A2(n_735),
.A3(n_732),
.B(n_734),
.Y(n_6278)
);

AOI21xp5_ASAP7_75t_L g6279 ( 
.A1(n_5934),
.A2(n_734),
.B(n_735),
.Y(n_6279)
);

NAND2xp5_ASAP7_75t_L g6280 ( 
.A(n_5893),
.B(n_736),
.Y(n_6280)
);

HB1xp67_ASAP7_75t_L g6281 ( 
.A(n_5891),
.Y(n_6281)
);

INVx2_ASAP7_75t_L g6282 ( 
.A(n_5851),
.Y(n_6282)
);

AOI22xp33_ASAP7_75t_L g6283 ( 
.A1(n_6008),
.A2(n_738),
.B1(n_736),
.B2(n_737),
.Y(n_6283)
);

OAI21xp5_ASAP7_75t_L g6284 ( 
.A1(n_5934),
.A2(n_738),
.B(n_739),
.Y(n_6284)
);

BUFx8_ASAP7_75t_L g6285 ( 
.A(n_5922),
.Y(n_6285)
);

AOI22xp33_ASAP7_75t_L g6286 ( 
.A1(n_6008),
.A2(n_741),
.B1(n_739),
.B2(n_740),
.Y(n_6286)
);

OAI21x1_ASAP7_75t_L g6287 ( 
.A1(n_5891),
.A2(n_740),
.B(n_741),
.Y(n_6287)
);

INVx2_ASAP7_75t_L g6288 ( 
.A(n_5851),
.Y(n_6288)
);

OA21x2_ASAP7_75t_L g6289 ( 
.A1(n_5885),
.A2(n_744),
.B(n_745),
.Y(n_6289)
);

NOR3xp33_ASAP7_75t_L g6290 ( 
.A(n_5934),
.B(n_744),
.C(n_745),
.Y(n_6290)
);

NAND3xp33_ASAP7_75t_L g6291 ( 
.A(n_6008),
.B(n_746),
.C(n_747),
.Y(n_6291)
);

INVx6_ASAP7_75t_L g6292 ( 
.A(n_5899),
.Y(n_6292)
);

OAI21xp33_ASAP7_75t_L g6293 ( 
.A1(n_6000),
.A2(n_746),
.B(n_748),
.Y(n_6293)
);

INVx1_ASAP7_75t_SL g6294 ( 
.A(n_5864),
.Y(n_6294)
);

INVx2_ASAP7_75t_L g6295 ( 
.A(n_5851),
.Y(n_6295)
);

HB1xp67_ASAP7_75t_L g6296 ( 
.A(n_5891),
.Y(n_6296)
);

O2A1O1Ixp33_ASAP7_75t_L g6297 ( 
.A1(n_5950),
.A2(n_751),
.B(n_752),
.C(n_750),
.Y(n_6297)
);

INVxp67_ASAP7_75t_L g6298 ( 
.A(n_5935),
.Y(n_6298)
);

BUFx2_ASAP7_75t_L g6299 ( 
.A(n_5898),
.Y(n_6299)
);

AOI21xp5_ASAP7_75t_L g6300 ( 
.A1(n_5934),
.A2(n_749),
.B(n_750),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_5853),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_5853),
.Y(n_6302)
);

NAND2xp5_ASAP7_75t_L g6303 ( 
.A(n_5893),
.B(n_749),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_5853),
.Y(n_6304)
);

BUFx8_ASAP7_75t_L g6305 ( 
.A(n_5922),
.Y(n_6305)
);

INVx5_ASAP7_75t_SL g6306 ( 
.A(n_6043),
.Y(n_6306)
);

NAND2xp5_ASAP7_75t_L g6307 ( 
.A(n_5893),
.B(n_751),
.Y(n_6307)
);

INVx1_ASAP7_75t_L g6308 ( 
.A(n_5853),
.Y(n_6308)
);

INVx2_ASAP7_75t_L g6309 ( 
.A(n_5851),
.Y(n_6309)
);

INVxp67_ASAP7_75t_L g6310 ( 
.A(n_5935),
.Y(n_6310)
);

AOI21xp5_ASAP7_75t_L g6311 ( 
.A1(n_5934),
.A2(n_753),
.B(n_755),
.Y(n_6311)
);

OA21x2_ASAP7_75t_L g6312 ( 
.A1(n_5885),
.A2(n_753),
.B(n_756),
.Y(n_6312)
);

NAND2xp5_ASAP7_75t_L g6313 ( 
.A(n_5893),
.B(n_756),
.Y(n_6313)
);

OAI221xp5_ASAP7_75t_L g6314 ( 
.A1(n_6072),
.A2(n_6145),
.B1(n_6277),
.B2(n_6076),
.C(n_6271),
.Y(n_6314)
);

INVx2_ASAP7_75t_L g6315 ( 
.A(n_6299),
.Y(n_6315)
);

OAI22xp5_ASAP7_75t_L g6316 ( 
.A1(n_6166),
.A2(n_759),
.B1(n_757),
.B2(n_758),
.Y(n_6316)
);

AND2x2_ASAP7_75t_L g6317 ( 
.A(n_6112),
.B(n_758),
.Y(n_6317)
);

AOI221xp5_ASAP7_75t_L g6318 ( 
.A1(n_6059),
.A2(n_6267),
.B1(n_6256),
.B2(n_6297),
.C(n_6105),
.Y(n_6318)
);

AOI221xp5_ASAP7_75t_L g6319 ( 
.A1(n_6291),
.A2(n_761),
.B1(n_759),
.B2(n_760),
.C(n_762),
.Y(n_6319)
);

BUFx3_ASAP7_75t_L g6320 ( 
.A(n_6292),
.Y(n_6320)
);

AND2x2_ASAP7_75t_L g6321 ( 
.A(n_6062),
.B(n_760),
.Y(n_6321)
);

OAI31xp33_ASAP7_75t_SL g6322 ( 
.A1(n_6153),
.A2(n_763),
.A3(n_764),
.B(n_762),
.Y(n_6322)
);

INVx2_ASAP7_75t_L g6323 ( 
.A(n_6078),
.Y(n_6323)
);

BUFx6f_ASAP7_75t_L g6324 ( 
.A(n_6063),
.Y(n_6324)
);

OR2x2_ASAP7_75t_L g6325 ( 
.A(n_6252),
.B(n_6310),
.Y(n_6325)
);

BUFx3_ASAP7_75t_L g6326 ( 
.A(n_6292),
.Y(n_6326)
);

AND2x2_ASAP7_75t_L g6327 ( 
.A(n_6186),
.B(n_761),
.Y(n_6327)
);

AO21x2_ASAP7_75t_L g6328 ( 
.A1(n_6164),
.A2(n_763),
.B(n_765),
.Y(n_6328)
);

AOI221xp5_ASAP7_75t_L g6329 ( 
.A1(n_6070),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.C(n_769),
.Y(n_6329)
);

HB1xp67_ASAP7_75t_L g6330 ( 
.A(n_6114),
.Y(n_6330)
);

AND2x2_ASAP7_75t_L g6331 ( 
.A(n_6194),
.B(n_766),
.Y(n_6331)
);

INVx1_ASAP7_75t_L g6332 ( 
.A(n_6128),
.Y(n_6332)
);

AND2x2_ASAP7_75t_L g6333 ( 
.A(n_6159),
.B(n_767),
.Y(n_6333)
);

INVxp33_ASAP7_75t_L g6334 ( 
.A(n_6123),
.Y(n_6334)
);

INVxp67_ASAP7_75t_L g6335 ( 
.A(n_6195),
.Y(n_6335)
);

INVx2_ASAP7_75t_L g6336 ( 
.A(n_6254),
.Y(n_6336)
);

AND2x4_ASAP7_75t_L g6337 ( 
.A(n_6177),
.B(n_768),
.Y(n_6337)
);

INVx2_ASAP7_75t_L g6338 ( 
.A(n_6130),
.Y(n_6338)
);

NAND2xp5_ASAP7_75t_L g6339 ( 
.A(n_6143),
.B(n_770),
.Y(n_6339)
);

INVxp67_ASAP7_75t_SL g6340 ( 
.A(n_6225),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_6067),
.Y(n_6341)
);

BUFx3_ASAP7_75t_L g6342 ( 
.A(n_6285),
.Y(n_6342)
);

INVx2_ASAP7_75t_L g6343 ( 
.A(n_6130),
.Y(n_6343)
);

AND2x2_ASAP7_75t_L g6344 ( 
.A(n_6060),
.B(n_770),
.Y(n_6344)
);

OAI221xp5_ASAP7_75t_L g6345 ( 
.A1(n_6203),
.A2(n_773),
.B1(n_771),
.B2(n_772),
.C(n_775),
.Y(n_6345)
);

OAI33xp33_ASAP7_75t_L g6346 ( 
.A1(n_6221),
.A2(n_775),
.A3(n_777),
.B1(n_771),
.B2(n_772),
.B3(n_776),
.Y(n_6346)
);

INVx1_ASAP7_75t_L g6347 ( 
.A(n_6069),
.Y(n_6347)
);

CKINVDCx5p33_ASAP7_75t_R g6348 ( 
.A(n_6305),
.Y(n_6348)
);

HB1xp67_ASAP7_75t_L g6349 ( 
.A(n_6073),
.Y(n_6349)
);

BUFx2_ASAP7_75t_L g6350 ( 
.A(n_6205),
.Y(n_6350)
);

NAND2xp5_ASAP7_75t_L g6351 ( 
.A(n_6298),
.B(n_6213),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_6077),
.Y(n_6352)
);

NOR2xp33_ASAP7_75t_L g6353 ( 
.A(n_6294),
.B(n_776),
.Y(n_6353)
);

INVx3_ASAP7_75t_L g6354 ( 
.A(n_6306),
.Y(n_6354)
);

AND2x2_ASAP7_75t_L g6355 ( 
.A(n_6251),
.B(n_778),
.Y(n_6355)
);

OAI22xp5_ASAP7_75t_L g6356 ( 
.A1(n_6210),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_6356)
);

NOR2x1_ASAP7_75t_L g6357 ( 
.A(n_6262),
.B(n_779),
.Y(n_6357)
);

CKINVDCx5p33_ASAP7_75t_R g6358 ( 
.A(n_6180),
.Y(n_6358)
);

INVx2_ASAP7_75t_L g6359 ( 
.A(n_6130),
.Y(n_6359)
);

INVx2_ASAP7_75t_L g6360 ( 
.A(n_6130),
.Y(n_6360)
);

OAI31xp33_ASAP7_75t_SL g6361 ( 
.A1(n_6236),
.A2(n_783),
.A3(n_784),
.B(n_781),
.Y(n_6361)
);

INVx2_ASAP7_75t_L g6362 ( 
.A(n_6257),
.Y(n_6362)
);

INVx3_ASAP7_75t_L g6363 ( 
.A(n_6306),
.Y(n_6363)
);

NAND2xp5_ASAP7_75t_L g6364 ( 
.A(n_6197),
.B(n_6201),
.Y(n_6364)
);

OA222x2_ASAP7_75t_L g6365 ( 
.A1(n_6223),
.A2(n_784),
.B1(n_787),
.B2(n_780),
.C1(n_783),
.C2(n_785),
.Y(n_6365)
);

OAI321xp33_ASAP7_75t_L g6366 ( 
.A1(n_6094),
.A2(n_788),
.A3(n_790),
.B1(n_785),
.B2(n_787),
.C(n_789),
.Y(n_6366)
);

AND2x4_ASAP7_75t_L g6367 ( 
.A(n_6266),
.B(n_788),
.Y(n_6367)
);

INVxp67_ASAP7_75t_SL g6368 ( 
.A(n_6238),
.Y(n_6368)
);

OR2x2_ASAP7_75t_L g6369 ( 
.A(n_6209),
.B(n_791),
.Y(n_6369)
);

AND2x4_ASAP7_75t_L g6370 ( 
.A(n_6107),
.B(n_791),
.Y(n_6370)
);

NAND2xp5_ASAP7_75t_L g6371 ( 
.A(n_6202),
.B(n_792),
.Y(n_6371)
);

NAND2xp5_ASAP7_75t_L g6372 ( 
.A(n_6206),
.B(n_792),
.Y(n_6372)
);

INVxp67_ASAP7_75t_L g6373 ( 
.A(n_6126),
.Y(n_6373)
);

INVx2_ASAP7_75t_L g6374 ( 
.A(n_6184),
.Y(n_6374)
);

AOI22xp5_ASAP7_75t_L g6375 ( 
.A1(n_6290),
.A2(n_795),
.B1(n_793),
.B2(n_794),
.Y(n_6375)
);

INVx1_ASAP7_75t_L g6376 ( 
.A(n_6096),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_6099),
.Y(n_6377)
);

AO21x2_ASAP7_75t_L g6378 ( 
.A1(n_6091),
.A2(n_6270),
.B(n_6057),
.Y(n_6378)
);

INVx2_ASAP7_75t_L g6379 ( 
.A(n_6184),
.Y(n_6379)
);

INVx2_ASAP7_75t_L g6380 ( 
.A(n_6230),
.Y(n_6380)
);

AND2x2_ASAP7_75t_L g6381 ( 
.A(n_6255),
.B(n_793),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_6115),
.Y(n_6382)
);

INVx2_ASAP7_75t_L g6383 ( 
.A(n_6261),
.Y(n_6383)
);

INVxp67_ASAP7_75t_SL g6384 ( 
.A(n_6243),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_6127),
.Y(n_6385)
);

NAND2xp5_ASAP7_75t_L g6386 ( 
.A(n_6211),
.B(n_794),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_6131),
.Y(n_6387)
);

NAND2x1_ASAP7_75t_L g6388 ( 
.A(n_6263),
.B(n_796),
.Y(n_6388)
);

AND2x2_ASAP7_75t_L g6389 ( 
.A(n_6275),
.B(n_796),
.Y(n_6389)
);

INVx1_ASAP7_75t_L g6390 ( 
.A(n_6136),
.Y(n_6390)
);

AND2x2_ASAP7_75t_L g6391 ( 
.A(n_6282),
.B(n_797),
.Y(n_6391)
);

AND2x2_ASAP7_75t_L g6392 ( 
.A(n_6288),
.B(n_798),
.Y(n_6392)
);

INVx1_ASAP7_75t_SL g6393 ( 
.A(n_6180),
.Y(n_6393)
);

AO21x2_ASAP7_75t_L g6394 ( 
.A1(n_6280),
.A2(n_798),
.B(n_800),
.Y(n_6394)
);

AND2x2_ASAP7_75t_L g6395 ( 
.A(n_6295),
.B(n_800),
.Y(n_6395)
);

AND2x2_ASAP7_75t_L g6396 ( 
.A(n_6309),
.B(n_801),
.Y(n_6396)
);

INVx2_ASAP7_75t_L g6397 ( 
.A(n_6205),
.Y(n_6397)
);

INVx1_ASAP7_75t_L g6398 ( 
.A(n_6138),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_6139),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_6250),
.Y(n_6400)
);

HB1xp67_ASAP7_75t_L g6401 ( 
.A(n_6058),
.Y(n_6401)
);

INVx2_ASAP7_75t_L g6402 ( 
.A(n_6065),
.Y(n_6402)
);

OR2x2_ASAP7_75t_L g6403 ( 
.A(n_6178),
.B(n_802),
.Y(n_6403)
);

AND2x2_ASAP7_75t_L g6404 ( 
.A(n_6154),
.B(n_802),
.Y(n_6404)
);

HB1xp67_ASAP7_75t_L g6405 ( 
.A(n_6253),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_6260),
.Y(n_6406)
);

AND2x2_ASAP7_75t_L g6407 ( 
.A(n_6167),
.B(n_803),
.Y(n_6407)
);

AOI221xp5_ASAP7_75t_L g6408 ( 
.A1(n_6155),
.A2(n_805),
.B1(n_803),
.B2(n_804),
.C(n_806),
.Y(n_6408)
);

AND2x2_ASAP7_75t_L g6409 ( 
.A(n_6188),
.B(n_805),
.Y(n_6409)
);

AO21x2_ASAP7_75t_L g6410 ( 
.A1(n_6303),
.A2(n_807),
.B(n_808),
.Y(n_6410)
);

INVx2_ASAP7_75t_L g6411 ( 
.A(n_6089),
.Y(n_6411)
);

INVx2_ASAP7_75t_L g6412 ( 
.A(n_6163),
.Y(n_6412)
);

NAND2xp5_ASAP7_75t_L g6413 ( 
.A(n_6183),
.B(n_810),
.Y(n_6413)
);

INVx2_ASAP7_75t_L g6414 ( 
.A(n_6129),
.Y(n_6414)
);

AND2x2_ASAP7_75t_L g6415 ( 
.A(n_6185),
.B(n_811),
.Y(n_6415)
);

INVx2_ASAP7_75t_L g6416 ( 
.A(n_6222),
.Y(n_6416)
);

NAND2xp5_ASAP7_75t_L g6417 ( 
.A(n_6242),
.B(n_6152),
.Y(n_6417)
);

NAND2xp5_ASAP7_75t_L g6418 ( 
.A(n_6207),
.B(n_811),
.Y(n_6418)
);

INVx2_ASAP7_75t_L g6419 ( 
.A(n_6068),
.Y(n_6419)
);

BUFx2_ASAP7_75t_L g6420 ( 
.A(n_6272),
.Y(n_6420)
);

INVxp67_ASAP7_75t_SL g6421 ( 
.A(n_6082),
.Y(n_6421)
);

NAND2xp5_ASAP7_75t_L g6422 ( 
.A(n_6187),
.B(n_813),
.Y(n_6422)
);

OAI21xp5_ASAP7_75t_SL g6423 ( 
.A1(n_6284),
.A2(n_817),
.B(n_816),
.Y(n_6423)
);

OR2x2_ASAP7_75t_L g6424 ( 
.A(n_6150),
.B(n_814),
.Y(n_6424)
);

AOI22xp33_ASAP7_75t_L g6425 ( 
.A1(n_6064),
.A2(n_818),
.B1(n_814),
.B2(n_817),
.Y(n_6425)
);

HB1xp67_ASAP7_75t_L g6426 ( 
.A(n_6281),
.Y(n_6426)
);

INVx2_ASAP7_75t_L g6427 ( 
.A(n_6080),
.Y(n_6427)
);

OAI221xp5_ASAP7_75t_L g6428 ( 
.A1(n_6208),
.A2(n_820),
.B1(n_818),
.B2(n_819),
.C(n_821),
.Y(n_6428)
);

OAI22xp5_ASAP7_75t_L g6429 ( 
.A1(n_6056),
.A2(n_821),
.B1(n_819),
.B2(n_820),
.Y(n_6429)
);

INVx4_ASAP7_75t_L g6430 ( 
.A(n_6103),
.Y(n_6430)
);

NAND3xp33_ASAP7_75t_L g6431 ( 
.A(n_6071),
.B(n_822),
.C(n_823),
.Y(n_6431)
);

INVx2_ASAP7_75t_L g6432 ( 
.A(n_6084),
.Y(n_6432)
);

INVx3_ASAP7_75t_L g6433 ( 
.A(n_6158),
.Y(n_6433)
);

AOI22xp33_ASAP7_75t_L g6434 ( 
.A1(n_6100),
.A2(n_824),
.B1(n_822),
.B2(n_823),
.Y(n_6434)
);

NAND4xp25_ASAP7_75t_L g6435 ( 
.A(n_6124),
.B(n_6098),
.C(n_6234),
.D(n_6066),
.Y(n_6435)
);

AND2x4_ASAP7_75t_L g6436 ( 
.A(n_6169),
.B(n_824),
.Y(n_6436)
);

AOI322xp5_ASAP7_75t_L g6437 ( 
.A1(n_6176),
.A2(n_831),
.A3(n_830),
.B1(n_827),
.B2(n_825),
.C1(n_826),
.C2(n_828),
.Y(n_6437)
);

AND2x2_ASAP7_75t_L g6438 ( 
.A(n_6232),
.B(n_826),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6264),
.Y(n_6439)
);

INVx1_ASAP7_75t_L g6440 ( 
.A(n_6274),
.Y(n_6440)
);

HB1xp67_ASAP7_75t_L g6441 ( 
.A(n_6296),
.Y(n_6441)
);

INVx2_ASAP7_75t_L g6442 ( 
.A(n_6087),
.Y(n_6442)
);

AND2x2_ASAP7_75t_L g6443 ( 
.A(n_6245),
.B(n_828),
.Y(n_6443)
);

AND2x2_ASAP7_75t_L g6444 ( 
.A(n_6165),
.B(n_831),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_6301),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_6302),
.Y(n_6446)
);

INVxp67_ASAP7_75t_L g6447 ( 
.A(n_6248),
.Y(n_6447)
);

INVxp67_ASAP7_75t_L g6448 ( 
.A(n_6249),
.Y(n_6448)
);

AND2x2_ASAP7_75t_L g6449 ( 
.A(n_6239),
.B(n_832),
.Y(n_6449)
);

INVx1_ASAP7_75t_SL g6450 ( 
.A(n_6079),
.Y(n_6450)
);

AND2x2_ASAP7_75t_L g6451 ( 
.A(n_6172),
.B(n_832),
.Y(n_6451)
);

CKINVDCx5p33_ASAP7_75t_R g6452 ( 
.A(n_6193),
.Y(n_6452)
);

BUFx3_ASAP7_75t_L g6453 ( 
.A(n_6061),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_6304),
.Y(n_6454)
);

INVx1_ASAP7_75t_L g6455 ( 
.A(n_6308),
.Y(n_6455)
);

AND2x2_ASAP7_75t_L g6456 ( 
.A(n_6174),
.B(n_833),
.Y(n_6456)
);

AND2x2_ASAP7_75t_L g6457 ( 
.A(n_6175),
.B(n_833),
.Y(n_6457)
);

INVx2_ASAP7_75t_L g6458 ( 
.A(n_6090),
.Y(n_6458)
);

INVx2_ASAP7_75t_L g6459 ( 
.A(n_6102),
.Y(n_6459)
);

OR2x2_ASAP7_75t_L g6460 ( 
.A(n_6110),
.B(n_834),
.Y(n_6460)
);

NAND2xp5_ASAP7_75t_L g6461 ( 
.A(n_6182),
.B(n_834),
.Y(n_6461)
);

OR2x2_ASAP7_75t_L g6462 ( 
.A(n_6146),
.B(n_6117),
.Y(n_6462)
);

HB1xp67_ASAP7_75t_L g6463 ( 
.A(n_6104),
.Y(n_6463)
);

BUFx2_ASAP7_75t_L g6464 ( 
.A(n_6162),
.Y(n_6464)
);

INVx1_ASAP7_75t_SL g6465 ( 
.A(n_6133),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_6132),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_6149),
.Y(n_6467)
);

NAND2xp5_ASAP7_75t_L g6468 ( 
.A(n_6121),
.B(n_836),
.Y(n_6468)
);

AOI221xp5_ASAP7_75t_L g6469 ( 
.A1(n_6093),
.A2(n_838),
.B1(n_836),
.B2(n_837),
.C(n_839),
.Y(n_6469)
);

AND2x4_ASAP7_75t_L g6470 ( 
.A(n_6156),
.B(n_839),
.Y(n_6470)
);

AND2x2_ASAP7_75t_L g6471 ( 
.A(n_6235),
.B(n_840),
.Y(n_6471)
);

INVx1_ASAP7_75t_L g6472 ( 
.A(n_6122),
.Y(n_6472)
);

OAI221xp5_ASAP7_75t_L g6473 ( 
.A1(n_6293),
.A2(n_842),
.B1(n_840),
.B2(n_841),
.C(n_843),
.Y(n_6473)
);

HB1xp67_ASAP7_75t_L g6474 ( 
.A(n_6289),
.Y(n_6474)
);

INVx1_ASAP7_75t_SL g6475 ( 
.A(n_6265),
.Y(n_6475)
);

INVx1_ASAP7_75t_L g6476 ( 
.A(n_6125),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_6119),
.Y(n_6477)
);

AND2x2_ASAP7_75t_L g6478 ( 
.A(n_6157),
.B(n_841),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_6055),
.Y(n_6479)
);

INVx2_ASAP7_75t_L g6480 ( 
.A(n_6160),
.Y(n_6480)
);

INVx1_ASAP7_75t_L g6481 ( 
.A(n_6055),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_6278),
.Y(n_6482)
);

BUFx3_ASAP7_75t_L g6483 ( 
.A(n_6199),
.Y(n_6483)
);

OR2x2_ASAP7_75t_L g6484 ( 
.A(n_6075),
.B(n_842),
.Y(n_6484)
);

OAI322xp33_ASAP7_75t_L g6485 ( 
.A1(n_6190),
.A2(n_6101),
.A3(n_6231),
.B1(n_6140),
.B2(n_6120),
.C1(n_6226),
.C2(n_6113),
.Y(n_6485)
);

INVx1_ASAP7_75t_L g6486 ( 
.A(n_6278),
.Y(n_6486)
);

OAI21xp33_ASAP7_75t_L g6487 ( 
.A1(n_6081),
.A2(n_843),
.B(n_844),
.Y(n_6487)
);

AOI21xp33_ASAP7_75t_L g6488 ( 
.A1(n_6095),
.A2(n_844),
.B(n_846),
.Y(n_6488)
);

INVx3_ASAP7_75t_L g6489 ( 
.A(n_6137),
.Y(n_6489)
);

HB1xp67_ASAP7_75t_L g6490 ( 
.A(n_6312),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_6258),
.Y(n_6491)
);

INVx1_ASAP7_75t_L g6492 ( 
.A(n_6111),
.Y(n_6492)
);

INVx3_ASAP7_75t_L g6493 ( 
.A(n_6092),
.Y(n_6493)
);

AO221x2_ASAP7_75t_L g6494 ( 
.A1(n_6219),
.A2(n_848),
.B1(n_846),
.B2(n_847),
.C(n_849),
.Y(n_6494)
);

BUFx2_ASAP7_75t_L g6495 ( 
.A(n_6215),
.Y(n_6495)
);

INVx2_ASAP7_75t_L g6496 ( 
.A(n_6196),
.Y(n_6496)
);

AND2x2_ASAP7_75t_L g6497 ( 
.A(n_6269),
.B(n_847),
.Y(n_6497)
);

OAI33xp33_ASAP7_75t_L g6498 ( 
.A1(n_6218),
.A2(n_851),
.A3(n_854),
.B1(n_848),
.B2(n_850),
.B3(n_853),
.Y(n_6498)
);

INVx1_ASAP7_75t_L g6499 ( 
.A(n_6200),
.Y(n_6499)
);

INVx4_ASAP7_75t_L g6500 ( 
.A(n_6142),
.Y(n_6500)
);

AND2x2_ASAP7_75t_L g6501 ( 
.A(n_6320),
.B(n_6326),
.Y(n_6501)
);

INVx2_ASAP7_75t_L g6502 ( 
.A(n_6324),
.Y(n_6502)
);

INVx1_ASAP7_75t_L g6503 ( 
.A(n_6349),
.Y(n_6503)
);

NAND2xp5_ASAP7_75t_L g6504 ( 
.A(n_6421),
.B(n_6240),
.Y(n_6504)
);

OR2x2_ASAP7_75t_L g6505 ( 
.A(n_6325),
.B(n_6179),
.Y(n_6505)
);

AND2x2_ASAP7_75t_L g6506 ( 
.A(n_6350),
.B(n_6240),
.Y(n_6506)
);

NAND2xp5_ASAP7_75t_L g6507 ( 
.A(n_6450),
.B(n_6170),
.Y(n_6507)
);

INVx1_ASAP7_75t_L g6508 ( 
.A(n_6401),
.Y(n_6508)
);

AND2x2_ASAP7_75t_L g6509 ( 
.A(n_6323),
.B(n_6276),
.Y(n_6509)
);

INVx2_ASAP7_75t_L g6510 ( 
.A(n_6324),
.Y(n_6510)
);

AND2x2_ASAP7_75t_L g6511 ( 
.A(n_6336),
.B(n_6074),
.Y(n_6511)
);

AND2x2_ASAP7_75t_L g6512 ( 
.A(n_6397),
.B(n_6134),
.Y(n_6512)
);

NAND2xp5_ASAP7_75t_L g6513 ( 
.A(n_6318),
.B(n_6173),
.Y(n_6513)
);

INVx2_ASAP7_75t_L g6514 ( 
.A(n_6483),
.Y(n_6514)
);

NAND2xp5_ASAP7_75t_L g6515 ( 
.A(n_6465),
.B(n_6307),
.Y(n_6515)
);

NAND2xp5_ASAP7_75t_L g6516 ( 
.A(n_6475),
.B(n_6313),
.Y(n_6516)
);

AND2x2_ASAP7_75t_L g6517 ( 
.A(n_6354),
.B(n_6106),
.Y(n_6517)
);

NAND2xp5_ASAP7_75t_L g6518 ( 
.A(n_6315),
.B(n_6244),
.Y(n_6518)
);

AND2x2_ASAP7_75t_L g6519 ( 
.A(n_6363),
.B(n_6220),
.Y(n_6519)
);

NAND2xp5_ASAP7_75t_L g6520 ( 
.A(n_6474),
.B(n_6181),
.Y(n_6520)
);

OR2x2_ASAP7_75t_L g6521 ( 
.A(n_6351),
.B(n_6086),
.Y(n_6521)
);

OR2x2_ASAP7_75t_L g6522 ( 
.A(n_6368),
.B(n_6214),
.Y(n_6522)
);

NOR2xp33_ASAP7_75t_L g6523 ( 
.A(n_6393),
.B(n_6227),
.Y(n_6523)
);

AND2x4_ASAP7_75t_L g6524 ( 
.A(n_6430),
.B(n_6168),
.Y(n_6524)
);

INVx3_ASAP7_75t_L g6525 ( 
.A(n_6342),
.Y(n_6525)
);

AND2x2_ASAP7_75t_L g6526 ( 
.A(n_6362),
.B(n_6233),
.Y(n_6526)
);

NAND2xp5_ASAP7_75t_L g6527 ( 
.A(n_6490),
.B(n_6447),
.Y(n_6527)
);

AND2x2_ASAP7_75t_L g6528 ( 
.A(n_6374),
.B(n_6217),
.Y(n_6528)
);

INVx2_ASAP7_75t_L g6529 ( 
.A(n_6453),
.Y(n_6529)
);

INVx1_ASAP7_75t_SL g6530 ( 
.A(n_6348),
.Y(n_6530)
);

INVx3_ASAP7_75t_L g6531 ( 
.A(n_6358),
.Y(n_6531)
);

AND2x4_ASAP7_75t_L g6532 ( 
.A(n_6379),
.B(n_6216),
.Y(n_6532)
);

AND2x2_ASAP7_75t_L g6533 ( 
.A(n_6493),
.B(n_6237),
.Y(n_6533)
);

AND2x2_ASAP7_75t_L g6534 ( 
.A(n_6433),
.B(n_6108),
.Y(n_6534)
);

OR2x2_ASAP7_75t_L g6535 ( 
.A(n_6384),
.B(n_6147),
.Y(n_6535)
);

INVx1_ASAP7_75t_L g6536 ( 
.A(n_6405),
.Y(n_6536)
);

HB1xp67_ASAP7_75t_L g6537 ( 
.A(n_6330),
.Y(n_6537)
);

INVx1_ASAP7_75t_L g6538 ( 
.A(n_6426),
.Y(n_6538)
);

INVx1_ASAP7_75t_L g6539 ( 
.A(n_6441),
.Y(n_6539)
);

INVx1_ASAP7_75t_SL g6540 ( 
.A(n_6452),
.Y(n_6540)
);

AND2x2_ASAP7_75t_L g6541 ( 
.A(n_6335),
.B(n_6085),
.Y(n_6541)
);

AND2x2_ASAP7_75t_L g6542 ( 
.A(n_6380),
.B(n_6224),
.Y(n_6542)
);

AND2x4_ASAP7_75t_L g6543 ( 
.A(n_6489),
.B(n_6241),
.Y(n_6543)
);

INVx1_ASAP7_75t_L g6544 ( 
.A(n_6420),
.Y(n_6544)
);

AND2x2_ASAP7_75t_L g6545 ( 
.A(n_6340),
.B(n_6500),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_6448),
.B(n_6464),
.Y(n_6546)
);

NAND2xp5_ASAP7_75t_L g6547 ( 
.A(n_6499),
.B(n_6141),
.Y(n_6547)
);

NAND2xp5_ASAP7_75t_L g6548 ( 
.A(n_6394),
.B(n_6141),
.Y(n_6548)
);

INVx2_ASAP7_75t_L g6549 ( 
.A(n_6462),
.Y(n_6549)
);

NAND3xp33_ASAP7_75t_L g6550 ( 
.A(n_6322),
.B(n_6361),
.C(n_6495),
.Y(n_6550)
);

AND2x2_ASAP7_75t_L g6551 ( 
.A(n_6373),
.B(n_6083),
.Y(n_6551)
);

INVx1_ASAP7_75t_L g6552 ( 
.A(n_6463),
.Y(n_6552)
);

INVxp67_ASAP7_75t_L g6553 ( 
.A(n_6357),
.Y(n_6553)
);

INVxp67_ASAP7_75t_SL g6554 ( 
.A(n_6334),
.Y(n_6554)
);

INVx1_ASAP7_75t_L g6555 ( 
.A(n_6472),
.Y(n_6555)
);

NAND2x1_ASAP7_75t_SL g6556 ( 
.A(n_6496),
.B(n_6228),
.Y(n_6556)
);

INVx2_ASAP7_75t_L g6557 ( 
.A(n_6338),
.Y(n_6557)
);

OR2x2_ASAP7_75t_L g6558 ( 
.A(n_6417),
.B(n_6212),
.Y(n_6558)
);

AND2x2_ASAP7_75t_L g6559 ( 
.A(n_6492),
.B(n_6246),
.Y(n_6559)
);

AND2x2_ASAP7_75t_L g6560 ( 
.A(n_6491),
.B(n_6198),
.Y(n_6560)
);

NAND3xp33_ASAP7_75t_L g6561 ( 
.A(n_6431),
.B(n_6118),
.C(n_6054),
.Y(n_6561)
);

INVx2_ASAP7_75t_L g6562 ( 
.A(n_6343),
.Y(n_6562)
);

AND2x4_ASAP7_75t_L g6563 ( 
.A(n_6317),
.B(n_6171),
.Y(n_6563)
);

AND2x4_ASAP7_75t_L g6564 ( 
.A(n_6414),
.B(n_6204),
.Y(n_6564)
);

INVx1_ASAP7_75t_L g6565 ( 
.A(n_6476),
.Y(n_6565)
);

AND2x4_ASAP7_75t_L g6566 ( 
.A(n_6337),
.B(n_6287),
.Y(n_6566)
);

OR2x2_ASAP7_75t_L g6567 ( 
.A(n_6383),
.B(n_6229),
.Y(n_6567)
);

AND2x2_ASAP7_75t_L g6568 ( 
.A(n_6412),
.B(n_6109),
.Y(n_6568)
);

OR2x2_ASAP7_75t_L g6569 ( 
.A(n_6416),
.B(n_6189),
.Y(n_6569)
);

INVx1_ASAP7_75t_L g6570 ( 
.A(n_6341),
.Y(n_6570)
);

BUFx2_ASAP7_75t_L g6571 ( 
.A(n_6359),
.Y(n_6571)
);

INVx1_ASAP7_75t_SL g6572 ( 
.A(n_6321),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_6347),
.Y(n_6573)
);

INVx1_ASAP7_75t_L g6574 ( 
.A(n_6352),
.Y(n_6574)
);

INVx1_ASAP7_75t_SL g6575 ( 
.A(n_6370),
.Y(n_6575)
);

AND2x2_ASAP7_75t_L g6576 ( 
.A(n_6480),
.B(n_6116),
.Y(n_6576)
);

NAND2xp5_ASAP7_75t_L g6577 ( 
.A(n_6410),
.B(n_6279),
.Y(n_6577)
);

AND2x4_ASAP7_75t_L g6578 ( 
.A(n_6333),
.B(n_6192),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_6376),
.Y(n_6579)
);

INVx2_ASAP7_75t_L g6580 ( 
.A(n_6360),
.Y(n_6580)
);

NOR2x1p5_ASAP7_75t_L g6581 ( 
.A(n_6388),
.B(n_6135),
.Y(n_6581)
);

AND2x2_ASAP7_75t_L g6582 ( 
.A(n_6443),
.B(n_6144),
.Y(n_6582)
);

AND2x2_ASAP7_75t_L g6583 ( 
.A(n_6438),
.B(n_6161),
.Y(n_6583)
);

NOR2x1_ASAP7_75t_L g6584 ( 
.A(n_6424),
.B(n_6191),
.Y(n_6584)
);

INVx1_ASAP7_75t_L g6585 ( 
.A(n_6377),
.Y(n_6585)
);

INVx2_ASAP7_75t_L g6586 ( 
.A(n_6460),
.Y(n_6586)
);

AND2x2_ASAP7_75t_L g6587 ( 
.A(n_6471),
.B(n_6148),
.Y(n_6587)
);

AND2x2_ASAP7_75t_L g6588 ( 
.A(n_6478),
.B(n_6300),
.Y(n_6588)
);

OR2x2_ASAP7_75t_L g6589 ( 
.A(n_6364),
.B(n_6311),
.Y(n_6589)
);

INVx2_ASAP7_75t_L g6590 ( 
.A(n_6402),
.Y(n_6590)
);

NAND2xp5_ASAP7_75t_L g6591 ( 
.A(n_6479),
.B(n_6259),
.Y(n_6591)
);

INVx1_ASAP7_75t_L g6592 ( 
.A(n_6382),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_6385),
.Y(n_6593)
);

INVx2_ASAP7_75t_L g6594 ( 
.A(n_6411),
.Y(n_6594)
);

OR2x2_ASAP7_75t_L g6595 ( 
.A(n_6403),
.B(n_6332),
.Y(n_6595)
);

OR2x2_ASAP7_75t_L g6596 ( 
.A(n_6419),
.B(n_6427),
.Y(n_6596)
);

AND2x2_ASAP7_75t_L g6597 ( 
.A(n_6407),
.B(n_6088),
.Y(n_6597)
);

NAND2xp5_ASAP7_75t_L g6598 ( 
.A(n_6481),
.B(n_6268),
.Y(n_6598)
);

OAI211xp5_ASAP7_75t_SL g6599 ( 
.A1(n_6314),
.A2(n_6273),
.B(n_6286),
.C(n_6283),
.Y(n_6599)
);

NAND2xp5_ASAP7_75t_L g6600 ( 
.A(n_6482),
.B(n_6486),
.Y(n_6600)
);

NAND2xp5_ASAP7_75t_L g6601 ( 
.A(n_6378),
.B(n_6097),
.Y(n_6601)
);

AOI21xp5_ASAP7_75t_L g6602 ( 
.A1(n_6485),
.A2(n_6356),
.B(n_6422),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_6387),
.Y(n_6603)
);

AND2x2_ASAP7_75t_L g6604 ( 
.A(n_6444),
.B(n_6151),
.Y(n_6604)
);

AND2x4_ASAP7_75t_L g6605 ( 
.A(n_6367),
.B(n_6247),
.Y(n_6605)
);

AND2x2_ASAP7_75t_L g6606 ( 
.A(n_6451),
.B(n_850),
.Y(n_6606)
);

AND2x2_ASAP7_75t_L g6607 ( 
.A(n_6456),
.B(n_851),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6390),
.Y(n_6608)
);

AND2x2_ASAP7_75t_L g6609 ( 
.A(n_6457),
.B(n_854),
.Y(n_6609)
);

INVx3_ASAP7_75t_L g6610 ( 
.A(n_6436),
.Y(n_6610)
);

INVx2_ASAP7_75t_L g6611 ( 
.A(n_6369),
.Y(n_6611)
);

INVx1_ASAP7_75t_L g6612 ( 
.A(n_6398),
.Y(n_6612)
);

OR2x2_ASAP7_75t_L g6613 ( 
.A(n_6432),
.B(n_6442),
.Y(n_6613)
);

BUFx2_ASAP7_75t_L g6614 ( 
.A(n_6328),
.Y(n_6614)
);

AND2x2_ASAP7_75t_L g6615 ( 
.A(n_6449),
.B(n_855),
.Y(n_6615)
);

INVx2_ASAP7_75t_L g6616 ( 
.A(n_6458),
.Y(n_6616)
);

INVx1_ASAP7_75t_L g6617 ( 
.A(n_6399),
.Y(n_6617)
);

INVx2_ASAP7_75t_L g6618 ( 
.A(n_6459),
.Y(n_6618)
);

INVx1_ASAP7_75t_L g6619 ( 
.A(n_6400),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6406),
.Y(n_6620)
);

NAND2xp5_ASAP7_75t_L g6621 ( 
.A(n_6415),
.B(n_855),
.Y(n_6621)
);

AND2x2_ASAP7_75t_L g6622 ( 
.A(n_6327),
.B(n_856),
.Y(n_6622)
);

NAND2xp5_ASAP7_75t_L g6623 ( 
.A(n_6409),
.B(n_856),
.Y(n_6623)
);

NAND2xp5_ASAP7_75t_SL g6624 ( 
.A(n_6366),
.B(n_6429),
.Y(n_6624)
);

OR2x2_ASAP7_75t_L g6625 ( 
.A(n_6477),
.B(n_857),
.Y(n_6625)
);

NAND4xp25_ASAP7_75t_L g6626 ( 
.A(n_6435),
.B(n_860),
.C(n_858),
.D(n_859),
.Y(n_6626)
);

NAND2xp5_ASAP7_75t_L g6627 ( 
.A(n_6418),
.B(n_860),
.Y(n_6627)
);

INVx2_ASAP7_75t_L g6628 ( 
.A(n_6404),
.Y(n_6628)
);

INVx1_ASAP7_75t_L g6629 ( 
.A(n_6439),
.Y(n_6629)
);

AND2x2_ASAP7_75t_L g6630 ( 
.A(n_6331),
.B(n_6497),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_6344),
.B(n_861),
.Y(n_6631)
);

AND2x2_ASAP7_75t_L g6632 ( 
.A(n_6355),
.B(n_861),
.Y(n_6632)
);

HB1xp67_ASAP7_75t_L g6633 ( 
.A(n_6466),
.Y(n_6633)
);

AND2x2_ASAP7_75t_L g6634 ( 
.A(n_6381),
.B(n_862),
.Y(n_6634)
);

INVx1_ASAP7_75t_L g6635 ( 
.A(n_6440),
.Y(n_6635)
);

INVx2_ASAP7_75t_L g6636 ( 
.A(n_6389),
.Y(n_6636)
);

INVx1_ASAP7_75t_L g6637 ( 
.A(n_6537),
.Y(n_6637)
);

NAND2xp5_ASAP7_75t_L g6638 ( 
.A(n_6554),
.B(n_6461),
.Y(n_6638)
);

NAND4xp75_ASAP7_75t_SL g6639 ( 
.A(n_6506),
.B(n_6353),
.C(n_6392),
.D(n_6391),
.Y(n_6639)
);

HB1xp67_ASAP7_75t_L g6640 ( 
.A(n_6553),
.Y(n_6640)
);

AND2x2_ASAP7_75t_L g6641 ( 
.A(n_6525),
.B(n_6395),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_6503),
.Y(n_6642)
);

INVx4_ASAP7_75t_L g6643 ( 
.A(n_6531),
.Y(n_6643)
);

OR2x2_ASAP7_75t_L g6644 ( 
.A(n_6572),
.B(n_6467),
.Y(n_6644)
);

XNOR2x2_ASAP7_75t_L g6645 ( 
.A(n_6550),
.B(n_6413),
.Y(n_6645)
);

XOR2x2_ASAP7_75t_L g6646 ( 
.A(n_6561),
.B(n_6345),
.Y(n_6646)
);

NAND4xp75_ASAP7_75t_L g6647 ( 
.A(n_6584),
.B(n_6546),
.C(n_6527),
.D(n_6601),
.Y(n_6647)
);

NAND4xp75_ASAP7_75t_SL g6648 ( 
.A(n_6501),
.B(n_6396),
.C(n_6365),
.D(n_6423),
.Y(n_6648)
);

AND2x2_ASAP7_75t_L g6649 ( 
.A(n_6517),
.B(n_6470),
.Y(n_6649)
);

INVx1_ASAP7_75t_L g6650 ( 
.A(n_6508),
.Y(n_6650)
);

INVx2_ASAP7_75t_L g6651 ( 
.A(n_6519),
.Y(n_6651)
);

INVx1_ASAP7_75t_L g6652 ( 
.A(n_6536),
.Y(n_6652)
);

OR2x2_ASAP7_75t_L g6653 ( 
.A(n_6535),
.B(n_6371),
.Y(n_6653)
);

AND2x4_ASAP7_75t_L g6654 ( 
.A(n_6530),
.B(n_6339),
.Y(n_6654)
);

NAND3xp33_ASAP7_75t_L g6655 ( 
.A(n_6614),
.B(n_6319),
.C(n_6437),
.Y(n_6655)
);

XNOR2xp5_ASAP7_75t_L g6656 ( 
.A(n_6581),
.B(n_6425),
.Y(n_6656)
);

INVx2_ASAP7_75t_L g6657 ( 
.A(n_6502),
.Y(n_6657)
);

OR2x2_ASAP7_75t_L g6658 ( 
.A(n_6504),
.B(n_6522),
.Y(n_6658)
);

INVx1_ASAP7_75t_L g6659 ( 
.A(n_6538),
.Y(n_6659)
);

NOR2xp33_ASAP7_75t_L g6660 ( 
.A(n_6540),
.B(n_6575),
.Y(n_6660)
);

AOI22xp5_ASAP7_75t_L g6661 ( 
.A1(n_6513),
.A2(n_6494),
.B1(n_6346),
.B2(n_6498),
.Y(n_6661)
);

AND2x2_ASAP7_75t_L g6662 ( 
.A(n_6551),
.B(n_6445),
.Y(n_6662)
);

INVx2_ASAP7_75t_L g6663 ( 
.A(n_6510),
.Y(n_6663)
);

NAND2xp5_ASAP7_75t_L g6664 ( 
.A(n_6582),
.B(n_6372),
.Y(n_6664)
);

INVx1_ASAP7_75t_L g6665 ( 
.A(n_6539),
.Y(n_6665)
);

INVx1_ASAP7_75t_L g6666 ( 
.A(n_6552),
.Y(n_6666)
);

BUFx2_ASAP7_75t_L g6667 ( 
.A(n_6556),
.Y(n_6667)
);

INVx2_ASAP7_75t_L g6668 ( 
.A(n_6543),
.Y(n_6668)
);

INVx1_ASAP7_75t_L g6669 ( 
.A(n_6633),
.Y(n_6669)
);

INVx2_ASAP7_75t_SL g6670 ( 
.A(n_6545),
.Y(n_6670)
);

NOR4xp25_ASAP7_75t_L g6671 ( 
.A(n_6599),
.B(n_6488),
.C(n_6428),
.D(n_6473),
.Y(n_6671)
);

XOR2x2_ASAP7_75t_L g6672 ( 
.A(n_6624),
.B(n_6375),
.Y(n_6672)
);

INVx1_ASAP7_75t_L g6673 ( 
.A(n_6625),
.Y(n_6673)
);

INVx1_ASAP7_75t_L g6674 ( 
.A(n_6611),
.Y(n_6674)
);

INVx1_ASAP7_75t_L g6675 ( 
.A(n_6595),
.Y(n_6675)
);

NAND4xp75_ASAP7_75t_SL g6676 ( 
.A(n_6523),
.B(n_6408),
.C(n_6487),
.D(n_6329),
.Y(n_6676)
);

INVx4_ASAP7_75t_L g6677 ( 
.A(n_6622),
.Y(n_6677)
);

NAND4xp75_ASAP7_75t_SL g6678 ( 
.A(n_6541),
.B(n_6469),
.C(n_6434),
.D(n_6316),
.Y(n_6678)
);

NOR4xp25_ASAP7_75t_L g6679 ( 
.A(n_6626),
.B(n_6468),
.C(n_6386),
.D(n_6484),
.Y(n_6679)
);

AND2x2_ASAP7_75t_L g6680 ( 
.A(n_6630),
.B(n_6446),
.Y(n_6680)
);

AND2x2_ASAP7_75t_L g6681 ( 
.A(n_6509),
.B(n_6454),
.Y(n_6681)
);

NAND4xp75_ASAP7_75t_L g6682 ( 
.A(n_6602),
.B(n_6455),
.C(n_864),
.D(n_862),
.Y(n_6682)
);

XNOR2xp5_ASAP7_75t_L g6683 ( 
.A(n_6511),
.B(n_863),
.Y(n_6683)
);

AND2x2_ASAP7_75t_L g6684 ( 
.A(n_6512),
.B(n_863),
.Y(n_6684)
);

INVxp67_ASAP7_75t_SL g6685 ( 
.A(n_6610),
.Y(n_6685)
);

XNOR2x2_ASAP7_75t_L g6686 ( 
.A(n_6577),
.B(n_866),
.Y(n_6686)
);

AND2x2_ASAP7_75t_L g6687 ( 
.A(n_6529),
.B(n_864),
.Y(n_6687)
);

NOR3xp33_ASAP7_75t_L g6688 ( 
.A(n_6591),
.B(n_866),
.C(n_867),
.Y(n_6688)
);

AND2x2_ASAP7_75t_L g6689 ( 
.A(n_6514),
.B(n_868),
.Y(n_6689)
);

NOR2xp33_ASAP7_75t_L g6690 ( 
.A(n_6605),
.B(n_868),
.Y(n_6690)
);

AOI22xp5_ASAP7_75t_SL g6691 ( 
.A1(n_6548),
.A2(n_6563),
.B1(n_6578),
.B2(n_6566),
.Y(n_6691)
);

NAND2xp5_ASAP7_75t_L g6692 ( 
.A(n_6526),
.B(n_869),
.Y(n_6692)
);

NOR3xp33_ASAP7_75t_L g6693 ( 
.A(n_6598),
.B(n_6520),
.C(n_6518),
.Y(n_6693)
);

NAND4xp75_ASAP7_75t_L g6694 ( 
.A(n_6544),
.B(n_871),
.C(n_869),
.D(n_870),
.Y(n_6694)
);

INVx1_ASAP7_75t_L g6695 ( 
.A(n_6586),
.Y(n_6695)
);

INVx2_ASAP7_75t_SL g6696 ( 
.A(n_6559),
.Y(n_6696)
);

NAND4xp75_ASAP7_75t_SL g6697 ( 
.A(n_6576),
.B(n_872),
.C(n_870),
.D(n_871),
.Y(n_6697)
);

NAND2xp5_ASAP7_75t_L g6698 ( 
.A(n_6533),
.B(n_872),
.Y(n_6698)
);

AOI22xp5_ASAP7_75t_L g6699 ( 
.A1(n_6524),
.A2(n_875),
.B1(n_873),
.B2(n_874),
.Y(n_6699)
);

NAND2xp5_ASAP7_75t_L g6700 ( 
.A(n_6588),
.B(n_875),
.Y(n_6700)
);

NAND4xp75_ASAP7_75t_L g6701 ( 
.A(n_6600),
.B(n_878),
.C(n_876),
.D(n_877),
.Y(n_6701)
);

INVx1_ASAP7_75t_SL g6702 ( 
.A(n_6534),
.Y(n_6702)
);

INVx2_ASAP7_75t_L g6703 ( 
.A(n_6528),
.Y(n_6703)
);

INVx1_ASAP7_75t_L g6704 ( 
.A(n_6549),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_6570),
.Y(n_6705)
);

AOI211x1_ASAP7_75t_L g6706 ( 
.A1(n_6507),
.A2(n_879),
.B(n_876),
.C(n_878),
.Y(n_6706)
);

INVx2_ASAP7_75t_L g6707 ( 
.A(n_6636),
.Y(n_6707)
);

INVx2_ASAP7_75t_L g6708 ( 
.A(n_6532),
.Y(n_6708)
);

NAND2xp5_ASAP7_75t_L g6709 ( 
.A(n_6583),
.B(n_880),
.Y(n_6709)
);

XOR2x2_ASAP7_75t_L g6710 ( 
.A(n_6597),
.B(n_881),
.Y(n_6710)
);

NAND4xp75_ASAP7_75t_SL g6711 ( 
.A(n_6568),
.B(n_883),
.C(n_881),
.D(n_882),
.Y(n_6711)
);

HB1xp67_ASAP7_75t_L g6712 ( 
.A(n_6564),
.Y(n_6712)
);

AND2x4_ASAP7_75t_L g6713 ( 
.A(n_6628),
.B(n_882),
.Y(n_6713)
);

OR2x6_ASAP7_75t_L g6714 ( 
.A(n_6515),
.B(n_6516),
.Y(n_6714)
);

INVx1_ASAP7_75t_L g6715 ( 
.A(n_6573),
.Y(n_6715)
);

AND2x2_ASAP7_75t_L g6716 ( 
.A(n_6542),
.B(n_884),
.Y(n_6716)
);

AND2x2_ASAP7_75t_L g6717 ( 
.A(n_6560),
.B(n_884),
.Y(n_6717)
);

INVx1_ASAP7_75t_L g6718 ( 
.A(n_6574),
.Y(n_6718)
);

INVx1_ASAP7_75t_L g6719 ( 
.A(n_6579),
.Y(n_6719)
);

HB1xp67_ASAP7_75t_L g6720 ( 
.A(n_6571),
.Y(n_6720)
);

INVx2_ASAP7_75t_L g6721 ( 
.A(n_6596),
.Y(n_6721)
);

NAND4xp75_ASAP7_75t_SL g6722 ( 
.A(n_6604),
.B(n_887),
.C(n_885),
.D(n_886),
.Y(n_6722)
);

INVx1_ASAP7_75t_L g6723 ( 
.A(n_6585),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_6592),
.Y(n_6724)
);

AND2x2_ASAP7_75t_L g6725 ( 
.A(n_6587),
.B(n_889),
.Y(n_6725)
);

NAND2xp5_ASAP7_75t_L g6726 ( 
.A(n_6616),
.B(n_889),
.Y(n_6726)
);

NAND4xp75_ASAP7_75t_L g6727 ( 
.A(n_6547),
.B(n_894),
.C(n_891),
.D(n_892),
.Y(n_6727)
);

INVx2_ASAP7_75t_L g6728 ( 
.A(n_6613),
.Y(n_6728)
);

NAND2xp5_ASAP7_75t_L g6729 ( 
.A(n_6618),
.B(n_891),
.Y(n_6729)
);

NOR2xp33_ASAP7_75t_L g6730 ( 
.A(n_6521),
.B(n_894),
.Y(n_6730)
);

XOR2x2_ASAP7_75t_L g6731 ( 
.A(n_6505),
.B(n_895),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_6593),
.Y(n_6732)
);

XNOR2xp5_ASAP7_75t_L g6733 ( 
.A(n_6615),
.B(n_895),
.Y(n_6733)
);

NAND4xp75_ASAP7_75t_L g6734 ( 
.A(n_6594),
.B(n_899),
.C(n_897),
.D(n_898),
.Y(n_6734)
);

NAND4xp75_ASAP7_75t_SL g6735 ( 
.A(n_6631),
.B(n_900),
.C(n_897),
.D(n_899),
.Y(n_6735)
);

NAND2xp5_ASAP7_75t_L g6736 ( 
.A(n_6590),
.B(n_901),
.Y(n_6736)
);

INVx1_ASAP7_75t_L g6737 ( 
.A(n_6603),
.Y(n_6737)
);

BUFx3_ASAP7_75t_L g6738 ( 
.A(n_6632),
.Y(n_6738)
);

OR2x2_ASAP7_75t_L g6739 ( 
.A(n_6558),
.B(n_901),
.Y(n_6739)
);

INVx2_ASAP7_75t_L g6740 ( 
.A(n_6567),
.Y(n_6740)
);

NOR4xp75_ASAP7_75t_L g6741 ( 
.A(n_6627),
.B(n_905),
.C(n_902),
.D(n_904),
.Y(n_6741)
);

AND2x4_ASAP7_75t_SL g6742 ( 
.A(n_6634),
.B(n_902),
.Y(n_6742)
);

INVx1_ASAP7_75t_L g6743 ( 
.A(n_6608),
.Y(n_6743)
);

AND2x2_ASAP7_75t_L g6744 ( 
.A(n_6606),
.B(n_904),
.Y(n_6744)
);

INVx1_ASAP7_75t_SL g6745 ( 
.A(n_6607),
.Y(n_6745)
);

XNOR2xp5_ASAP7_75t_L g6746 ( 
.A(n_6609),
.B(n_905),
.Y(n_6746)
);

INVx3_ASAP7_75t_SL g6747 ( 
.A(n_6569),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_6557),
.Y(n_6748)
);

AND2x2_ASAP7_75t_L g6749 ( 
.A(n_6562),
.B(n_906),
.Y(n_6749)
);

INVx1_ASAP7_75t_L g6750 ( 
.A(n_6612),
.Y(n_6750)
);

INVx1_ASAP7_75t_L g6751 ( 
.A(n_6617),
.Y(n_6751)
);

AND2x2_ASAP7_75t_L g6752 ( 
.A(n_6580),
.B(n_908),
.Y(n_6752)
);

XOR2x1_ASAP7_75t_L g6753 ( 
.A(n_6589),
.B(n_6555),
.Y(n_6753)
);

NAND4xp75_ASAP7_75t_L g6754 ( 
.A(n_6565),
.B(n_911),
.C(n_909),
.D(n_910),
.Y(n_6754)
);

NAND4xp75_ASAP7_75t_L g6755 ( 
.A(n_6619),
.B(n_911),
.C(n_909),
.D(n_910),
.Y(n_6755)
);

INVx1_ASAP7_75t_L g6756 ( 
.A(n_6620),
.Y(n_6756)
);

INVx3_ASAP7_75t_L g6757 ( 
.A(n_6629),
.Y(n_6757)
);

NOR4xp25_ASAP7_75t_L g6758 ( 
.A(n_6635),
.B(n_914),
.C(n_912),
.D(n_913),
.Y(n_6758)
);

AND4x1_ASAP7_75t_L g6759 ( 
.A(n_6623),
.B(n_916),
.C(n_912),
.D(n_914),
.Y(n_6759)
);

NAND3xp33_ASAP7_75t_L g6760 ( 
.A(n_6621),
.B(n_918),
.C(n_917),
.Y(n_6760)
);

INVx2_ASAP7_75t_L g6761 ( 
.A(n_6525),
.Y(n_6761)
);

INVx2_ASAP7_75t_L g6762 ( 
.A(n_6525),
.Y(n_6762)
);

BUFx3_ASAP7_75t_L g6763 ( 
.A(n_6525),
.Y(n_6763)
);

INVx1_ASAP7_75t_L g6764 ( 
.A(n_6537),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_6537),
.Y(n_6765)
);

NAND4xp75_ASAP7_75t_L g6766 ( 
.A(n_6584),
.B(n_919),
.C(n_916),
.D(n_918),
.Y(n_6766)
);

BUFx3_ASAP7_75t_L g6767 ( 
.A(n_6525),
.Y(n_6767)
);

OR2x2_ASAP7_75t_L g6768 ( 
.A(n_6572),
.B(n_920),
.Y(n_6768)
);

AND2x2_ASAP7_75t_L g6769 ( 
.A(n_6763),
.B(n_920),
.Y(n_6769)
);

INVx1_ASAP7_75t_SL g6770 ( 
.A(n_6747),
.Y(n_6770)
);

INVx1_ASAP7_75t_L g6771 ( 
.A(n_6720),
.Y(n_6771)
);

INVxp67_ASAP7_75t_L g6772 ( 
.A(n_6667),
.Y(n_6772)
);

NAND2xp5_ASAP7_75t_L g6773 ( 
.A(n_6685),
.B(n_921),
.Y(n_6773)
);

INVx1_ASAP7_75t_L g6774 ( 
.A(n_6640),
.Y(n_6774)
);

INVx1_ASAP7_75t_L g6775 ( 
.A(n_6712),
.Y(n_6775)
);

AND2x2_ASAP7_75t_L g6776 ( 
.A(n_6767),
.B(n_922),
.Y(n_6776)
);

INVx1_ASAP7_75t_L g6777 ( 
.A(n_6637),
.Y(n_6777)
);

AND2x2_ASAP7_75t_L g6778 ( 
.A(n_6761),
.B(n_923),
.Y(n_6778)
);

NAND2xp5_ASAP7_75t_L g6779 ( 
.A(n_6670),
.B(n_923),
.Y(n_6779)
);

NAND2xp5_ASAP7_75t_L g6780 ( 
.A(n_6758),
.B(n_924),
.Y(n_6780)
);

OAI21xp5_ASAP7_75t_L g6781 ( 
.A1(n_6655),
.A2(n_924),
.B(n_925),
.Y(n_6781)
);

AO221x1_ASAP7_75t_L g6782 ( 
.A1(n_6757),
.A2(n_928),
.B1(n_930),
.B2(n_927),
.C(n_929),
.Y(n_6782)
);

INVx2_ASAP7_75t_L g6783 ( 
.A(n_6762),
.Y(n_6783)
);

INVx2_ASAP7_75t_L g6784 ( 
.A(n_6643),
.Y(n_6784)
);

OAI22xp5_ASAP7_75t_L g6785 ( 
.A1(n_6661),
.A2(n_928),
.B1(n_929),
.B2(n_927),
.Y(n_6785)
);

NAND2xp33_ASAP7_75t_SL g6786 ( 
.A(n_6656),
.B(n_926),
.Y(n_6786)
);

INVxp67_ASAP7_75t_SL g6787 ( 
.A(n_6753),
.Y(n_6787)
);

OR2x2_ASAP7_75t_L g6788 ( 
.A(n_6745),
.B(n_932),
.Y(n_6788)
);

NAND3xp33_ASAP7_75t_L g6789 ( 
.A(n_6693),
.B(n_932),
.C(n_933),
.Y(n_6789)
);

NAND2xp5_ASAP7_75t_L g6790 ( 
.A(n_6706),
.B(n_934),
.Y(n_6790)
);

AOI22xp5_ASAP7_75t_L g6791 ( 
.A1(n_6647),
.A2(n_936),
.B1(n_934),
.B2(n_935),
.Y(n_6791)
);

AND2x2_ASAP7_75t_L g6792 ( 
.A(n_6641),
.B(n_936),
.Y(n_6792)
);

NAND2xp5_ASAP7_75t_L g6793 ( 
.A(n_6691),
.B(n_938),
.Y(n_6793)
);

INVx2_ASAP7_75t_L g6794 ( 
.A(n_6738),
.Y(n_6794)
);

AND2x4_ASAP7_75t_L g6795 ( 
.A(n_6696),
.B(n_6649),
.Y(n_6795)
);

NAND2xp5_ASAP7_75t_L g6796 ( 
.A(n_6677),
.B(n_938),
.Y(n_6796)
);

AND2x2_ASAP7_75t_L g6797 ( 
.A(n_6668),
.B(n_939),
.Y(n_6797)
);

INVx1_ASAP7_75t_L g6798 ( 
.A(n_6764),
.Y(n_6798)
);

NAND2xp5_ASAP7_75t_L g6799 ( 
.A(n_6702),
.B(n_939),
.Y(n_6799)
);

AND2x2_ASAP7_75t_L g6800 ( 
.A(n_6651),
.B(n_6662),
.Y(n_6800)
);

OR2x2_ASAP7_75t_L g6801 ( 
.A(n_6714),
.B(n_940),
.Y(n_6801)
);

AND2x2_ASAP7_75t_L g6802 ( 
.A(n_6725),
.B(n_940),
.Y(n_6802)
);

AND2x4_ASAP7_75t_L g6803 ( 
.A(n_6703),
.B(n_941),
.Y(n_6803)
);

AND2x2_ASAP7_75t_L g6804 ( 
.A(n_6660),
.B(n_941),
.Y(n_6804)
);

NAND2x1p5_ASAP7_75t_L g6805 ( 
.A(n_6759),
.B(n_942),
.Y(n_6805)
);

AOI21xp5_ASAP7_75t_L g6806 ( 
.A1(n_6646),
.A2(n_943),
.B(n_945),
.Y(n_6806)
);

INVx2_ASAP7_75t_L g6807 ( 
.A(n_6708),
.Y(n_6807)
);

INVxp67_ASAP7_75t_L g6808 ( 
.A(n_6766),
.Y(n_6808)
);

AND2x2_ASAP7_75t_L g6809 ( 
.A(n_6654),
.B(n_946),
.Y(n_6809)
);

OAI322xp33_ASAP7_75t_L g6810 ( 
.A1(n_6645),
.A2(n_953),
.A3(n_952),
.B1(n_948),
.B2(n_946),
.C1(n_947),
.C2(n_951),
.Y(n_6810)
);

HB1xp67_ASAP7_75t_L g6811 ( 
.A(n_6639),
.Y(n_6811)
);

INVxp67_ASAP7_75t_SL g6812 ( 
.A(n_6686),
.Y(n_6812)
);

NOR2x1_ASAP7_75t_L g6813 ( 
.A(n_6682),
.B(n_948),
.Y(n_6813)
);

INVx1_ASAP7_75t_L g6814 ( 
.A(n_6765),
.Y(n_6814)
);

INVxp67_ASAP7_75t_L g6815 ( 
.A(n_6727),
.Y(n_6815)
);

AND2x2_ASAP7_75t_L g6816 ( 
.A(n_6680),
.B(n_951),
.Y(n_6816)
);

NAND2xp5_ASAP7_75t_L g6817 ( 
.A(n_6671),
.B(n_952),
.Y(n_6817)
);

NAND2xp5_ASAP7_75t_L g6818 ( 
.A(n_6716),
.B(n_6688),
.Y(n_6818)
);

INVx1_ASAP7_75t_L g6819 ( 
.A(n_6675),
.Y(n_6819)
);

NAND2xp5_ASAP7_75t_L g6820 ( 
.A(n_6717),
.B(n_953),
.Y(n_6820)
);

INVx1_ASAP7_75t_SL g6821 ( 
.A(n_6742),
.Y(n_6821)
);

AND2x2_ASAP7_75t_L g6822 ( 
.A(n_6657),
.B(n_954),
.Y(n_6822)
);

NAND2xp5_ASAP7_75t_L g6823 ( 
.A(n_6710),
.B(n_954),
.Y(n_6823)
);

INVx2_ASAP7_75t_L g6824 ( 
.A(n_6684),
.Y(n_6824)
);

NAND2xp5_ASAP7_75t_L g6825 ( 
.A(n_6679),
.B(n_955),
.Y(n_6825)
);

OAI21xp33_ASAP7_75t_SL g6826 ( 
.A1(n_6648),
.A2(n_955),
.B(n_956),
.Y(n_6826)
);

NAND2xp5_ASAP7_75t_L g6827 ( 
.A(n_6749),
.B(n_956),
.Y(n_6827)
);

OR2x2_ASAP7_75t_L g6828 ( 
.A(n_6714),
.B(n_957),
.Y(n_6828)
);

OR2x2_ASAP7_75t_L g6829 ( 
.A(n_6658),
.B(n_957),
.Y(n_6829)
);

NAND2xp5_ASAP7_75t_L g6830 ( 
.A(n_6752),
.B(n_958),
.Y(n_6830)
);

OAI22xp33_ASAP7_75t_R g6831 ( 
.A1(n_6663),
.A2(n_960),
.B1(n_958),
.B2(n_959),
.Y(n_6831)
);

INVx1_ASAP7_75t_L g6832 ( 
.A(n_6768),
.Y(n_6832)
);

NAND2xp5_ASAP7_75t_L g6833 ( 
.A(n_6690),
.B(n_959),
.Y(n_6833)
);

INVx2_ASAP7_75t_L g6834 ( 
.A(n_6713),
.Y(n_6834)
);

HB1xp67_ASAP7_75t_L g6835 ( 
.A(n_6669),
.Y(n_6835)
);

AND2x2_ASAP7_75t_L g6836 ( 
.A(n_6681),
.B(n_961),
.Y(n_6836)
);

OR2x2_ASAP7_75t_L g6837 ( 
.A(n_6638),
.B(n_961),
.Y(n_6837)
);

INVx1_ASAP7_75t_L g6838 ( 
.A(n_6644),
.Y(n_6838)
);

AND2x4_ASAP7_75t_L g6839 ( 
.A(n_6721),
.B(n_963),
.Y(n_6839)
);

NOR2xp33_ASAP7_75t_L g6840 ( 
.A(n_6709),
.B(n_963),
.Y(n_6840)
);

INVx2_ASAP7_75t_L g6841 ( 
.A(n_6687),
.Y(n_6841)
);

NAND2xp5_ASAP7_75t_L g6842 ( 
.A(n_6673),
.B(n_964),
.Y(n_6842)
);

AND2x2_ASAP7_75t_L g6843 ( 
.A(n_6740),
.B(n_964),
.Y(n_6843)
);

NAND2xp5_ASAP7_75t_L g6844 ( 
.A(n_6731),
.B(n_965),
.Y(n_6844)
);

INVx1_ASAP7_75t_L g6845 ( 
.A(n_6726),
.Y(n_6845)
);

INVx2_ASAP7_75t_SL g6846 ( 
.A(n_6689),
.Y(n_6846)
);

OR2x2_ASAP7_75t_L g6847 ( 
.A(n_6664),
.B(n_966),
.Y(n_6847)
);

NAND2xp5_ASAP7_75t_L g6848 ( 
.A(n_6730),
.B(n_967),
.Y(n_6848)
);

AND2x2_ASAP7_75t_L g6849 ( 
.A(n_6728),
.B(n_968),
.Y(n_6849)
);

INVx2_ASAP7_75t_L g6850 ( 
.A(n_6744),
.Y(n_6850)
);

AO21x1_ASAP7_75t_L g6851 ( 
.A1(n_6700),
.A2(n_970),
.B(n_971),
.Y(n_6851)
);

INVx2_ASAP7_75t_L g6852 ( 
.A(n_6707),
.Y(n_6852)
);

OR2x2_ASAP7_75t_L g6853 ( 
.A(n_6653),
.B(n_970),
.Y(n_6853)
);

INVx2_ASAP7_75t_L g6854 ( 
.A(n_6748),
.Y(n_6854)
);

INVx1_ASAP7_75t_L g6855 ( 
.A(n_6729),
.Y(n_6855)
);

NAND2xp5_ASAP7_75t_L g6856 ( 
.A(n_6699),
.B(n_971),
.Y(n_6856)
);

OR2x2_ASAP7_75t_L g6857 ( 
.A(n_6704),
.B(n_972),
.Y(n_6857)
);

AND2x2_ASAP7_75t_L g6858 ( 
.A(n_6695),
.B(n_972),
.Y(n_6858)
);

NAND2x1p5_ASAP7_75t_L g6859 ( 
.A(n_6739),
.B(n_6674),
.Y(n_6859)
);

INVx1_ASAP7_75t_L g6860 ( 
.A(n_6736),
.Y(n_6860)
);

AND2x2_ASAP7_75t_L g6861 ( 
.A(n_6642),
.B(n_973),
.Y(n_6861)
);

NAND2x1p5_ASAP7_75t_L g6862 ( 
.A(n_6650),
.B(n_973),
.Y(n_6862)
);

HB1xp67_ASAP7_75t_L g6863 ( 
.A(n_6734),
.Y(n_6863)
);

AND2x2_ASAP7_75t_L g6864 ( 
.A(n_6652),
.B(n_974),
.Y(n_6864)
);

OR2x2_ASAP7_75t_L g6865 ( 
.A(n_6659),
.B(n_975),
.Y(n_6865)
);

NAND2x1p5_ASAP7_75t_L g6866 ( 
.A(n_6665),
.B(n_976),
.Y(n_6866)
);

INVx1_ASAP7_75t_L g6867 ( 
.A(n_6666),
.Y(n_6867)
);

NAND2xp5_ASAP7_75t_L g6868 ( 
.A(n_6692),
.B(n_976),
.Y(n_6868)
);

INVx1_ASAP7_75t_L g6869 ( 
.A(n_6698),
.Y(n_6869)
);

NAND2xp5_ASAP7_75t_L g6870 ( 
.A(n_6683),
.B(n_977),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_6705),
.Y(n_6871)
);

INVx2_ASAP7_75t_L g6872 ( 
.A(n_6694),
.Y(n_6872)
);

INVx2_ASAP7_75t_L g6873 ( 
.A(n_6715),
.Y(n_6873)
);

INVx2_ASAP7_75t_L g6874 ( 
.A(n_6718),
.Y(n_6874)
);

AND2x2_ASAP7_75t_L g6875 ( 
.A(n_6746),
.B(n_978),
.Y(n_6875)
);

INVx1_ASAP7_75t_L g6876 ( 
.A(n_6719),
.Y(n_6876)
);

AND2x2_ASAP7_75t_L g6877 ( 
.A(n_6733),
.B(n_978),
.Y(n_6877)
);

NAND2xp5_ASAP7_75t_L g6878 ( 
.A(n_6672),
.B(n_979),
.Y(n_6878)
);

NAND2xp5_ASAP7_75t_L g6879 ( 
.A(n_6760),
.B(n_979),
.Y(n_6879)
);

OR2x2_ASAP7_75t_L g6880 ( 
.A(n_6723),
.B(n_980),
.Y(n_6880)
);

INVx1_ASAP7_75t_SL g6881 ( 
.A(n_6735),
.Y(n_6881)
);

NAND2xp5_ASAP7_75t_L g6882 ( 
.A(n_6701),
.B(n_6724),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_6732),
.Y(n_6883)
);

NAND2xp5_ASAP7_75t_L g6884 ( 
.A(n_6737),
.B(n_980),
.Y(n_6884)
);

INVxp67_ASAP7_75t_L g6885 ( 
.A(n_6754),
.Y(n_6885)
);

OR4x1_ASAP7_75t_L g6886 ( 
.A(n_6743),
.B(n_984),
.C(n_982),
.D(n_983),
.Y(n_6886)
);

NAND2xp5_ASAP7_75t_L g6887 ( 
.A(n_6750),
.B(n_982),
.Y(n_6887)
);

OR2x2_ASAP7_75t_L g6888 ( 
.A(n_6751),
.B(n_983),
.Y(n_6888)
);

AND2x2_ASAP7_75t_SL g6889 ( 
.A(n_6678),
.B(n_984),
.Y(n_6889)
);

INVxp67_ASAP7_75t_L g6890 ( 
.A(n_6755),
.Y(n_6890)
);

INVx1_ASAP7_75t_L g6891 ( 
.A(n_6756),
.Y(n_6891)
);

AOI22xp5_ASAP7_75t_L g6892 ( 
.A1(n_6676),
.A2(n_987),
.B1(n_985),
.B2(n_986),
.Y(n_6892)
);

HB1xp67_ASAP7_75t_L g6893 ( 
.A(n_6711),
.Y(n_6893)
);

INVx1_ASAP7_75t_L g6894 ( 
.A(n_6741),
.Y(n_6894)
);

OR2x2_ASAP7_75t_L g6895 ( 
.A(n_6697),
.B(n_986),
.Y(n_6895)
);

INVxp67_ASAP7_75t_L g6896 ( 
.A(n_6722),
.Y(n_6896)
);

HB1xp67_ASAP7_75t_L g6897 ( 
.A(n_6720),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6720),
.Y(n_6898)
);

INVx2_ASAP7_75t_L g6899 ( 
.A(n_6763),
.Y(n_6899)
);

INVx1_ASAP7_75t_L g6900 ( 
.A(n_6720),
.Y(n_6900)
);

AOI22xp5_ASAP7_75t_L g6901 ( 
.A1(n_6812),
.A2(n_989),
.B1(n_987),
.B2(n_988),
.Y(n_6901)
);

OAI21xp5_ASAP7_75t_SL g6902 ( 
.A1(n_6791),
.A2(n_988),
.B(n_990),
.Y(n_6902)
);

AOI21xp33_ASAP7_75t_SL g6903 ( 
.A1(n_6889),
.A2(n_991),
.B(n_992),
.Y(n_6903)
);

HB1xp67_ASAP7_75t_L g6904 ( 
.A(n_6897),
.Y(n_6904)
);

OR2x2_ASAP7_75t_L g6905 ( 
.A(n_6775),
.B(n_991),
.Y(n_6905)
);

INVx1_ASAP7_75t_L g6906 ( 
.A(n_6835),
.Y(n_6906)
);

AOI22xp5_ASAP7_75t_L g6907 ( 
.A1(n_6787),
.A2(n_994),
.B1(n_992),
.B2(n_993),
.Y(n_6907)
);

INVx1_ASAP7_75t_L g6908 ( 
.A(n_6771),
.Y(n_6908)
);

INVx1_ASAP7_75t_L g6909 ( 
.A(n_6898),
.Y(n_6909)
);

OAI22xp5_ASAP7_75t_L g6910 ( 
.A1(n_6892),
.A2(n_996),
.B1(n_994),
.B2(n_995),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_6900),
.Y(n_6911)
);

INVx1_ASAP7_75t_L g6912 ( 
.A(n_6774),
.Y(n_6912)
);

AOI22x1_ASAP7_75t_L g6913 ( 
.A1(n_6770),
.A2(n_997),
.B1(n_995),
.B2(n_996),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_6788),
.Y(n_6914)
);

A2O1A1Ixp33_ASAP7_75t_L g6915 ( 
.A1(n_6826),
.A2(n_1000),
.B(n_998),
.C(n_999),
.Y(n_6915)
);

OAI211xp5_ASAP7_75t_L g6916 ( 
.A1(n_6817),
.A2(n_1000),
.B(n_998),
.C(n_999),
.Y(n_6916)
);

OAI21xp33_ASAP7_75t_L g6917 ( 
.A1(n_6899),
.A2(n_1001),
.B(n_1002),
.Y(n_6917)
);

INVxp67_ASAP7_75t_L g6918 ( 
.A(n_6813),
.Y(n_6918)
);

AOI21xp5_ASAP7_75t_L g6919 ( 
.A1(n_6825),
.A2(n_1001),
.B(n_1002),
.Y(n_6919)
);

OAI21xp5_ASAP7_75t_L g6920 ( 
.A1(n_6781),
.A2(n_6789),
.B(n_6785),
.Y(n_6920)
);

NAND2xp5_ASAP7_75t_L g6921 ( 
.A(n_6821),
.B(n_1003),
.Y(n_6921)
);

OA21x2_ASAP7_75t_L g6922 ( 
.A1(n_6793),
.A2(n_1003),
.B(n_1004),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_6773),
.Y(n_6923)
);

OAI22xp5_ASAP7_75t_SL g6924 ( 
.A1(n_6886),
.A2(n_1006),
.B1(n_1004),
.B2(n_1005),
.Y(n_6924)
);

OA21x2_ASAP7_75t_L g6925 ( 
.A1(n_6878),
.A2(n_1006),
.B(n_1007),
.Y(n_6925)
);

AOI21xp33_ASAP7_75t_L g6926 ( 
.A1(n_6811),
.A2(n_1007),
.B(n_1008),
.Y(n_6926)
);

INVx1_ASAP7_75t_L g6927 ( 
.A(n_6802),
.Y(n_6927)
);

HB1xp67_ASAP7_75t_L g6928 ( 
.A(n_6862),
.Y(n_6928)
);

NOR3xp33_ASAP7_75t_L g6929 ( 
.A(n_6772),
.B(n_1009),
.C(n_1010),
.Y(n_6929)
);

INVx2_ASAP7_75t_L g6930 ( 
.A(n_6795),
.Y(n_6930)
);

AO21x1_ASAP7_75t_L g6931 ( 
.A1(n_6786),
.A2(n_1012),
.B(n_1011),
.Y(n_6931)
);

OAI22xp33_ASAP7_75t_L g6932 ( 
.A1(n_6780),
.A2(n_1012),
.B1(n_1009),
.B2(n_1011),
.Y(n_6932)
);

XNOR2xp5_ASAP7_75t_L g6933 ( 
.A(n_6805),
.B(n_6893),
.Y(n_6933)
);

OAI21xp5_ASAP7_75t_L g6934 ( 
.A1(n_6806),
.A2(n_6808),
.B(n_6815),
.Y(n_6934)
);

AOI21xp5_ASAP7_75t_L g6935 ( 
.A1(n_6810),
.A2(n_1013),
.B(n_1014),
.Y(n_6935)
);

NAND2xp5_ASAP7_75t_L g6936 ( 
.A(n_6894),
.B(n_1013),
.Y(n_6936)
);

XNOR2xp5_ASAP7_75t_L g6937 ( 
.A(n_6881),
.B(n_1014),
.Y(n_6937)
);

AOI22xp33_ASAP7_75t_L g6938 ( 
.A1(n_6863),
.A2(n_1017),
.B1(n_1015),
.B2(n_1016),
.Y(n_6938)
);

OAI22xp5_ASAP7_75t_L g6939 ( 
.A1(n_6885),
.A2(n_1019),
.B1(n_1015),
.B2(n_1018),
.Y(n_6939)
);

AOI22xp5_ASAP7_75t_L g6940 ( 
.A1(n_6890),
.A2(n_1021),
.B1(n_1018),
.B2(n_1019),
.Y(n_6940)
);

AOI21xp5_ASAP7_75t_L g6941 ( 
.A1(n_6818),
.A2(n_1022),
.B(n_1023),
.Y(n_6941)
);

AND2x2_ASAP7_75t_L g6942 ( 
.A(n_6784),
.B(n_1022),
.Y(n_6942)
);

INVx2_ASAP7_75t_L g6943 ( 
.A(n_6859),
.Y(n_6943)
);

OAI22xp5_ASAP7_75t_L g6944 ( 
.A1(n_6896),
.A2(n_1025),
.B1(n_1023),
.B2(n_1024),
.Y(n_6944)
);

AOI21xp33_ASAP7_75t_L g6945 ( 
.A1(n_6838),
.A2(n_6832),
.B(n_6794),
.Y(n_6945)
);

AOI22xp5_ASAP7_75t_L g6946 ( 
.A1(n_6872),
.A2(n_1026),
.B1(n_1024),
.B2(n_1025),
.Y(n_6946)
);

OAI221xp5_ASAP7_75t_L g6947 ( 
.A1(n_6882),
.A2(n_1031),
.B1(n_1027),
.B2(n_1030),
.C(n_1032),
.Y(n_6947)
);

INVx2_ASAP7_75t_L g6948 ( 
.A(n_6866),
.Y(n_6948)
);

INVx2_ASAP7_75t_L g6949 ( 
.A(n_6769),
.Y(n_6949)
);

AND2x2_ASAP7_75t_L g6950 ( 
.A(n_6800),
.B(n_1031),
.Y(n_6950)
);

INVx1_ASAP7_75t_L g6951 ( 
.A(n_6836),
.Y(n_6951)
);

AND2x2_ASAP7_75t_L g6952 ( 
.A(n_6804),
.B(n_1032),
.Y(n_6952)
);

AND2x2_ASAP7_75t_L g6953 ( 
.A(n_6834),
.B(n_6850),
.Y(n_6953)
);

INVx2_ASAP7_75t_SL g6954 ( 
.A(n_6776),
.Y(n_6954)
);

AOI22xp33_ASAP7_75t_SL g6955 ( 
.A1(n_6782),
.A2(n_1035),
.B1(n_1033),
.B2(n_1034),
.Y(n_6955)
);

AOI211xp5_ASAP7_75t_SL g6956 ( 
.A1(n_6777),
.A2(n_1037),
.B(n_1035),
.C(n_1036),
.Y(n_6956)
);

NAND4xp25_ASAP7_75t_SL g6957 ( 
.A(n_6851),
.B(n_1040),
.C(n_1038),
.D(n_1039),
.Y(n_6957)
);

NAND2xp5_ASAP7_75t_L g6958 ( 
.A(n_6846),
.B(n_6792),
.Y(n_6958)
);

OAI22xp33_ASAP7_75t_L g6959 ( 
.A1(n_6790),
.A2(n_1040),
.B1(n_1038),
.B2(n_1039),
.Y(n_6959)
);

INVx2_ASAP7_75t_L g6960 ( 
.A(n_6809),
.Y(n_6960)
);

INVx1_ASAP7_75t_L g6961 ( 
.A(n_6849),
.Y(n_6961)
);

INVx2_ASAP7_75t_SL g6962 ( 
.A(n_6803),
.Y(n_6962)
);

INVxp67_ASAP7_75t_L g6963 ( 
.A(n_6801),
.Y(n_6963)
);

INVx1_ASAP7_75t_L g6964 ( 
.A(n_6816),
.Y(n_6964)
);

INVx1_ASAP7_75t_L g6965 ( 
.A(n_6779),
.Y(n_6965)
);

OAI21xp33_ASAP7_75t_L g6966 ( 
.A1(n_6783),
.A2(n_1041),
.B(n_1042),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6843),
.Y(n_6967)
);

AOI22xp33_ASAP7_75t_SL g6968 ( 
.A1(n_6824),
.A2(n_1045),
.B1(n_1043),
.B2(n_1044),
.Y(n_6968)
);

AOI22xp5_ASAP7_75t_L g6969 ( 
.A1(n_6831),
.A2(n_1045),
.B1(n_1043),
.B2(n_1044),
.Y(n_6969)
);

INVx1_ASAP7_75t_SL g6970 ( 
.A(n_6828),
.Y(n_6970)
);

OAI21xp33_ASAP7_75t_SL g6971 ( 
.A1(n_6819),
.A2(n_1046),
.B(n_1047),
.Y(n_6971)
);

NAND2xp5_ASAP7_75t_L g6972 ( 
.A(n_6839),
.B(n_1046),
.Y(n_6972)
);

NAND3xp33_ASAP7_75t_L g6973 ( 
.A(n_6798),
.B(n_1048),
.C(n_1049),
.Y(n_6973)
);

OAI22xp5_ASAP7_75t_L g6974 ( 
.A1(n_6823),
.A2(n_1051),
.B1(n_1048),
.B2(n_1050),
.Y(n_6974)
);

AOI21xp33_ASAP7_75t_L g6975 ( 
.A1(n_6845),
.A2(n_6860),
.B(n_6855),
.Y(n_6975)
);

INVx2_ASAP7_75t_L g6976 ( 
.A(n_6797),
.Y(n_6976)
);

INVx2_ASAP7_75t_SL g6977 ( 
.A(n_6822),
.Y(n_6977)
);

NAND4xp25_ASAP7_75t_L g6978 ( 
.A(n_6807),
.B(n_1052),
.C(n_1050),
.D(n_1051),
.Y(n_6978)
);

OAI21xp33_ASAP7_75t_SL g6979 ( 
.A1(n_6814),
.A2(n_1053),
.B(n_1054),
.Y(n_6979)
);

OR2x2_ASAP7_75t_L g6980 ( 
.A(n_6829),
.B(n_1053),
.Y(n_6980)
);

INVx1_ASAP7_75t_SL g6981 ( 
.A(n_6895),
.Y(n_6981)
);

AOI22xp5_ASAP7_75t_L g6982 ( 
.A1(n_6841),
.A2(n_1056),
.B1(n_1054),
.B2(n_1055),
.Y(n_6982)
);

INVx1_ASAP7_75t_L g6983 ( 
.A(n_6827),
.Y(n_6983)
);

AOI21xp33_ASAP7_75t_L g6984 ( 
.A1(n_6869),
.A2(n_1055),
.B(n_1056),
.Y(n_6984)
);

INVx1_ASAP7_75t_SL g6985 ( 
.A(n_6875),
.Y(n_6985)
);

INVx1_ASAP7_75t_L g6986 ( 
.A(n_6830),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_6857),
.Y(n_6987)
);

OR2x2_ASAP7_75t_L g6988 ( 
.A(n_6837),
.B(n_1057),
.Y(n_6988)
);

INVx1_ASAP7_75t_L g6989 ( 
.A(n_6858),
.Y(n_6989)
);

INVxp67_ASAP7_75t_L g6990 ( 
.A(n_6844),
.Y(n_6990)
);

AOI22xp5_ASAP7_75t_L g6991 ( 
.A1(n_6852),
.A2(n_1060),
.B1(n_1057),
.B2(n_1058),
.Y(n_6991)
);

NAND4xp25_ASAP7_75t_SL g6992 ( 
.A(n_6879),
.B(n_1065),
.C(n_1061),
.D(n_1062),
.Y(n_6992)
);

INVxp67_ASAP7_75t_L g6993 ( 
.A(n_6778),
.Y(n_6993)
);

INVx1_ASAP7_75t_L g6994 ( 
.A(n_6880),
.Y(n_6994)
);

XOR2x2_ASAP7_75t_L g6995 ( 
.A(n_6870),
.B(n_1061),
.Y(n_6995)
);

OAI21xp33_ASAP7_75t_L g6996 ( 
.A1(n_6854),
.A2(n_1062),
.B(n_1065),
.Y(n_6996)
);

INVx1_ASAP7_75t_SL g6997 ( 
.A(n_6877),
.Y(n_6997)
);

NAND4xp75_ASAP7_75t_L g6998 ( 
.A(n_6867),
.B(n_1068),
.C(n_1066),
.D(n_1067),
.Y(n_6998)
);

OAI21xp33_ASAP7_75t_L g6999 ( 
.A1(n_6891),
.A2(n_1068),
.B(n_1069),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6888),
.Y(n_7000)
);

INVx2_ASAP7_75t_SL g7001 ( 
.A(n_6861),
.Y(n_7001)
);

XOR2xp5_ASAP7_75t_L g7002 ( 
.A(n_6847),
.B(n_1070),
.Y(n_7002)
);

INVx3_ASAP7_75t_L g7003 ( 
.A(n_6873),
.Y(n_7003)
);

A2O1A1Ixp33_ASAP7_75t_L g7004 ( 
.A1(n_6856),
.A2(n_1072),
.B(n_1070),
.C(n_1071),
.Y(n_7004)
);

OAI21xp33_ASAP7_75t_SL g7005 ( 
.A1(n_6871),
.A2(n_1072),
.B(n_1073),
.Y(n_7005)
);

AND2x4_ASAP7_75t_L g7006 ( 
.A(n_6874),
.B(n_1074),
.Y(n_7006)
);

INVx1_ASAP7_75t_L g7007 ( 
.A(n_6796),
.Y(n_7007)
);

INVx1_ASAP7_75t_L g7008 ( 
.A(n_6864),
.Y(n_7008)
);

BUFx2_ASAP7_75t_L g7009 ( 
.A(n_6799),
.Y(n_7009)
);

INVx1_ASAP7_75t_L g7010 ( 
.A(n_6865),
.Y(n_7010)
);

INVx2_ASAP7_75t_L g7011 ( 
.A(n_6853),
.Y(n_7011)
);

AOI22xp5_ASAP7_75t_L g7012 ( 
.A1(n_6840),
.A2(n_1076),
.B1(n_1074),
.B2(n_1075),
.Y(n_7012)
);

NAND3xp33_ASAP7_75t_L g7013 ( 
.A(n_6876),
.B(n_1075),
.C(n_1077),
.Y(n_7013)
);

INVx1_ASAP7_75t_L g7014 ( 
.A(n_6820),
.Y(n_7014)
);

INVx1_ASAP7_75t_L g7015 ( 
.A(n_6842),
.Y(n_7015)
);

AOI22xp5_ASAP7_75t_L g7016 ( 
.A1(n_6883),
.A2(n_1079),
.B1(n_1077),
.B2(n_1078),
.Y(n_7016)
);

NAND2xp5_ASAP7_75t_L g7017 ( 
.A(n_6868),
.B(n_1078),
.Y(n_7017)
);

INVx2_ASAP7_75t_L g7018 ( 
.A(n_6884),
.Y(n_7018)
);

INVx1_ASAP7_75t_L g7019 ( 
.A(n_6887),
.Y(n_7019)
);

INVxp67_ASAP7_75t_L g7020 ( 
.A(n_6833),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6848),
.Y(n_7021)
);

AOI22xp33_ASAP7_75t_L g7022 ( 
.A1(n_6889),
.A2(n_1081),
.B1(n_1079),
.B2(n_1080),
.Y(n_7022)
);

NAND2xp5_ASAP7_75t_L g7023 ( 
.A(n_6812),
.B(n_1081),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6897),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6897),
.Y(n_7025)
);

OAI21xp33_ASAP7_75t_L g7026 ( 
.A1(n_6787),
.A2(n_1082),
.B(n_1083),
.Y(n_7026)
);

OAI22xp33_ASAP7_75t_L g7027 ( 
.A1(n_6787),
.A2(n_1084),
.B1(n_1082),
.B2(n_1083),
.Y(n_7027)
);

XOR2x2_ASAP7_75t_L g7028 ( 
.A(n_6889),
.B(n_1084),
.Y(n_7028)
);

INVxp67_ASAP7_75t_L g7029 ( 
.A(n_6897),
.Y(n_7029)
);

INVx2_ASAP7_75t_L g7030 ( 
.A(n_6795),
.Y(n_7030)
);

OAI221xp5_ASAP7_75t_SL g7031 ( 
.A1(n_6826),
.A2(n_1101),
.B1(n_1109),
.B2(n_1093),
.C(n_1085),
.Y(n_7031)
);

INVx1_ASAP7_75t_SL g7032 ( 
.A(n_6770),
.Y(n_7032)
);

OAI22xp33_ASAP7_75t_L g7033 ( 
.A1(n_6787),
.A2(n_1087),
.B1(n_1085),
.B2(n_1086),
.Y(n_7033)
);

OAI21xp5_ASAP7_75t_L g7034 ( 
.A1(n_6826),
.A2(n_1087),
.B(n_1088),
.Y(n_7034)
);

INVx2_ASAP7_75t_L g7035 ( 
.A(n_6795),
.Y(n_7035)
);

OAI22xp5_ASAP7_75t_L g7036 ( 
.A1(n_6787),
.A2(n_1090),
.B1(n_1088),
.B2(n_1089),
.Y(n_7036)
);

OA22x2_ASAP7_75t_L g7037 ( 
.A1(n_6791),
.A2(n_1092),
.B1(n_1089),
.B2(n_1091),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6897),
.Y(n_7038)
);

OAI21xp33_ASAP7_75t_L g7039 ( 
.A1(n_6787),
.A2(n_1091),
.B(n_1092),
.Y(n_7039)
);

AND2x2_ASAP7_75t_L g7040 ( 
.A(n_6821),
.B(n_1093),
.Y(n_7040)
);

INVx1_ASAP7_75t_L g7041 ( 
.A(n_6897),
.Y(n_7041)
);

AOI22xp5_ASAP7_75t_L g7042 ( 
.A1(n_6812),
.A2(n_1096),
.B1(n_1094),
.B2(n_1095),
.Y(n_7042)
);

AOI21xp5_ASAP7_75t_L g7043 ( 
.A1(n_6787),
.A2(n_1094),
.B(n_1095),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_6897),
.Y(n_7044)
);

NAND2xp5_ASAP7_75t_L g7045 ( 
.A(n_6812),
.B(n_1097),
.Y(n_7045)
);

XNOR2xp5_ASAP7_75t_L g7046 ( 
.A(n_6892),
.B(n_1097),
.Y(n_7046)
);

XNOR2x1_ASAP7_75t_L g7047 ( 
.A(n_6892),
.B(n_1098),
.Y(n_7047)
);

NAND2xp5_ASAP7_75t_L g7048 ( 
.A(n_6812),
.B(n_1099),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_6897),
.Y(n_7049)
);

XOR2xp5_ASAP7_75t_L g7050 ( 
.A(n_6892),
.B(n_1100),
.Y(n_7050)
);

XOR2x2_ASAP7_75t_L g7051 ( 
.A(n_6889),
.B(n_1100),
.Y(n_7051)
);

AOI22xp5_ASAP7_75t_L g7052 ( 
.A1(n_6812),
.A2(n_1103),
.B1(n_1101),
.B2(n_1102),
.Y(n_7052)
);

OAI22xp5_ASAP7_75t_L g7053 ( 
.A1(n_6787),
.A2(n_1105),
.B1(n_1102),
.B2(n_1104),
.Y(n_7053)
);

INVx1_ASAP7_75t_L g7054 ( 
.A(n_6897),
.Y(n_7054)
);

INVx2_ASAP7_75t_L g7055 ( 
.A(n_6795),
.Y(n_7055)
);

AO22x1_ASAP7_75t_L g7056 ( 
.A1(n_6812),
.A2(n_1108),
.B1(n_1106),
.B2(n_1107),
.Y(n_7056)
);

AO22x1_ASAP7_75t_L g7057 ( 
.A1(n_6812),
.A2(n_1111),
.B1(n_1109),
.B2(n_1110),
.Y(n_7057)
);

AOI22xp5_ASAP7_75t_L g7058 ( 
.A1(n_6812),
.A2(n_1113),
.B1(n_1110),
.B2(n_1111),
.Y(n_7058)
);

AOI221xp5_ASAP7_75t_L g7059 ( 
.A1(n_6812),
.A2(n_1130),
.B1(n_1138),
.B2(n_1122),
.C(n_1114),
.Y(n_7059)
);

OAI21xp5_ASAP7_75t_L g7060 ( 
.A1(n_6826),
.A2(n_1115),
.B(n_1116),
.Y(n_7060)
);

INVx1_ASAP7_75t_L g7061 ( 
.A(n_6897),
.Y(n_7061)
);

AND2x2_ASAP7_75t_L g7062 ( 
.A(n_6821),
.B(n_1115),
.Y(n_7062)
);

INVx1_ASAP7_75t_L g7063 ( 
.A(n_6897),
.Y(n_7063)
);

INVx1_ASAP7_75t_L g7064 ( 
.A(n_6897),
.Y(n_7064)
);

AOI21xp33_ASAP7_75t_SL g7065 ( 
.A1(n_6889),
.A2(n_1116),
.B(n_1117),
.Y(n_7065)
);

OAI211xp5_ASAP7_75t_L g7066 ( 
.A1(n_6812),
.A2(n_1119),
.B(n_1117),
.C(n_1118),
.Y(n_7066)
);

OAI21xp33_ASAP7_75t_SL g7067 ( 
.A1(n_6812),
.A2(n_1120),
.B(n_1121),
.Y(n_7067)
);

NAND2xp5_ASAP7_75t_L g7068 ( 
.A(n_6812),
.B(n_1121),
.Y(n_7068)
);

XNOR2x1_ASAP7_75t_L g7069 ( 
.A(n_6892),
.B(n_1122),
.Y(n_7069)
);

NAND2xp5_ASAP7_75t_L g7070 ( 
.A(n_6812),
.B(n_1123),
.Y(n_7070)
);

INVx1_ASAP7_75t_L g7071 ( 
.A(n_6897),
.Y(n_7071)
);

INVx2_ASAP7_75t_L g7072 ( 
.A(n_6795),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_6897),
.Y(n_7073)
);

INVx3_ASAP7_75t_L g7074 ( 
.A(n_6795),
.Y(n_7074)
);

OAI22xp5_ASAP7_75t_L g7075 ( 
.A1(n_6787),
.A2(n_1126),
.B1(n_1124),
.B2(n_1125),
.Y(n_7075)
);

AOI211xp5_ASAP7_75t_SL g7076 ( 
.A1(n_6812),
.A2(n_1128),
.B(n_1126),
.C(n_1127),
.Y(n_7076)
);

INVx1_ASAP7_75t_L g7077 ( 
.A(n_6897),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_6897),
.Y(n_7078)
);

OAI211xp5_ASAP7_75t_L g7079 ( 
.A1(n_6812),
.A2(n_1129),
.B(n_1127),
.C(n_1128),
.Y(n_7079)
);

AOI22xp33_ASAP7_75t_L g7080 ( 
.A1(n_6889),
.A2(n_1132),
.B1(n_1130),
.B2(n_1131),
.Y(n_7080)
);

OAI22xp5_ASAP7_75t_L g7081 ( 
.A1(n_6787),
.A2(n_1134),
.B1(n_1131),
.B2(n_1133),
.Y(n_7081)
);

AOI21xp33_ASAP7_75t_SL g7082 ( 
.A1(n_6889),
.A2(n_1133),
.B(n_1134),
.Y(n_7082)
);

AOI22xp33_ASAP7_75t_L g7083 ( 
.A1(n_6889),
.A2(n_1137),
.B1(n_1135),
.B2(n_1136),
.Y(n_7083)
);

AOI22xp5_ASAP7_75t_L g7084 ( 
.A1(n_6812),
.A2(n_1137),
.B1(n_1135),
.B2(n_1136),
.Y(n_7084)
);

INVx2_ASAP7_75t_SL g7085 ( 
.A(n_6897),
.Y(n_7085)
);

O2A1O1Ixp33_ASAP7_75t_L g7086 ( 
.A1(n_6812),
.A2(n_1141),
.B(n_1139),
.C(n_1140),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_6897),
.Y(n_7087)
);

OAI21xp33_ASAP7_75t_L g7088 ( 
.A1(n_6787),
.A2(n_1140),
.B(n_1141),
.Y(n_7088)
);

INVx2_ASAP7_75t_L g7089 ( 
.A(n_6795),
.Y(n_7089)
);

NOR3xp33_ASAP7_75t_L g7090 ( 
.A(n_6787),
.B(n_1142),
.C(n_1143),
.Y(n_7090)
);

XOR2xp5_ASAP7_75t_L g7091 ( 
.A(n_6892),
.B(n_1144),
.Y(n_7091)
);

OA21x2_ASAP7_75t_L g7092 ( 
.A1(n_6812),
.A2(n_1144),
.B(n_1145),
.Y(n_7092)
);

NAND3xp33_ASAP7_75t_L g7093 ( 
.A(n_7076),
.B(n_1147),
.C(n_1148),
.Y(n_7093)
);

OAI211xp5_ASAP7_75t_L g7094 ( 
.A1(n_7067),
.A2(n_1149),
.B(n_1147),
.C(n_1148),
.Y(n_7094)
);

INVx1_ASAP7_75t_SL g7095 ( 
.A(n_7032),
.Y(n_7095)
);

INVx1_ASAP7_75t_L g7096 ( 
.A(n_6904),
.Y(n_7096)
);

INVx2_ASAP7_75t_L g7097 ( 
.A(n_7074),
.Y(n_7097)
);

INVx1_ASAP7_75t_SL g7098 ( 
.A(n_7040),
.Y(n_7098)
);

NOR2xp33_ASAP7_75t_L g7099 ( 
.A(n_6918),
.B(n_1150),
.Y(n_7099)
);

OR2x2_ASAP7_75t_L g7100 ( 
.A(n_6981),
.B(n_1151),
.Y(n_7100)
);

INVx1_ASAP7_75t_L g7101 ( 
.A(n_7062),
.Y(n_7101)
);

NAND2xp5_ASAP7_75t_L g7102 ( 
.A(n_7056),
.B(n_1151),
.Y(n_7102)
);

INVx1_ASAP7_75t_L g7103 ( 
.A(n_6921),
.Y(n_7103)
);

OAI21xp33_ASAP7_75t_L g7104 ( 
.A1(n_6933),
.A2(n_1152),
.B(n_1153),
.Y(n_7104)
);

OAI21xp33_ASAP7_75t_L g7105 ( 
.A1(n_6934),
.A2(n_1152),
.B(n_1154),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_7085),
.Y(n_7106)
);

INVx3_ASAP7_75t_L g7107 ( 
.A(n_6930),
.Y(n_7107)
);

INVxp67_ASAP7_75t_L g7108 ( 
.A(n_7092),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6953),
.Y(n_7109)
);

NAND2xp5_ASAP7_75t_L g7110 ( 
.A(n_7057),
.B(n_1155),
.Y(n_7110)
);

AND2x2_ASAP7_75t_L g7111 ( 
.A(n_7030),
.B(n_1156),
.Y(n_7111)
);

NAND2xp5_ASAP7_75t_L g7112 ( 
.A(n_6955),
.B(n_1156),
.Y(n_7112)
);

OR2x6_ASAP7_75t_L g7113 ( 
.A(n_6954),
.B(n_1157),
.Y(n_7113)
);

OAI21xp33_ASAP7_75t_SL g7114 ( 
.A1(n_7023),
.A2(n_1158),
.B(n_1159),
.Y(n_7114)
);

AOI21xp5_ASAP7_75t_L g7115 ( 
.A1(n_7045),
.A2(n_1158),
.B(n_1160),
.Y(n_7115)
);

NAND3xp33_ASAP7_75t_L g7116 ( 
.A(n_7092),
.B(n_1161),
.C(n_1162),
.Y(n_7116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g7117 ( 
.A1(n_6915),
.A2(n_1181),
.B(n_1190),
.C(n_1172),
.D(n_1162),
.Y(n_7117)
);

NOR3xp33_ASAP7_75t_SL g7118 ( 
.A(n_6945),
.B(n_1163),
.C(n_1164),
.Y(n_7118)
);

AOI21xp5_ASAP7_75t_L g7119 ( 
.A1(n_7048),
.A2(n_1165),
.B(n_1166),
.Y(n_7119)
);

OAI211xp5_ASAP7_75t_L g7120 ( 
.A1(n_7068),
.A2(n_1167),
.B(n_1165),
.C(n_1166),
.Y(n_7120)
);

OR2x6_ASAP7_75t_L g7121 ( 
.A(n_6943),
.B(n_7029),
.Y(n_7121)
);

OAI21xp33_ASAP7_75t_SL g7122 ( 
.A1(n_7070),
.A2(n_1167),
.B(n_1168),
.Y(n_7122)
);

NAND2xp5_ASAP7_75t_L g7123 ( 
.A(n_7035),
.B(n_1168),
.Y(n_7123)
);

AOI21xp5_ASAP7_75t_L g7124 ( 
.A1(n_7086),
.A2(n_1171),
.B(n_1173),
.Y(n_7124)
);

INVx1_ASAP7_75t_L g7125 ( 
.A(n_6950),
.Y(n_7125)
);

INVxp67_ASAP7_75t_L g7126 ( 
.A(n_6928),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_7024),
.Y(n_7127)
);

NOR2xp33_ASAP7_75t_L g7128 ( 
.A(n_6903),
.B(n_1171),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_7025),
.Y(n_7129)
);

INVx2_ASAP7_75t_L g7130 ( 
.A(n_7055),
.Y(n_7130)
);

OAI22xp5_ASAP7_75t_L g7131 ( 
.A1(n_7031),
.A2(n_1176),
.B1(n_1173),
.B2(n_1174),
.Y(n_7131)
);

OR2x2_ASAP7_75t_L g7132 ( 
.A(n_6985),
.B(n_1174),
.Y(n_7132)
);

NAND2xp5_ASAP7_75t_L g7133 ( 
.A(n_7072),
.B(n_1176),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_7038),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_7041),
.Y(n_7135)
);

NAND2xp5_ASAP7_75t_L g7136 ( 
.A(n_7089),
.B(n_1177),
.Y(n_7136)
);

AOI221xp5_ASAP7_75t_L g7137 ( 
.A1(n_6920),
.A2(n_1179),
.B1(n_1177),
.B2(n_1178),
.C(n_1180),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_7044),
.Y(n_7138)
);

INVx1_ASAP7_75t_L g7139 ( 
.A(n_7049),
.Y(n_7139)
);

AND2x4_ASAP7_75t_L g7140 ( 
.A(n_6962),
.B(n_1178),
.Y(n_7140)
);

AND2x2_ASAP7_75t_L g7141 ( 
.A(n_6997),
.B(n_1179),
.Y(n_7141)
);

INVx1_ASAP7_75t_L g7142 ( 
.A(n_7054),
.Y(n_7142)
);

INVx1_ASAP7_75t_L g7143 ( 
.A(n_7061),
.Y(n_7143)
);

INVx1_ASAP7_75t_L g7144 ( 
.A(n_7063),
.Y(n_7144)
);

AOI21xp5_ASAP7_75t_L g7145 ( 
.A1(n_7028),
.A2(n_1180),
.B(n_1181),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_7064),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_7071),
.Y(n_7147)
);

AND2x2_ASAP7_75t_L g7148 ( 
.A(n_6948),
.B(n_1182),
.Y(n_7148)
);

INVx1_ASAP7_75t_L g7149 ( 
.A(n_7073),
.Y(n_7149)
);

INVxp67_ASAP7_75t_L g7150 ( 
.A(n_6957),
.Y(n_7150)
);

INVx3_ASAP7_75t_L g7151 ( 
.A(n_7003),
.Y(n_7151)
);

OAI21xp33_ASAP7_75t_L g7152 ( 
.A1(n_6958),
.A2(n_1182),
.B(n_1183),
.Y(n_7152)
);

OAI22xp5_ASAP7_75t_L g7153 ( 
.A1(n_7022),
.A2(n_1186),
.B1(n_1183),
.B2(n_1185),
.Y(n_7153)
);

INVx1_ASAP7_75t_L g7154 ( 
.A(n_7077),
.Y(n_7154)
);

INVx1_ASAP7_75t_L g7155 ( 
.A(n_7078),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_7087),
.Y(n_7156)
);

OAI21xp5_ASAP7_75t_SL g7157 ( 
.A1(n_7034),
.A2(n_1185),
.B(n_1186),
.Y(n_7157)
);

O2A1O1Ixp33_ASAP7_75t_L g7158 ( 
.A1(n_7065),
.A2(n_1189),
.B(n_1187),
.C(n_1188),
.Y(n_7158)
);

AOI22xp5_ASAP7_75t_L g7159 ( 
.A1(n_6924),
.A2(n_1189),
.B1(n_1187),
.B2(n_1188),
.Y(n_7159)
);

NAND2xp5_ASAP7_75t_L g7160 ( 
.A(n_7082),
.B(n_1191),
.Y(n_7160)
);

NAND2xp5_ASAP7_75t_L g7161 ( 
.A(n_6956),
.B(n_7080),
.Y(n_7161)
);

AND2x2_ASAP7_75t_L g7162 ( 
.A(n_6949),
.B(n_1191),
.Y(n_7162)
);

OR2x2_ASAP7_75t_L g7163 ( 
.A(n_7001),
.B(n_1192),
.Y(n_7163)
);

NAND2xp5_ASAP7_75t_L g7164 ( 
.A(n_7083),
.B(n_1192),
.Y(n_7164)
);

AND2x2_ASAP7_75t_L g7165 ( 
.A(n_6976),
.B(n_1193),
.Y(n_7165)
);

OAI211xp5_ASAP7_75t_L g7166 ( 
.A1(n_7066),
.A2(n_7079),
.B(n_7060),
.C(n_7042),
.Y(n_7166)
);

INVx1_ASAP7_75t_L g7167 ( 
.A(n_6952),
.Y(n_7167)
);

INVx2_ASAP7_75t_L g7168 ( 
.A(n_6980),
.Y(n_7168)
);

OAI22xp5_ASAP7_75t_L g7169 ( 
.A1(n_6901),
.A2(n_1195),
.B1(n_1193),
.B2(n_1194),
.Y(n_7169)
);

INVx2_ASAP7_75t_L g7170 ( 
.A(n_6905),
.Y(n_7170)
);

INVx3_ASAP7_75t_L g7171 ( 
.A(n_6960),
.Y(n_7171)
);

AND2x2_ASAP7_75t_L g7172 ( 
.A(n_6927),
.B(n_1194),
.Y(n_7172)
);

NAND2xp5_ASAP7_75t_L g7173 ( 
.A(n_6969),
.B(n_1196),
.Y(n_7173)
);

NAND2xp5_ASAP7_75t_L g7174 ( 
.A(n_6935),
.B(n_1196),
.Y(n_7174)
);

NAND2xp5_ASAP7_75t_L g7175 ( 
.A(n_7052),
.B(n_1197),
.Y(n_7175)
);

INVx1_ASAP7_75t_L g7176 ( 
.A(n_6936),
.Y(n_7176)
);

INVxp67_ASAP7_75t_SL g7177 ( 
.A(n_6931),
.Y(n_7177)
);

INVx2_ASAP7_75t_L g7178 ( 
.A(n_7006),
.Y(n_7178)
);

AND2x4_ASAP7_75t_L g7179 ( 
.A(n_6977),
.B(n_1197),
.Y(n_7179)
);

INVx1_ASAP7_75t_L g7180 ( 
.A(n_6906),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_6988),
.Y(n_7181)
);

NAND2xp5_ASAP7_75t_L g7182 ( 
.A(n_7058),
.B(n_1198),
.Y(n_7182)
);

OAI22xp33_ASAP7_75t_SL g7183 ( 
.A1(n_6908),
.A2(n_1201),
.B1(n_1198),
.B2(n_1199),
.Y(n_7183)
);

INVx1_ASAP7_75t_L g7184 ( 
.A(n_6942),
.Y(n_7184)
);

AOI22xp5_ASAP7_75t_L g7185 ( 
.A1(n_7090),
.A2(n_1202),
.B1(n_1199),
.B2(n_1201),
.Y(n_7185)
);

INVx2_ASAP7_75t_L g7186 ( 
.A(n_7006),
.Y(n_7186)
);

AOI21xp5_ASAP7_75t_L g7187 ( 
.A1(n_7051),
.A2(n_1202),
.B(n_1203),
.Y(n_7187)
);

OR2x2_ASAP7_75t_L g7188 ( 
.A(n_6970),
.B(n_1203),
.Y(n_7188)
);

NAND2xp5_ASAP7_75t_SL g7189 ( 
.A(n_6971),
.B(n_6979),
.Y(n_7189)
);

OAI32xp33_ASAP7_75t_L g7190 ( 
.A1(n_7005),
.A2(n_1221),
.A3(n_1230),
.B1(n_1212),
.B2(n_1204),
.Y(n_7190)
);

INVx1_ASAP7_75t_L g7191 ( 
.A(n_6972),
.Y(n_7191)
);

INVx1_ASAP7_75t_L g7192 ( 
.A(n_6951),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_6964),
.Y(n_7193)
);

AOI22xp5_ASAP7_75t_L g7194 ( 
.A1(n_7084),
.A2(n_1206),
.B1(n_1204),
.B2(n_1205),
.Y(n_7194)
);

INVx1_ASAP7_75t_L g7195 ( 
.A(n_6989),
.Y(n_7195)
);

HB1xp67_ASAP7_75t_L g7196 ( 
.A(n_6925),
.Y(n_7196)
);

NAND2xp5_ASAP7_75t_L g7197 ( 
.A(n_7043),
.B(n_1205),
.Y(n_7197)
);

INVx1_ASAP7_75t_L g7198 ( 
.A(n_7008),
.Y(n_7198)
);

AOI33xp33_ASAP7_75t_L g7199 ( 
.A1(n_6912),
.A2(n_1208),
.A3(n_1210),
.B1(n_1206),
.B2(n_1207),
.B3(n_1209),
.Y(n_7199)
);

AOI22xp33_ASAP7_75t_L g7200 ( 
.A1(n_6961),
.A2(n_1210),
.B1(n_1207),
.B2(n_1208),
.Y(n_7200)
);

INVx1_ASAP7_75t_L g7201 ( 
.A(n_6967),
.Y(n_7201)
);

OR2x2_ASAP7_75t_L g7202 ( 
.A(n_6914),
.B(n_1211),
.Y(n_7202)
);

INVx2_ASAP7_75t_L g7203 ( 
.A(n_7011),
.Y(n_7203)
);

OR2x2_ASAP7_75t_L g7204 ( 
.A(n_6909),
.B(n_1211),
.Y(n_7204)
);

AOI22xp33_ASAP7_75t_L g7205 ( 
.A1(n_7021),
.A2(n_1215),
.B1(n_1213),
.B2(n_1214),
.Y(n_7205)
);

NOR3xp33_ASAP7_75t_L g7206 ( 
.A(n_6975),
.B(n_6990),
.C(n_6963),
.Y(n_7206)
);

AOI32xp33_ASAP7_75t_L g7207 ( 
.A1(n_7059),
.A2(n_1216),
.A3(n_1213),
.B1(n_1214),
.B2(n_1217),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_6937),
.Y(n_7208)
);

INVx1_ASAP7_75t_L g7209 ( 
.A(n_6911),
.Y(n_7209)
);

AOI22xp5_ASAP7_75t_L g7210 ( 
.A1(n_7026),
.A2(n_1218),
.B1(n_1216),
.B2(n_1217),
.Y(n_7210)
);

INVx1_ASAP7_75t_L g7211 ( 
.A(n_7002),
.Y(n_7211)
);

AOI21xp33_ASAP7_75t_SL g7212 ( 
.A1(n_6932),
.A2(n_1218),
.B(n_1219),
.Y(n_7212)
);

OAI21xp5_ASAP7_75t_L g7213 ( 
.A1(n_6919),
.A2(n_1224),
.B(n_1223),
.Y(n_7213)
);

AND2x2_ASAP7_75t_L g7214 ( 
.A(n_6993),
.B(n_1222),
.Y(n_7214)
);

NAND2xp5_ASAP7_75t_L g7215 ( 
.A(n_7047),
.B(n_1222),
.Y(n_7215)
);

INVx2_ASAP7_75t_L g7216 ( 
.A(n_6913),
.Y(n_7216)
);

NAND2xp5_ASAP7_75t_L g7217 ( 
.A(n_7069),
.B(n_1223),
.Y(n_7217)
);

OAI221xp5_ASAP7_75t_L g7218 ( 
.A1(n_7039),
.A2(n_1228),
.B1(n_1225),
.B2(n_1226),
.C(n_1229),
.Y(n_7218)
);

NAND2xp5_ASAP7_75t_L g7219 ( 
.A(n_7027),
.B(n_1226),
.Y(n_7219)
);

NAND2xp5_ASAP7_75t_L g7220 ( 
.A(n_7033),
.B(n_1228),
.Y(n_7220)
);

NOR2xp33_ASAP7_75t_L g7221 ( 
.A(n_7088),
.B(n_1229),
.Y(n_7221)
);

OAI21xp5_ASAP7_75t_L g7222 ( 
.A1(n_6941),
.A2(n_1232),
.B(n_1231),
.Y(n_7222)
);

OAI21xp33_ASAP7_75t_L g7223 ( 
.A1(n_7014),
.A2(n_1230),
.B(n_1231),
.Y(n_7223)
);

INVx1_ASAP7_75t_L g7224 ( 
.A(n_7009),
.Y(n_7224)
);

BUFx2_ASAP7_75t_L g7225 ( 
.A(n_6925),
.Y(n_7225)
);

INVxp33_ASAP7_75t_L g7226 ( 
.A(n_7050),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_6987),
.Y(n_7227)
);

AND2x2_ASAP7_75t_L g7228 ( 
.A(n_6994),
.B(n_1232),
.Y(n_7228)
);

INVx2_ASAP7_75t_L g7229 ( 
.A(n_7000),
.Y(n_7229)
);

NAND2xp5_ASAP7_75t_L g7230 ( 
.A(n_6907),
.B(n_1235),
.Y(n_7230)
);

AOI211xp5_ASAP7_75t_L g7231 ( 
.A1(n_6959),
.A2(n_1243),
.B(n_1254),
.C(n_1235),
.Y(n_7231)
);

INVx1_ASAP7_75t_L g7232 ( 
.A(n_7010),
.Y(n_7232)
);

NAND2xp5_ASAP7_75t_L g7233 ( 
.A(n_6902),
.B(n_6929),
.Y(n_7233)
);

AOI222xp33_ASAP7_75t_SL g7234 ( 
.A1(n_7020),
.A2(n_6923),
.B1(n_6965),
.B2(n_6983),
.C1(n_6986),
.C2(n_7007),
.Y(n_7234)
);

INVx2_ASAP7_75t_L g7235 ( 
.A(n_7018),
.Y(n_7235)
);

AOI322xp5_ASAP7_75t_L g7236 ( 
.A1(n_6926),
.A2(n_6938),
.A3(n_7015),
.B1(n_7019),
.B2(n_6999),
.C1(n_6917),
.C2(n_6966),
.Y(n_7236)
);

AOI222xp33_ASAP7_75t_L g7237 ( 
.A1(n_6947),
.A2(n_1238),
.B1(n_1240),
.B2(n_1236),
.C1(n_1237),
.C2(n_1239),
.Y(n_7237)
);

INVx1_ASAP7_75t_L g7238 ( 
.A(n_7017),
.Y(n_7238)
);

OAI222xp33_ASAP7_75t_L g7239 ( 
.A1(n_7177),
.A2(n_6968),
.B1(n_7037),
.B2(n_7075),
.C1(n_7053),
.C2(n_7036),
.Y(n_7239)
);

AOI21xp5_ASAP7_75t_L g7240 ( 
.A1(n_7108),
.A2(n_6916),
.B(n_7081),
.Y(n_7240)
);

AOI22xp33_ASAP7_75t_L g7241 ( 
.A1(n_7095),
.A2(n_6992),
.B1(n_6922),
.B2(n_7091),
.Y(n_7241)
);

O2A1O1Ixp33_ASAP7_75t_L g7242 ( 
.A1(n_7196),
.A2(n_7004),
.B(n_6939),
.C(n_6984),
.Y(n_7242)
);

AO21x1_ASAP7_75t_L g7243 ( 
.A1(n_7112),
.A2(n_6974),
.B(n_6944),
.Y(n_7243)
);

AND2x2_ASAP7_75t_L g7244 ( 
.A(n_7097),
.B(n_7107),
.Y(n_7244)
);

INVx1_ASAP7_75t_L g7245 ( 
.A(n_7225),
.Y(n_7245)
);

OAI22xp5_ASAP7_75t_L g7246 ( 
.A1(n_7159),
.A2(n_6946),
.B1(n_6940),
.B2(n_7046),
.Y(n_7246)
);

NAND2xp5_ASAP7_75t_L g7247 ( 
.A(n_7098),
.B(n_6922),
.Y(n_7247)
);

AOI22xp5_ASAP7_75t_L g7248 ( 
.A1(n_7150),
.A2(n_6910),
.B1(n_6995),
.B2(n_6996),
.Y(n_7248)
);

OAI22xp33_ASAP7_75t_L g7249 ( 
.A1(n_7117),
.A2(n_7174),
.B1(n_7093),
.B2(n_7216),
.Y(n_7249)
);

AOI221xp5_ASAP7_75t_L g7250 ( 
.A1(n_7206),
.A2(n_6973),
.B1(n_7013),
.B2(n_6978),
.C(n_6991),
.Y(n_7250)
);

OAI211xp5_ASAP7_75t_SL g7251 ( 
.A1(n_7126),
.A2(n_7012),
.B(n_6982),
.C(n_7016),
.Y(n_7251)
);

INVxp67_ASAP7_75t_L g7252 ( 
.A(n_7189),
.Y(n_7252)
);

NAND2xp5_ASAP7_75t_L g7253 ( 
.A(n_7140),
.B(n_6998),
.Y(n_7253)
);

INVx1_ASAP7_75t_L g7254 ( 
.A(n_7113),
.Y(n_7254)
);

OR2x2_ASAP7_75t_L g7255 ( 
.A(n_7121),
.B(n_1236),
.Y(n_7255)
);

NAND4xp25_ASAP7_75t_L g7256 ( 
.A(n_7236),
.B(n_1241),
.C(n_1238),
.D(n_1239),
.Y(n_7256)
);

INVx1_ASAP7_75t_L g7257 ( 
.A(n_7113),
.Y(n_7257)
);

INVx1_ASAP7_75t_L g7258 ( 
.A(n_7178),
.Y(n_7258)
);

NAND2xp5_ASAP7_75t_L g7259 ( 
.A(n_7186),
.B(n_1242),
.Y(n_7259)
);

AOI21xp5_ASAP7_75t_L g7260 ( 
.A1(n_7124),
.A2(n_1242),
.B(n_1243),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_7100),
.Y(n_7261)
);

INVx1_ASAP7_75t_L g7262 ( 
.A(n_7111),
.Y(n_7262)
);

INVx3_ASAP7_75t_L g7263 ( 
.A(n_7151),
.Y(n_7263)
);

BUFx2_ASAP7_75t_SL g7264 ( 
.A(n_7096),
.Y(n_7264)
);

AO21x1_ASAP7_75t_L g7265 ( 
.A1(n_7102),
.A2(n_1244),
.B(n_1245),
.Y(n_7265)
);

INVx2_ASAP7_75t_L g7266 ( 
.A(n_7121),
.Y(n_7266)
);

OAI211xp5_ASAP7_75t_SL g7267 ( 
.A1(n_7224),
.A2(n_1248),
.B(n_1245),
.C(n_1247),
.Y(n_7267)
);

INVx1_ASAP7_75t_L g7268 ( 
.A(n_7141),
.Y(n_7268)
);

INVx2_ASAP7_75t_L g7269 ( 
.A(n_7179),
.Y(n_7269)
);

OAI21xp33_ASAP7_75t_L g7270 ( 
.A1(n_7226),
.A2(n_1247),
.B(n_1248),
.Y(n_7270)
);

INVx2_ASAP7_75t_SL g7271 ( 
.A(n_7163),
.Y(n_7271)
);

INVx1_ASAP7_75t_L g7272 ( 
.A(n_7109),
.Y(n_7272)
);

INVx1_ASAP7_75t_L g7273 ( 
.A(n_7188),
.Y(n_7273)
);

INVx1_ASAP7_75t_L g7274 ( 
.A(n_7106),
.Y(n_7274)
);

INVxp33_ASAP7_75t_L g7275 ( 
.A(n_7128),
.Y(n_7275)
);

AND2x2_ASAP7_75t_L g7276 ( 
.A(n_7130),
.B(n_1250),
.Y(n_7276)
);

INVx1_ASAP7_75t_SL g7277 ( 
.A(n_7132),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_7101),
.Y(n_7278)
);

INVx1_ASAP7_75t_L g7279 ( 
.A(n_7172),
.Y(n_7279)
);

AOI222xp33_ASAP7_75t_L g7280 ( 
.A1(n_7161),
.A2(n_1254),
.B1(n_1256),
.B2(n_1251),
.C1(n_1253),
.C2(n_1255),
.Y(n_7280)
);

INVx1_ASAP7_75t_L g7281 ( 
.A(n_7148),
.Y(n_7281)
);

INVx2_ASAP7_75t_L g7282 ( 
.A(n_7171),
.Y(n_7282)
);

AOI21xp33_ASAP7_75t_L g7283 ( 
.A1(n_7208),
.A2(n_1253),
.B(n_1255),
.Y(n_7283)
);

INVx1_ASAP7_75t_L g7284 ( 
.A(n_7228),
.Y(n_7284)
);

AOI21xp33_ASAP7_75t_L g7285 ( 
.A1(n_7166),
.A2(n_1256),
.B(n_1257),
.Y(n_7285)
);

INVx2_ASAP7_75t_L g7286 ( 
.A(n_7202),
.Y(n_7286)
);

AOI32xp33_ASAP7_75t_L g7287 ( 
.A1(n_7131),
.A2(n_1262),
.A3(n_1259),
.B1(n_1260),
.B2(n_1263),
.Y(n_7287)
);

AND2x4_ASAP7_75t_L g7288 ( 
.A(n_7125),
.B(n_1259),
.Y(n_7288)
);

OR2x6_ASAP7_75t_L g7289 ( 
.A(n_7203),
.B(n_1262),
.Y(n_7289)
);

OAI31xp33_ASAP7_75t_L g7290 ( 
.A1(n_7094),
.A2(n_7116),
.A3(n_7120),
.B(n_7183),
.Y(n_7290)
);

NOR2xp33_ASAP7_75t_L g7291 ( 
.A(n_7114),
.B(n_1263),
.Y(n_7291)
);

OAI22xp5_ASAP7_75t_L g7292 ( 
.A1(n_7185),
.A2(n_7210),
.B1(n_7217),
.B2(n_7215),
.Y(n_7292)
);

AND2x2_ASAP7_75t_L g7293 ( 
.A(n_7167),
.B(n_1264),
.Y(n_7293)
);

O2A1O1Ixp33_ASAP7_75t_L g7294 ( 
.A1(n_7190),
.A2(n_1267),
.B(n_1265),
.C(n_1266),
.Y(n_7294)
);

INVx1_ASAP7_75t_L g7295 ( 
.A(n_7162),
.Y(n_7295)
);

OAI221xp5_ASAP7_75t_L g7296 ( 
.A1(n_7157),
.A2(n_1269),
.B1(n_1266),
.B2(n_1268),
.C(n_1270),
.Y(n_7296)
);

INVx2_ASAP7_75t_SL g7297 ( 
.A(n_7165),
.Y(n_7297)
);

OAI22xp5_ASAP7_75t_L g7298 ( 
.A1(n_7233),
.A2(n_1271),
.B1(n_1269),
.B2(n_1270),
.Y(n_7298)
);

AND2x2_ASAP7_75t_L g7299 ( 
.A(n_7184),
.B(n_1271),
.Y(n_7299)
);

OAI221xp5_ASAP7_75t_L g7300 ( 
.A1(n_7122),
.A2(n_1274),
.B1(n_1272),
.B2(n_1273),
.C(n_1275),
.Y(n_7300)
);

AOI21xp33_ASAP7_75t_SL g7301 ( 
.A1(n_7110),
.A2(n_1275),
.B(n_1274),
.Y(n_7301)
);

OR2x2_ASAP7_75t_L g7302 ( 
.A(n_7123),
.B(n_1273),
.Y(n_7302)
);

INVxp67_ASAP7_75t_SL g7303 ( 
.A(n_7158),
.Y(n_7303)
);

OAI22xp5_ASAP7_75t_L g7304 ( 
.A1(n_7194),
.A2(n_1278),
.B1(n_1276),
.B2(n_1277),
.Y(n_7304)
);

OAI21xp5_ASAP7_75t_SL g7305 ( 
.A1(n_7211),
.A2(n_1276),
.B(n_1277),
.Y(n_7305)
);

AOI222xp33_ASAP7_75t_L g7306 ( 
.A1(n_7127),
.A2(n_7138),
.B1(n_7129),
.B2(n_7139),
.C1(n_7135),
.C2(n_7134),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_7214),
.Y(n_7307)
);

AOI321xp33_ASAP7_75t_L g7308 ( 
.A1(n_7192),
.A2(n_1280),
.A3(n_1282),
.B1(n_1278),
.B2(n_1279),
.C(n_1281),
.Y(n_7308)
);

OR2x2_ASAP7_75t_L g7309 ( 
.A(n_7133),
.B(n_1279),
.Y(n_7309)
);

INVx1_ASAP7_75t_L g7310 ( 
.A(n_7204),
.Y(n_7310)
);

AND2x4_ASAP7_75t_L g7311 ( 
.A(n_7170),
.B(n_1280),
.Y(n_7311)
);

INVx1_ASAP7_75t_L g7312 ( 
.A(n_7136),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_7099),
.Y(n_7313)
);

AOI222xp33_ASAP7_75t_L g7314 ( 
.A1(n_7142),
.A2(n_1285),
.B1(n_1287),
.B2(n_1283),
.C1(n_1284),
.C2(n_1286),
.Y(n_7314)
);

OR2x2_ASAP7_75t_L g7315 ( 
.A(n_7193),
.B(n_1283),
.Y(n_7315)
);

INVx1_ASAP7_75t_L g7316 ( 
.A(n_7143),
.Y(n_7316)
);

BUFx2_ASAP7_75t_L g7317 ( 
.A(n_7229),
.Y(n_7317)
);

OAI222xp33_ASAP7_75t_L g7318 ( 
.A1(n_7144),
.A2(n_1286),
.B1(n_1289),
.B2(n_1284),
.C1(n_1285),
.C2(n_1288),
.Y(n_7318)
);

INVx1_ASAP7_75t_L g7319 ( 
.A(n_7146),
.Y(n_7319)
);

NAND2xp5_ASAP7_75t_L g7320 ( 
.A(n_7145),
.B(n_1288),
.Y(n_7320)
);

OAI32xp33_ASAP7_75t_L g7321 ( 
.A1(n_7147),
.A2(n_1292),
.A3(n_1294),
.B1(n_1291),
.B2(n_1293),
.Y(n_7321)
);

INVx1_ASAP7_75t_L g7322 ( 
.A(n_7149),
.Y(n_7322)
);

AOI221xp5_ASAP7_75t_L g7323 ( 
.A1(n_7154),
.A2(n_1293),
.B1(n_1290),
.B2(n_1291),
.C(n_1295),
.Y(n_7323)
);

NAND3xp33_ASAP7_75t_SL g7324 ( 
.A(n_7118),
.B(n_1297),
.C(n_1296),
.Y(n_7324)
);

AOI22xp33_ASAP7_75t_L g7325 ( 
.A1(n_7176),
.A2(n_1297),
.B1(n_1290),
.B2(n_1296),
.Y(n_7325)
);

OAI21xp33_ASAP7_75t_SL g7326 ( 
.A1(n_7155),
.A2(n_1298),
.B(n_1300),
.Y(n_7326)
);

NOR2xp67_ASAP7_75t_L g7327 ( 
.A(n_7168),
.B(n_1298),
.Y(n_7327)
);

A2O1A1Ixp33_ASAP7_75t_L g7328 ( 
.A1(n_7207),
.A2(n_1310),
.B(n_1319),
.C(n_1301),
.Y(n_7328)
);

AOI221xp5_ASAP7_75t_L g7329 ( 
.A1(n_7156),
.A2(n_1305),
.B1(n_1302),
.B2(n_1304),
.C(n_1306),
.Y(n_7329)
);

AND2x2_ASAP7_75t_L g7330 ( 
.A(n_7181),
.B(n_1305),
.Y(n_7330)
);

AOI22xp33_ASAP7_75t_L g7331 ( 
.A1(n_7103),
.A2(n_1308),
.B1(n_1306),
.B2(n_1307),
.Y(n_7331)
);

AND2x2_ASAP7_75t_L g7332 ( 
.A(n_7195),
.B(n_1307),
.Y(n_7332)
);

OAI221xp5_ASAP7_75t_L g7333 ( 
.A1(n_7222),
.A2(n_1311),
.B1(n_1309),
.B2(n_1310),
.C(n_1312),
.Y(n_7333)
);

NAND2xp5_ASAP7_75t_L g7334 ( 
.A(n_7187),
.B(n_1309),
.Y(n_7334)
);

NAND2xp5_ASAP7_75t_L g7335 ( 
.A(n_7115),
.B(n_1313),
.Y(n_7335)
);

OAI221xp5_ASAP7_75t_L g7336 ( 
.A1(n_7105),
.A2(n_1315),
.B1(n_1313),
.B2(n_1314),
.C(n_1317),
.Y(n_7336)
);

OAI22xp5_ASAP7_75t_L g7337 ( 
.A1(n_7218),
.A2(n_1319),
.B1(n_1317),
.B2(n_1318),
.Y(n_7337)
);

INVx1_ASAP7_75t_L g7338 ( 
.A(n_7160),
.Y(n_7338)
);

INVx1_ASAP7_75t_L g7339 ( 
.A(n_7180),
.Y(n_7339)
);

NOR2xp67_ASAP7_75t_SL g7340 ( 
.A(n_7119),
.B(n_1321),
.Y(n_7340)
);

NAND2xp5_ASAP7_75t_L g7341 ( 
.A(n_7237),
.B(n_1318),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_L g7342 ( 
.A(n_7104),
.B(n_1321),
.Y(n_7342)
);

AOI22xp5_ASAP7_75t_L g7343 ( 
.A1(n_7234),
.A2(n_1324),
.B1(n_1322),
.B2(n_1323),
.Y(n_7343)
);

INVx1_ASAP7_75t_L g7344 ( 
.A(n_7227),
.Y(n_7344)
);

NAND2x1p5_ASAP7_75t_L g7345 ( 
.A(n_7232),
.B(n_1322),
.Y(n_7345)
);

AOI21xp5_ASAP7_75t_L g7346 ( 
.A1(n_7197),
.A2(n_1323),
.B(n_1324),
.Y(n_7346)
);

OAI21xp33_ASAP7_75t_L g7347 ( 
.A1(n_7238),
.A2(n_7198),
.B(n_7201),
.Y(n_7347)
);

NAND2xp5_ASAP7_75t_L g7348 ( 
.A(n_7221),
.B(n_1325),
.Y(n_7348)
);

AOI221xp5_ASAP7_75t_L g7349 ( 
.A1(n_7212),
.A2(n_1327),
.B1(n_1325),
.B2(n_1326),
.C(n_1328),
.Y(n_7349)
);

AOI311xp33_ASAP7_75t_L g7350 ( 
.A1(n_7209),
.A2(n_1328),
.A3(n_1326),
.B(n_1327),
.C(n_1329),
.Y(n_7350)
);

INVx1_ASAP7_75t_L g7351 ( 
.A(n_7219),
.Y(n_7351)
);

O2A1O1Ixp33_ASAP7_75t_L g7352 ( 
.A1(n_7213),
.A2(n_1331),
.B(n_1329),
.C(n_1330),
.Y(n_7352)
);

INVx1_ASAP7_75t_L g7353 ( 
.A(n_7220),
.Y(n_7353)
);

AOI21xp33_ASAP7_75t_L g7354 ( 
.A1(n_7191),
.A2(n_1330),
.B(n_1331),
.Y(n_7354)
);

INVx2_ASAP7_75t_L g7355 ( 
.A(n_7235),
.Y(n_7355)
);

INVx1_ASAP7_75t_L g7356 ( 
.A(n_7199),
.Y(n_7356)
);

OAI332xp33_ASAP7_75t_L g7357 ( 
.A1(n_7153),
.A2(n_1338),
.A3(n_1337),
.B1(n_1334),
.B2(n_1339),
.B3(n_1332),
.C1(n_1333),
.C2(n_1336),
.Y(n_7357)
);

NAND2xp5_ASAP7_75t_L g7358 ( 
.A(n_7231),
.B(n_1332),
.Y(n_7358)
);

AOI22xp5_ASAP7_75t_L g7359 ( 
.A1(n_7152),
.A2(n_1337),
.B1(n_1334),
.B2(n_1336),
.Y(n_7359)
);

A2O1A1Ixp33_ASAP7_75t_SL g7360 ( 
.A1(n_7205),
.A2(n_1340),
.B(n_1338),
.C(n_1339),
.Y(n_7360)
);

NAND2xp5_ASAP7_75t_L g7361 ( 
.A(n_7223),
.B(n_1341),
.Y(n_7361)
);

OAI22xp33_ASAP7_75t_L g7362 ( 
.A1(n_7173),
.A2(n_1345),
.B1(n_1342),
.B2(n_1343),
.Y(n_7362)
);

INVx1_ASAP7_75t_L g7363 ( 
.A(n_7175),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_7182),
.Y(n_7364)
);

INVx1_ASAP7_75t_L g7365 ( 
.A(n_7230),
.Y(n_7365)
);

INVxp67_ASAP7_75t_L g7366 ( 
.A(n_7164),
.Y(n_7366)
);

AOI21xp33_ASAP7_75t_L g7367 ( 
.A1(n_7169),
.A2(n_1342),
.B(n_1343),
.Y(n_7367)
);

INVx1_ASAP7_75t_L g7368 ( 
.A(n_7200),
.Y(n_7368)
);

INVx2_ASAP7_75t_L g7369 ( 
.A(n_7137),
.Y(n_7369)
);

AOI22xp5_ASAP7_75t_L g7370 ( 
.A1(n_7095),
.A2(n_1348),
.B1(n_1345),
.B2(n_1347),
.Y(n_7370)
);

AOI22xp5_ASAP7_75t_L g7371 ( 
.A1(n_7095),
.A2(n_1350),
.B1(n_1348),
.B2(n_1349),
.Y(n_7371)
);

NAND2xp5_ASAP7_75t_L g7372 ( 
.A(n_7095),
.B(n_1350),
.Y(n_7372)
);

OA22x2_ASAP7_75t_L g7373 ( 
.A1(n_7095),
.A2(n_1353),
.B1(n_1351),
.B2(n_1352),
.Y(n_7373)
);

BUFx2_ASAP7_75t_L g7374 ( 
.A(n_7113),
.Y(n_7374)
);

AND2x2_ASAP7_75t_L g7375 ( 
.A(n_7095),
.B(n_1352),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_7196),
.Y(n_7376)
);

NAND2xp5_ASAP7_75t_L g7377 ( 
.A(n_7095),
.B(n_1353),
.Y(n_7377)
);

AND2x4_ASAP7_75t_L g7378 ( 
.A(n_7095),
.B(n_1354),
.Y(n_7378)
);

INVx1_ASAP7_75t_L g7379 ( 
.A(n_7196),
.Y(n_7379)
);

AOI22xp5_ASAP7_75t_L g7380 ( 
.A1(n_7095),
.A2(n_1356),
.B1(n_1354),
.B2(n_1355),
.Y(n_7380)
);

O2A1O1Ixp33_ASAP7_75t_L g7381 ( 
.A1(n_7177),
.A2(n_1357),
.B(n_1355),
.C(n_1356),
.Y(n_7381)
);

OAI221xp5_ASAP7_75t_L g7382 ( 
.A1(n_7177),
.A2(n_1359),
.B1(n_1357),
.B2(n_1358),
.C(n_1360),
.Y(n_7382)
);

AOI21xp5_ASAP7_75t_L g7383 ( 
.A1(n_7177),
.A2(n_1359),
.B(n_1360),
.Y(n_7383)
);

OAI22xp5_ASAP7_75t_L g7384 ( 
.A1(n_7177),
.A2(n_1363),
.B1(n_1361),
.B2(n_1362),
.Y(n_7384)
);

AND2x4_ASAP7_75t_L g7385 ( 
.A(n_7095),
.B(n_1361),
.Y(n_7385)
);

INVx2_ASAP7_75t_L g7386 ( 
.A(n_7113),
.Y(n_7386)
);

A2O1A1Ixp33_ASAP7_75t_L g7387 ( 
.A1(n_7177),
.A2(n_1371),
.B(n_1380),
.C(n_1363),
.Y(n_7387)
);

NAND2xp5_ASAP7_75t_L g7388 ( 
.A(n_7095),
.B(n_1364),
.Y(n_7388)
);

NAND2xp5_ASAP7_75t_L g7389 ( 
.A(n_7095),
.B(n_1365),
.Y(n_7389)
);

O2A1O1Ixp33_ASAP7_75t_L g7390 ( 
.A1(n_7177),
.A2(n_1367),
.B(n_1365),
.C(n_1366),
.Y(n_7390)
);

OAI21xp33_ASAP7_75t_SL g7391 ( 
.A1(n_7177),
.A2(n_1366),
.B(n_1368),
.Y(n_7391)
);

INVx2_ASAP7_75t_L g7392 ( 
.A(n_7113),
.Y(n_7392)
);

OAI222xp33_ASAP7_75t_L g7393 ( 
.A1(n_7177),
.A2(n_1370),
.B1(n_1373),
.B2(n_1368),
.C1(n_1369),
.C2(n_1372),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_7196),
.Y(n_7394)
);

NAND3xp33_ASAP7_75t_SL g7395 ( 
.A(n_7095),
.B(n_1373),
.C(n_1372),
.Y(n_7395)
);

INVx1_ASAP7_75t_L g7396 ( 
.A(n_7196),
.Y(n_7396)
);

NAND2xp5_ASAP7_75t_L g7397 ( 
.A(n_7095),
.B(n_1369),
.Y(n_7397)
);

NOR2xp33_ASAP7_75t_L g7398 ( 
.A(n_7095),
.B(n_1374),
.Y(n_7398)
);

NAND2xp5_ASAP7_75t_L g7399 ( 
.A(n_7095),
.B(n_1375),
.Y(n_7399)
);

AOI22xp5_ASAP7_75t_L g7400 ( 
.A1(n_7095),
.A2(n_1377),
.B1(n_1375),
.B2(n_1376),
.Y(n_7400)
);

OAI21xp33_ASAP7_75t_SL g7401 ( 
.A1(n_7177),
.A2(n_1376),
.B(n_1377),
.Y(n_7401)
);

INVx1_ASAP7_75t_L g7402 ( 
.A(n_7196),
.Y(n_7402)
);

NAND2xp5_ASAP7_75t_SL g7403 ( 
.A(n_7374),
.B(n_1378),
.Y(n_7403)
);

INVx1_ASAP7_75t_L g7404 ( 
.A(n_7255),
.Y(n_7404)
);

NAND3xp33_ASAP7_75t_L g7405 ( 
.A(n_7245),
.B(n_1378),
.C(n_1380),
.Y(n_7405)
);

NAND2xp5_ASAP7_75t_L g7406 ( 
.A(n_7252),
.B(n_1381),
.Y(n_7406)
);

OR2x2_ASAP7_75t_L g7407 ( 
.A(n_7395),
.B(n_1381),
.Y(n_7407)
);

NOR2xp33_ASAP7_75t_L g7408 ( 
.A(n_7239),
.B(n_7266),
.Y(n_7408)
);

NAND3xp33_ASAP7_75t_L g7409 ( 
.A(n_7343),
.B(n_1382),
.C(n_1383),
.Y(n_7409)
);

NOR2xp67_ASAP7_75t_L g7410 ( 
.A(n_7326),
.B(n_1382),
.Y(n_7410)
);

OR2x2_ASAP7_75t_L g7411 ( 
.A(n_7247),
.B(n_1384),
.Y(n_7411)
);

NAND2xp5_ASAP7_75t_L g7412 ( 
.A(n_7378),
.B(n_7254),
.Y(n_7412)
);

NAND2xp5_ASAP7_75t_SL g7413 ( 
.A(n_7327),
.B(n_1385),
.Y(n_7413)
);

NAND2xp5_ASAP7_75t_L g7414 ( 
.A(n_7378),
.B(n_1385),
.Y(n_7414)
);

AOI211xp5_ASAP7_75t_L g7415 ( 
.A1(n_7249),
.A2(n_1388),
.B(n_1386),
.C(n_1387),
.Y(n_7415)
);

NAND2xp5_ASAP7_75t_L g7416 ( 
.A(n_7257),
.B(n_1386),
.Y(n_7416)
);

OAI21xp33_ASAP7_75t_L g7417 ( 
.A1(n_7241),
.A2(n_1398),
.B(n_1389),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_7376),
.Y(n_7418)
);

NAND2xp5_ASAP7_75t_L g7419 ( 
.A(n_7386),
.B(n_1389),
.Y(n_7419)
);

AO21x1_ASAP7_75t_L g7420 ( 
.A1(n_7379),
.A2(n_1390),
.B(n_1392),
.Y(n_7420)
);

INVx1_ASAP7_75t_L g7421 ( 
.A(n_7394),
.Y(n_7421)
);

INVx1_ASAP7_75t_L g7422 ( 
.A(n_7396),
.Y(n_7422)
);

NAND2xp5_ASAP7_75t_L g7423 ( 
.A(n_7392),
.B(n_1390),
.Y(n_7423)
);

OR2x2_ASAP7_75t_L g7424 ( 
.A(n_7256),
.B(n_1392),
.Y(n_7424)
);

NOR2xp33_ASAP7_75t_L g7425 ( 
.A(n_7275),
.B(n_1393),
.Y(n_7425)
);

OAI21xp33_ASAP7_75t_SL g7426 ( 
.A1(n_7402),
.A2(n_1393),
.B(n_1394),
.Y(n_7426)
);

INVx2_ASAP7_75t_L g7427 ( 
.A(n_7345),
.Y(n_7427)
);

NAND3xp33_ASAP7_75t_SL g7428 ( 
.A(n_7290),
.B(n_1394),
.C(n_1395),
.Y(n_7428)
);

INVx2_ASAP7_75t_SL g7429 ( 
.A(n_7244),
.Y(n_7429)
);

NOR3x1_ASAP7_75t_L g7430 ( 
.A(n_7324),
.B(n_1395),
.C(n_1396),
.Y(n_7430)
);

INVx1_ASAP7_75t_L g7431 ( 
.A(n_7375),
.Y(n_7431)
);

INVx1_ASAP7_75t_L g7432 ( 
.A(n_7264),
.Y(n_7432)
);

AND2x2_ASAP7_75t_L g7433 ( 
.A(n_7269),
.B(n_1396),
.Y(n_7433)
);

OAI21xp5_ASAP7_75t_L g7434 ( 
.A1(n_7240),
.A2(n_1397),
.B(n_1398),
.Y(n_7434)
);

OAI21xp5_ASAP7_75t_L g7435 ( 
.A1(n_7391),
.A2(n_1397),
.B(n_1399),
.Y(n_7435)
);

OAI21xp33_ASAP7_75t_L g7436 ( 
.A1(n_7248),
.A2(n_1408),
.B(n_1399),
.Y(n_7436)
);

NOR2xp33_ASAP7_75t_SL g7437 ( 
.A(n_7393),
.B(n_1400),
.Y(n_7437)
);

NAND2xp5_ASAP7_75t_L g7438 ( 
.A(n_7385),
.B(n_1402),
.Y(n_7438)
);

AOI21xp5_ASAP7_75t_L g7439 ( 
.A1(n_7242),
.A2(n_1402),
.B(n_1403),
.Y(n_7439)
);

INVx1_ASAP7_75t_L g7440 ( 
.A(n_7373),
.Y(n_7440)
);

OAI21xp33_ASAP7_75t_SL g7441 ( 
.A1(n_7303),
.A2(n_1404),
.B(n_1405),
.Y(n_7441)
);

AOI22xp5_ASAP7_75t_L g7442 ( 
.A1(n_7243),
.A2(n_1406),
.B1(n_1404),
.B2(n_1405),
.Y(n_7442)
);

AND2x4_ASAP7_75t_L g7443 ( 
.A(n_7271),
.B(n_1406),
.Y(n_7443)
);

INVx1_ASAP7_75t_L g7444 ( 
.A(n_7253),
.Y(n_7444)
);

INVx1_ASAP7_75t_SL g7445 ( 
.A(n_7317),
.Y(n_7445)
);

AND2x2_ASAP7_75t_L g7446 ( 
.A(n_7263),
.B(n_1407),
.Y(n_7446)
);

NOR2xp33_ASAP7_75t_L g7447 ( 
.A(n_7401),
.B(n_1407),
.Y(n_7447)
);

OAI21xp5_ASAP7_75t_SL g7448 ( 
.A1(n_7250),
.A2(n_1408),
.B(n_1409),
.Y(n_7448)
);

OAI21xp5_ASAP7_75t_L g7449 ( 
.A1(n_7328),
.A2(n_1410),
.B(n_1411),
.Y(n_7449)
);

INVxp67_ASAP7_75t_SL g7450 ( 
.A(n_7265),
.Y(n_7450)
);

AOI22xp5_ASAP7_75t_L g7451 ( 
.A1(n_7246),
.A2(n_1413),
.B1(n_1410),
.B2(n_1412),
.Y(n_7451)
);

AOI211xp5_ASAP7_75t_L g7452 ( 
.A1(n_7285),
.A2(n_1415),
.B(n_1412),
.C(n_1414),
.Y(n_7452)
);

AOI21xp33_ASAP7_75t_SL g7453 ( 
.A1(n_7294),
.A2(n_1417),
.B(n_1416),
.Y(n_7453)
);

AOI221xp5_ASAP7_75t_L g7454 ( 
.A1(n_7251),
.A2(n_7356),
.B1(n_7381),
.B2(n_7390),
.C(n_7347),
.Y(n_7454)
);

NAND2xp5_ASAP7_75t_L g7455 ( 
.A(n_7258),
.B(n_7291),
.Y(n_7455)
);

INVx1_ASAP7_75t_L g7456 ( 
.A(n_7293),
.Y(n_7456)
);

NOR3x1_ASAP7_75t_L g7457 ( 
.A(n_7360),
.B(n_7305),
.C(n_7300),
.Y(n_7457)
);

NAND2xp5_ASAP7_75t_L g7458 ( 
.A(n_7311),
.B(n_1414),
.Y(n_7458)
);

BUFx2_ASAP7_75t_L g7459 ( 
.A(n_7289),
.Y(n_7459)
);

NOR2xp33_ASAP7_75t_L g7460 ( 
.A(n_7301),
.B(n_1416),
.Y(n_7460)
);

AOI211xp5_ASAP7_75t_SL g7461 ( 
.A1(n_7292),
.A2(n_1420),
.B(n_1418),
.C(n_1419),
.Y(n_7461)
);

NOR3x1_ASAP7_75t_L g7462 ( 
.A(n_7297),
.B(n_1420),
.C(n_1421),
.Y(n_7462)
);

NAND2xp5_ASAP7_75t_L g7463 ( 
.A(n_7311),
.B(n_7398),
.Y(n_7463)
);

NAND3xp33_ASAP7_75t_L g7464 ( 
.A(n_7306),
.B(n_1421),
.C(n_1422),
.Y(n_7464)
);

NAND2xp5_ASAP7_75t_L g7465 ( 
.A(n_7330),
.B(n_1422),
.Y(n_7465)
);

INVx1_ASAP7_75t_L g7466 ( 
.A(n_7372),
.Y(n_7466)
);

AOI211xp5_ASAP7_75t_L g7467 ( 
.A1(n_7274),
.A2(n_1425),
.B(n_1423),
.C(n_1424),
.Y(n_7467)
);

NAND2xp33_ASAP7_75t_SL g7468 ( 
.A(n_7340),
.B(n_1423),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_7377),
.Y(n_7469)
);

OAI211xp5_ASAP7_75t_L g7470 ( 
.A1(n_7280),
.A2(n_1428),
.B(n_1426),
.C(n_1427),
.Y(n_7470)
);

INVx1_ASAP7_75t_L g7471 ( 
.A(n_7388),
.Y(n_7471)
);

AND2x2_ASAP7_75t_L g7472 ( 
.A(n_7282),
.B(n_1426),
.Y(n_7472)
);

NAND2xp5_ASAP7_75t_L g7473 ( 
.A(n_7276),
.B(n_1428),
.Y(n_7473)
);

INVx1_ASAP7_75t_L g7474 ( 
.A(n_7389),
.Y(n_7474)
);

NOR2xp67_ASAP7_75t_SL g7475 ( 
.A(n_7261),
.B(n_1429),
.Y(n_7475)
);

NAND3xp33_ASAP7_75t_SL g7476 ( 
.A(n_7277),
.B(n_1430),
.C(n_1431),
.Y(n_7476)
);

CKINVDCx20_ASAP7_75t_R g7477 ( 
.A(n_7268),
.Y(n_7477)
);

OAI22xp33_ASAP7_75t_SL g7478 ( 
.A1(n_7368),
.A2(n_1432),
.B1(n_1430),
.B2(n_1431),
.Y(n_7478)
);

NOR2xp33_ASAP7_75t_L g7479 ( 
.A(n_7296),
.B(n_1432),
.Y(n_7479)
);

INVx1_ASAP7_75t_L g7480 ( 
.A(n_7397),
.Y(n_7480)
);

AOI21xp33_ASAP7_75t_L g7481 ( 
.A1(n_7278),
.A2(n_7273),
.B(n_7281),
.Y(n_7481)
);

INVxp67_ASAP7_75t_L g7482 ( 
.A(n_7289),
.Y(n_7482)
);

NAND2xp5_ASAP7_75t_L g7483 ( 
.A(n_7383),
.B(n_1433),
.Y(n_7483)
);

NOR2xp33_ASAP7_75t_L g7484 ( 
.A(n_7270),
.B(n_1433),
.Y(n_7484)
);

AOI22xp5_ASAP7_75t_L g7485 ( 
.A1(n_7369),
.A2(n_1436),
.B1(n_1434),
.B2(n_1435),
.Y(n_7485)
);

NAND2xp5_ASAP7_75t_SL g7486 ( 
.A(n_7350),
.B(n_1436),
.Y(n_7486)
);

NAND2xp5_ASAP7_75t_SL g7487 ( 
.A(n_7308),
.B(n_1438),
.Y(n_7487)
);

NOR3x1_ASAP7_75t_L g7488 ( 
.A(n_7341),
.B(n_1438),
.C(n_1439),
.Y(n_7488)
);

NAND2xp5_ASAP7_75t_L g7489 ( 
.A(n_7299),
.B(n_1439),
.Y(n_7489)
);

AND2x2_ASAP7_75t_L g7490 ( 
.A(n_7279),
.B(n_7284),
.Y(n_7490)
);

NAND2xp5_ASAP7_75t_L g7491 ( 
.A(n_7332),
.B(n_1440),
.Y(n_7491)
);

INVx1_ASAP7_75t_L g7492 ( 
.A(n_7399),
.Y(n_7492)
);

INVx2_ASAP7_75t_L g7493 ( 
.A(n_7288),
.Y(n_7493)
);

NOR3xp33_ASAP7_75t_SL g7494 ( 
.A(n_7272),
.B(n_1440),
.C(n_1441),
.Y(n_7494)
);

NOR2xp33_ASAP7_75t_L g7495 ( 
.A(n_7382),
.B(n_1442),
.Y(n_7495)
);

NOR2xp67_ASAP7_75t_L g7496 ( 
.A(n_7286),
.B(n_1442),
.Y(n_7496)
);

INVx1_ASAP7_75t_L g7497 ( 
.A(n_7288),
.Y(n_7497)
);

OR2x2_ASAP7_75t_L g7498 ( 
.A(n_7259),
.B(n_1444),
.Y(n_7498)
);

NAND2xp5_ASAP7_75t_SL g7499 ( 
.A(n_7410),
.B(n_7287),
.Y(n_7499)
);

NAND2xp5_ASAP7_75t_L g7500 ( 
.A(n_7497),
.B(n_7447),
.Y(n_7500)
);

AOI221xp5_ASAP7_75t_L g7501 ( 
.A1(n_7408),
.A2(n_7454),
.B1(n_7450),
.B2(n_7428),
.C(n_7453),
.Y(n_7501)
);

OAI32xp33_ASAP7_75t_L g7502 ( 
.A1(n_7445),
.A2(n_7322),
.A3(n_7339),
.B1(n_7319),
.B2(n_7316),
.Y(n_7502)
);

AOI31xp33_ASAP7_75t_L g7503 ( 
.A1(n_7435),
.A2(n_7262),
.A3(n_7307),
.B(n_7295),
.Y(n_7503)
);

NOR2xp33_ASAP7_75t_L g7504 ( 
.A(n_7441),
.B(n_7482),
.Y(n_7504)
);

OAI32xp33_ASAP7_75t_L g7505 ( 
.A1(n_7440),
.A2(n_7344),
.A3(n_7355),
.B1(n_7353),
.B2(n_7351),
.Y(n_7505)
);

OAI21xp5_ASAP7_75t_SL g7506 ( 
.A1(n_7448),
.A2(n_7366),
.B(n_7338),
.Y(n_7506)
);

NAND4xp25_ASAP7_75t_L g7507 ( 
.A(n_7457),
.B(n_7313),
.C(n_7364),
.D(n_7363),
.Y(n_7507)
);

O2A1O1Ixp33_ASAP7_75t_L g7508 ( 
.A1(n_7487),
.A2(n_7387),
.B(n_7384),
.C(n_7318),
.Y(n_7508)
);

NAND2xp5_ASAP7_75t_L g7509 ( 
.A(n_7443),
.B(n_7260),
.Y(n_7509)
);

AOI222xp33_ASAP7_75t_L g7510 ( 
.A1(n_7417),
.A2(n_7365),
.B1(n_7310),
.B2(n_7312),
.C1(n_7329),
.C2(n_7323),
.Y(n_7510)
);

O2A1O1Ixp33_ASAP7_75t_L g7511 ( 
.A1(n_7486),
.A2(n_7267),
.B(n_7335),
.C(n_7321),
.Y(n_7511)
);

OAI21xp33_ASAP7_75t_SL g7512 ( 
.A1(n_7432),
.A2(n_7334),
.B(n_7320),
.Y(n_7512)
);

AOI221xp5_ASAP7_75t_L g7513 ( 
.A1(n_7464),
.A2(n_7367),
.B1(n_7362),
.B2(n_7352),
.C(n_7337),
.Y(n_7513)
);

NAND3xp33_ASAP7_75t_L g7514 ( 
.A(n_7415),
.B(n_7349),
.C(n_7346),
.Y(n_7514)
);

AOI221x1_ASAP7_75t_L g7515 ( 
.A1(n_7478),
.A2(n_7283),
.B1(n_7354),
.B2(n_7298),
.C(n_7358),
.Y(n_7515)
);

AOI221xp5_ASAP7_75t_L g7516 ( 
.A1(n_7439),
.A2(n_7357),
.B1(n_7304),
.B2(n_7333),
.C(n_7336),
.Y(n_7516)
);

AOI211xp5_ASAP7_75t_L g7517 ( 
.A1(n_7481),
.A2(n_7342),
.B(n_7348),
.C(n_7361),
.Y(n_7517)
);

O2A1O1Ixp33_ASAP7_75t_L g7518 ( 
.A1(n_7476),
.A2(n_7314),
.B(n_7315),
.C(n_7309),
.Y(n_7518)
);

AOI21xp33_ASAP7_75t_L g7519 ( 
.A1(n_7411),
.A2(n_7302),
.B(n_7359),
.Y(n_7519)
);

AOI22xp5_ASAP7_75t_L g7520 ( 
.A1(n_7477),
.A2(n_7400),
.B1(n_7371),
.B2(n_7380),
.Y(n_7520)
);

A2O1A1Ixp33_ASAP7_75t_L g7521 ( 
.A1(n_7442),
.A2(n_7370),
.B(n_7331),
.C(n_7325),
.Y(n_7521)
);

OAI211xp5_ASAP7_75t_L g7522 ( 
.A1(n_7426),
.A2(n_1453),
.B(n_1461),
.C(n_1444),
.Y(n_7522)
);

AND4x1_ASAP7_75t_L g7523 ( 
.A(n_7437),
.B(n_1447),
.C(n_1445),
.D(n_1446),
.Y(n_7523)
);

OAI221xp5_ASAP7_75t_L g7524 ( 
.A1(n_7434),
.A2(n_1449),
.B1(n_1446),
.B2(n_1447),
.C(n_1450),
.Y(n_7524)
);

AOI211xp5_ASAP7_75t_SL g7525 ( 
.A1(n_7470),
.A2(n_1451),
.B(n_1449),
.C(n_1450),
.Y(n_7525)
);

NOR3xp33_ASAP7_75t_L g7526 ( 
.A(n_7455),
.B(n_1452),
.C(n_1454),
.Y(n_7526)
);

AOI21xp5_ASAP7_75t_L g7527 ( 
.A1(n_7413),
.A2(n_1452),
.B(n_1454),
.Y(n_7527)
);

NOR2xp33_ASAP7_75t_L g7528 ( 
.A(n_7493),
.B(n_7459),
.Y(n_7528)
);

OAI211xp5_ASAP7_75t_L g7529 ( 
.A1(n_7412),
.A2(n_7406),
.B(n_7449),
.C(n_7421),
.Y(n_7529)
);

OAI211xp5_ASAP7_75t_L g7530 ( 
.A1(n_7418),
.A2(n_1463),
.B(n_1472),
.C(n_1455),
.Y(n_7530)
);

NOR2xp67_ASAP7_75t_L g7531 ( 
.A(n_7429),
.B(n_1456),
.Y(n_7531)
);

NAND2xp5_ASAP7_75t_L g7532 ( 
.A(n_7443),
.B(n_1456),
.Y(n_7532)
);

NAND3xp33_ASAP7_75t_SL g7533 ( 
.A(n_7452),
.B(n_1457),
.C(n_1458),
.Y(n_7533)
);

NAND2xp5_ASAP7_75t_L g7534 ( 
.A(n_7496),
.B(n_1459),
.Y(n_7534)
);

O2A1O1Ixp33_ASAP7_75t_L g7535 ( 
.A1(n_7407),
.A2(n_1461),
.B(n_1459),
.C(n_1460),
.Y(n_7535)
);

NAND3xp33_ASAP7_75t_L g7536 ( 
.A(n_7468),
.B(n_1460),
.C(n_1462),
.Y(n_7536)
);

NOR2xp33_ASAP7_75t_L g7537 ( 
.A(n_7403),
.B(n_1462),
.Y(n_7537)
);

OAI322xp33_ASAP7_75t_L g7538 ( 
.A1(n_7422),
.A2(n_1469),
.A3(n_1468),
.B1(n_1465),
.B2(n_1463),
.C1(n_1464),
.C2(n_1466),
.Y(n_7538)
);

NOR2xp33_ASAP7_75t_R g7539 ( 
.A(n_7431),
.B(n_7456),
.Y(n_7539)
);

O2A1O1Ixp33_ASAP7_75t_L g7540 ( 
.A1(n_7420),
.A2(n_1466),
.B(n_1464),
.C(n_1465),
.Y(n_7540)
);

O2A1O1Ixp33_ASAP7_75t_SL g7541 ( 
.A1(n_7414),
.A2(n_1471),
.B(n_1469),
.C(n_1470),
.Y(n_7541)
);

CKINVDCx5p33_ASAP7_75t_R g7542 ( 
.A(n_7494),
.Y(n_7542)
);

NAND2x1_ASAP7_75t_L g7543 ( 
.A(n_7475),
.B(n_1470),
.Y(n_7543)
);

AOI211xp5_ASAP7_75t_L g7544 ( 
.A1(n_7409),
.A2(n_7436),
.B(n_7444),
.C(n_7490),
.Y(n_7544)
);

OAI22xp5_ASAP7_75t_L g7545 ( 
.A1(n_7451),
.A2(n_1474),
.B1(n_1472),
.B2(n_1473),
.Y(n_7545)
);

NAND3xp33_ASAP7_75t_SL g7546 ( 
.A(n_7427),
.B(n_1473),
.C(n_1475),
.Y(n_7546)
);

OAI21xp5_ASAP7_75t_L g7547 ( 
.A1(n_7463),
.A2(n_1475),
.B(n_1476),
.Y(n_7547)
);

A2O1A1Ixp33_ASAP7_75t_L g7548 ( 
.A1(n_7461),
.A2(n_1480),
.B(n_1477),
.C(n_1478),
.Y(n_7548)
);

NAND4xp25_ASAP7_75t_L g7549 ( 
.A(n_7430),
.B(n_1480),
.C(n_1477),
.D(n_1478),
.Y(n_7549)
);

NAND3xp33_ASAP7_75t_SL g7550 ( 
.A(n_7467),
.B(n_1481),
.C(n_1482),
.Y(n_7550)
);

NAND2xp5_ASAP7_75t_SL g7551 ( 
.A(n_7446),
.B(n_1481),
.Y(n_7551)
);

AOI21xp5_ASAP7_75t_L g7552 ( 
.A1(n_7483),
.A2(n_1482),
.B(n_1483),
.Y(n_7552)
);

OAI21xp33_ASAP7_75t_SL g7553 ( 
.A1(n_7404),
.A2(n_1484),
.B(n_1485),
.Y(n_7553)
);

A2O1A1Ixp33_ASAP7_75t_L g7554 ( 
.A1(n_7479),
.A2(n_1486),
.B(n_1484),
.C(n_1485),
.Y(n_7554)
);

NAND3xp33_ASAP7_75t_SL g7555 ( 
.A(n_7424),
.B(n_1488),
.C(n_1489),
.Y(n_7555)
);

AND2x2_ASAP7_75t_L g7556 ( 
.A(n_7433),
.B(n_1488),
.Y(n_7556)
);

BUFx2_ASAP7_75t_L g7557 ( 
.A(n_7458),
.Y(n_7557)
);

OAI221xp5_ASAP7_75t_L g7558 ( 
.A1(n_7416),
.A2(n_1491),
.B1(n_1489),
.B2(n_1490),
.C(n_1492),
.Y(n_7558)
);

OAI22xp33_ASAP7_75t_L g7559 ( 
.A1(n_7419),
.A2(n_1495),
.B1(n_1496),
.B2(n_1493),
.Y(n_7559)
);

NOR2x1_ASAP7_75t_L g7560 ( 
.A(n_7405),
.B(n_1491),
.Y(n_7560)
);

NAND4xp75_ASAP7_75t_L g7561 ( 
.A(n_7488),
.B(n_7462),
.C(n_7469),
.D(n_7466),
.Y(n_7561)
);

INVx2_ASAP7_75t_L g7562 ( 
.A(n_7556),
.Y(n_7562)
);

INVxp67_ASAP7_75t_L g7563 ( 
.A(n_7504),
.Y(n_7563)
);

INVxp33_ASAP7_75t_SL g7564 ( 
.A(n_7528),
.Y(n_7564)
);

OAI22xp5_ASAP7_75t_L g7565 ( 
.A1(n_7520),
.A2(n_7485),
.B1(n_7423),
.B2(n_7495),
.Y(n_7565)
);

AOI31xp33_ASAP7_75t_L g7566 ( 
.A1(n_7525),
.A2(n_7471),
.A3(n_7480),
.B(n_7474),
.Y(n_7566)
);

OA22x2_ASAP7_75t_L g7567 ( 
.A1(n_7522),
.A2(n_7492),
.B1(n_7472),
.B2(n_7491),
.Y(n_7567)
);

INVx1_ASAP7_75t_L g7568 ( 
.A(n_7531),
.Y(n_7568)
);

OAI22xp5_ASAP7_75t_L g7569 ( 
.A1(n_7542),
.A2(n_7484),
.B1(n_7489),
.B2(n_7465),
.Y(n_7569)
);

AOI22xp5_ASAP7_75t_L g7570 ( 
.A1(n_7501),
.A2(n_7425),
.B1(n_7460),
.B2(n_7473),
.Y(n_7570)
);

AOI221xp5_ASAP7_75t_L g7571 ( 
.A1(n_7502),
.A2(n_7438),
.B1(n_7498),
.B2(n_1496),
.C(n_1493),
.Y(n_7571)
);

AOI22xp5_ASAP7_75t_L g7572 ( 
.A1(n_7499),
.A2(n_7516),
.B1(n_7514),
.B2(n_7513),
.Y(n_7572)
);

HB1xp67_ASAP7_75t_L g7573 ( 
.A(n_7543),
.Y(n_7573)
);

OAI22xp5_ASAP7_75t_L g7574 ( 
.A1(n_7536),
.A2(n_1498),
.B1(n_1495),
.B2(n_1497),
.Y(n_7574)
);

INVx1_ASAP7_75t_L g7575 ( 
.A(n_7500),
.Y(n_7575)
);

INVx2_ASAP7_75t_L g7576 ( 
.A(n_7561),
.Y(n_7576)
);

INVx1_ASAP7_75t_L g7577 ( 
.A(n_7532),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_7534),
.Y(n_7578)
);

BUFx2_ASAP7_75t_L g7579 ( 
.A(n_7553),
.Y(n_7579)
);

INVx1_ASAP7_75t_L g7580 ( 
.A(n_7509),
.Y(n_7580)
);

OAI22xp5_ASAP7_75t_L g7581 ( 
.A1(n_7521),
.A2(n_1499),
.B1(n_1497),
.B2(n_1498),
.Y(n_7581)
);

AOI221xp5_ASAP7_75t_L g7582 ( 
.A1(n_7505),
.A2(n_1502),
.B1(n_1500),
.B2(n_1501),
.C(n_1504),
.Y(n_7582)
);

AOI221xp5_ASAP7_75t_L g7583 ( 
.A1(n_7503),
.A2(n_1505),
.B1(n_1500),
.B2(n_1501),
.C(n_1507),
.Y(n_7583)
);

AOI22xp5_ASAP7_75t_L g7584 ( 
.A1(n_7549),
.A2(n_1509),
.B1(n_1505),
.B2(n_1508),
.Y(n_7584)
);

INVx1_ASAP7_75t_L g7585 ( 
.A(n_7523),
.Y(n_7585)
);

AOI22xp5_ASAP7_75t_L g7586 ( 
.A1(n_7533),
.A2(n_7507),
.B1(n_7550),
.B2(n_7506),
.Y(n_7586)
);

INVxp33_ASAP7_75t_L g7587 ( 
.A(n_7539),
.Y(n_7587)
);

OAI22xp5_ASAP7_75t_L g7588 ( 
.A1(n_7548),
.A2(n_1511),
.B1(n_1508),
.B2(n_1510),
.Y(n_7588)
);

A2O1A1Ixp33_ASAP7_75t_SL g7589 ( 
.A1(n_7544),
.A2(n_1513),
.B(n_1511),
.C(n_1512),
.Y(n_7589)
);

AOI22xp5_ASAP7_75t_L g7590 ( 
.A1(n_7529),
.A2(n_1515),
.B1(n_1512),
.B2(n_1514),
.Y(n_7590)
);

INVx2_ASAP7_75t_L g7591 ( 
.A(n_7557),
.Y(n_7591)
);

INVx1_ASAP7_75t_L g7592 ( 
.A(n_7541),
.Y(n_7592)
);

BUFx2_ASAP7_75t_L g7593 ( 
.A(n_7560),
.Y(n_7593)
);

INVx1_ASAP7_75t_L g7594 ( 
.A(n_7540),
.Y(n_7594)
);

NAND2xp5_ASAP7_75t_L g7595 ( 
.A(n_7537),
.B(n_1514),
.Y(n_7595)
);

INVx1_ASAP7_75t_L g7596 ( 
.A(n_7551),
.Y(n_7596)
);

OA22x2_ASAP7_75t_L g7597 ( 
.A1(n_7515),
.A2(n_1517),
.B1(n_1515),
.B2(n_1516),
.Y(n_7597)
);

OAI22x1_ASAP7_75t_L g7598 ( 
.A1(n_7508),
.A2(n_1518),
.B1(n_1516),
.B2(n_1517),
.Y(n_7598)
);

OA22x2_ASAP7_75t_L g7599 ( 
.A1(n_7547),
.A2(n_1522),
.B1(n_1520),
.B2(n_1521),
.Y(n_7599)
);

AOI221xp5_ASAP7_75t_L g7600 ( 
.A1(n_7519),
.A2(n_1522),
.B1(n_1520),
.B2(n_1521),
.C(n_1523),
.Y(n_7600)
);

AOI221xp5_ASAP7_75t_L g7601 ( 
.A1(n_7511),
.A2(n_1525),
.B1(n_1523),
.B2(n_1524),
.C(n_1526),
.Y(n_7601)
);

AOI221x1_ASAP7_75t_L g7602 ( 
.A1(n_7598),
.A2(n_7526),
.B1(n_7555),
.B2(n_7552),
.C(n_7546),
.Y(n_7602)
);

OAI21xp5_ASAP7_75t_SL g7603 ( 
.A1(n_7587),
.A2(n_7518),
.B(n_7510),
.Y(n_7603)
);

INVx1_ASAP7_75t_L g7604 ( 
.A(n_7579),
.Y(n_7604)
);

AOI33xp33_ASAP7_75t_L g7605 ( 
.A1(n_7576),
.A2(n_7592),
.A3(n_7594),
.B1(n_7568),
.B2(n_7585),
.B3(n_7572),
.Y(n_7605)
);

AOI221xp5_ASAP7_75t_SL g7606 ( 
.A1(n_7566),
.A2(n_7512),
.B1(n_7517),
.B2(n_7535),
.C(n_7527),
.Y(n_7606)
);

AOI321xp33_ASAP7_75t_L g7607 ( 
.A1(n_7565),
.A2(n_7524),
.A3(n_7545),
.B1(n_7554),
.B2(n_7558),
.C(n_7530),
.Y(n_7607)
);

OAI211xp5_ASAP7_75t_SL g7608 ( 
.A1(n_7563),
.A2(n_7559),
.B(n_7538),
.C(n_1527),
.Y(n_7608)
);

AOI211xp5_ASAP7_75t_L g7609 ( 
.A1(n_7582),
.A2(n_1527),
.B(n_1524),
.C(n_1525),
.Y(n_7609)
);

AOI22xp5_ASAP7_75t_L g7610 ( 
.A1(n_7564),
.A2(n_1530),
.B1(n_1528),
.B2(n_1529),
.Y(n_7610)
);

INVx1_ASAP7_75t_L g7611 ( 
.A(n_7573),
.Y(n_7611)
);

NAND4xp25_ASAP7_75t_L g7612 ( 
.A(n_7570),
.B(n_1531),
.C(n_1528),
.D(n_1529),
.Y(n_7612)
);

AOI31xp33_ASAP7_75t_L g7613 ( 
.A1(n_7571),
.A2(n_1533),
.A3(n_1531),
.B(n_1532),
.Y(n_7613)
);

AOI221xp5_ASAP7_75t_L g7614 ( 
.A1(n_7569),
.A2(n_1534),
.B1(n_1532),
.B2(n_1533),
.C(n_1535),
.Y(n_7614)
);

NAND2xp5_ASAP7_75t_SL g7615 ( 
.A(n_7583),
.B(n_1536),
.Y(n_7615)
);

AOI221x1_ASAP7_75t_L g7616 ( 
.A1(n_7581),
.A2(n_1538),
.B1(n_1536),
.B2(n_1537),
.C(n_1540),
.Y(n_7616)
);

OAI222xp33_ASAP7_75t_L g7617 ( 
.A1(n_7586),
.A2(n_1541),
.B1(n_1543),
.B2(n_1538),
.C1(n_1540),
.C2(n_1542),
.Y(n_7617)
);

OA22x2_ASAP7_75t_SL g7618 ( 
.A1(n_7596),
.A2(n_1543),
.B1(n_1541),
.B2(n_1542),
.Y(n_7618)
);

NAND3xp33_ASAP7_75t_L g7619 ( 
.A(n_7601),
.B(n_1544),
.C(n_1545),
.Y(n_7619)
);

INVx1_ASAP7_75t_L g7620 ( 
.A(n_7597),
.Y(n_7620)
);

NAND2xp5_ASAP7_75t_SL g7621 ( 
.A(n_7590),
.B(n_1544),
.Y(n_7621)
);

OAI21xp33_ASAP7_75t_L g7622 ( 
.A1(n_7575),
.A2(n_1545),
.B(n_1546),
.Y(n_7622)
);

OAI211xp5_ASAP7_75t_SL g7623 ( 
.A1(n_7580),
.A2(n_1548),
.B(n_1546),
.C(n_1547),
.Y(n_7623)
);

AOI221x1_ASAP7_75t_L g7624 ( 
.A1(n_7588),
.A2(n_1549),
.B1(n_1547),
.B2(n_1548),
.C(n_1550),
.Y(n_7624)
);

AOI221xp5_ASAP7_75t_L g7625 ( 
.A1(n_7593),
.A2(n_1553),
.B1(n_1549),
.B2(n_1552),
.C(n_1554),
.Y(n_7625)
);

AOI31xp33_ASAP7_75t_L g7626 ( 
.A1(n_7604),
.A2(n_7562),
.A3(n_7591),
.B(n_7578),
.Y(n_7626)
);

OR2x2_ASAP7_75t_L g7627 ( 
.A(n_7611),
.B(n_7589),
.Y(n_7627)
);

AOI221xp5_ASAP7_75t_L g7628 ( 
.A1(n_7613),
.A2(n_7577),
.B1(n_7574),
.B2(n_7600),
.C(n_7584),
.Y(n_7628)
);

AOI211xp5_ASAP7_75t_L g7629 ( 
.A1(n_7603),
.A2(n_7595),
.B(n_7567),
.C(n_7599),
.Y(n_7629)
);

AOI22xp5_ASAP7_75t_L g7630 ( 
.A1(n_7620),
.A2(n_1556),
.B1(n_1552),
.B2(n_1553),
.Y(n_7630)
);

NOR3xp33_ASAP7_75t_L g7631 ( 
.A(n_7606),
.B(n_7605),
.C(n_7608),
.Y(n_7631)
);

O2A1O1Ixp5_ASAP7_75t_L g7632 ( 
.A1(n_7615),
.A2(n_1558),
.B(n_1556),
.C(n_1557),
.Y(n_7632)
);

AOI222xp33_ASAP7_75t_L g7633 ( 
.A1(n_7621),
.A2(n_1559),
.B1(n_1562),
.B2(n_1557),
.C1(n_1558),
.C2(n_1561),
.Y(n_7633)
);

OAI221xp5_ASAP7_75t_L g7634 ( 
.A1(n_7607),
.A2(n_1563),
.B1(n_1561),
.B2(n_1562),
.C(n_1564),
.Y(n_7634)
);

AOI22xp5_ASAP7_75t_L g7635 ( 
.A1(n_7623),
.A2(n_7619),
.B1(n_7612),
.B2(n_7609),
.Y(n_7635)
);

OAI21xp33_ASAP7_75t_L g7636 ( 
.A1(n_7622),
.A2(n_1564),
.B(n_1565),
.Y(n_7636)
);

NOR3xp33_ASAP7_75t_L g7637 ( 
.A(n_7614),
.B(n_1565),
.C(n_1566),
.Y(n_7637)
);

NOR2xp33_ASAP7_75t_L g7638 ( 
.A(n_7617),
.B(n_1566),
.Y(n_7638)
);

AO22x2_ASAP7_75t_L g7639 ( 
.A1(n_7602),
.A2(n_7616),
.B1(n_7624),
.B2(n_7618),
.Y(n_7639)
);

NAND2xp5_ASAP7_75t_L g7640 ( 
.A(n_7610),
.B(n_7625),
.Y(n_7640)
);

OAI21xp33_ASAP7_75t_L g7641 ( 
.A1(n_7605),
.A2(n_1567),
.B(n_1568),
.Y(n_7641)
);

NOR2x1_ASAP7_75t_L g7642 ( 
.A(n_7612),
.B(n_1568),
.Y(n_7642)
);

OAI211xp5_ASAP7_75t_L g7643 ( 
.A1(n_7603),
.A2(n_1572),
.B(n_1569),
.C(n_1571),
.Y(n_7643)
);

AND3x1_ASAP7_75t_L g7644 ( 
.A(n_7605),
.B(n_1569),
.C(n_1571),
.Y(n_7644)
);

OAI32xp33_ASAP7_75t_L g7645 ( 
.A1(n_7627),
.A2(n_1574),
.A3(n_1572),
.B1(n_1573),
.B2(n_1575),
.Y(n_7645)
);

AOI222xp33_ASAP7_75t_L g7646 ( 
.A1(n_7641),
.A2(n_1577),
.B1(n_1579),
.B2(n_1573),
.C1(n_1576),
.C2(n_1578),
.Y(n_7646)
);

AOI21xp5_ASAP7_75t_L g7647 ( 
.A1(n_7626),
.A2(n_7639),
.B(n_7640),
.Y(n_7647)
);

AND2x2_ASAP7_75t_L g7648 ( 
.A(n_7639),
.B(n_1577),
.Y(n_7648)
);

INVx1_ASAP7_75t_L g7649 ( 
.A(n_7644),
.Y(n_7649)
);

NOR2x1p5_ASAP7_75t_L g7650 ( 
.A(n_7634),
.B(n_1578),
.Y(n_7650)
);

INVx2_ASAP7_75t_L g7651 ( 
.A(n_7632),
.Y(n_7651)
);

NAND3xp33_ASAP7_75t_L g7652 ( 
.A(n_7631),
.B(n_1580),
.C(n_1581),
.Y(n_7652)
);

AO211x2_ASAP7_75t_L g7653 ( 
.A1(n_7637),
.A2(n_7643),
.B(n_7629),
.C(n_7642),
.Y(n_7653)
);

AOI221xp5_ASAP7_75t_L g7654 ( 
.A1(n_7638),
.A2(n_1583),
.B1(n_1581),
.B2(n_1582),
.C(n_1584),
.Y(n_7654)
);

A2O1A1Ixp33_ASAP7_75t_L g7655 ( 
.A1(n_7636),
.A2(n_1585),
.B(n_1582),
.C(n_1583),
.Y(n_7655)
);

NAND3xp33_ASAP7_75t_L g7656 ( 
.A(n_7633),
.B(n_1585),
.C(n_1587),
.Y(n_7656)
);

INVx1_ASAP7_75t_L g7657 ( 
.A(n_7630),
.Y(n_7657)
);

NAND3xp33_ASAP7_75t_SL g7658 ( 
.A(n_7628),
.B(n_1587),
.C(n_1588),
.Y(n_7658)
);

AND2x2_ASAP7_75t_L g7659 ( 
.A(n_7648),
.B(n_7635),
.Y(n_7659)
);

INVx1_ASAP7_75t_L g7660 ( 
.A(n_7652),
.Y(n_7660)
);

INVx1_ASAP7_75t_SL g7661 ( 
.A(n_7651),
.Y(n_7661)
);

NAND3x2_ASAP7_75t_L g7662 ( 
.A(n_7649),
.B(n_7657),
.C(n_7653),
.Y(n_7662)
);

O2A1O1Ixp33_ASAP7_75t_L g7663 ( 
.A1(n_7658),
.A2(n_1591),
.B(n_1589),
.C(n_1590),
.Y(n_7663)
);

AND2x4_ASAP7_75t_L g7664 ( 
.A(n_7659),
.B(n_7650),
.Y(n_7664)
);

AOI22xp5_ASAP7_75t_L g7665 ( 
.A1(n_7661),
.A2(n_7654),
.B1(n_7656),
.B2(n_7647),
.Y(n_7665)
);

OAI211xp5_ASAP7_75t_L g7666 ( 
.A1(n_7662),
.A2(n_7646),
.B(n_7655),
.C(n_7645),
.Y(n_7666)
);

NOR4xp75_ASAP7_75t_L g7667 ( 
.A(n_7663),
.B(n_1594),
.C(n_1591),
.D(n_1592),
.Y(n_7667)
);

NOR3xp33_ASAP7_75t_L g7668 ( 
.A(n_7666),
.B(n_7660),
.C(n_1594),
.Y(n_7668)
);

AND4x2_ASAP7_75t_L g7669 ( 
.A(n_7667),
.B(n_1597),
.C(n_1595),
.D(n_1596),
.Y(n_7669)
);

OAI22x1_ASAP7_75t_L g7670 ( 
.A1(n_7669),
.A2(n_7665),
.B1(n_7664),
.B2(n_1599),
.Y(n_7670)
);

INVx1_ASAP7_75t_L g7671 ( 
.A(n_7668),
.Y(n_7671)
);

OAI22x1_ASAP7_75t_L g7672 ( 
.A1(n_7671),
.A2(n_1599),
.B1(n_1596),
.B2(n_1597),
.Y(n_7672)
);

INVx1_ASAP7_75t_L g7673 ( 
.A(n_7670),
.Y(n_7673)
);

NOR2x2_ASAP7_75t_L g7674 ( 
.A(n_7673),
.B(n_1600),
.Y(n_7674)
);

AOI22xp5_ASAP7_75t_L g7675 ( 
.A1(n_7672),
.A2(n_1602),
.B1(n_1600),
.B2(n_1601),
.Y(n_7675)
);

AOI22xp33_ASAP7_75t_L g7676 ( 
.A1(n_7675),
.A2(n_1605),
.B1(n_1602),
.B2(n_1604),
.Y(n_7676)
);

NOR2xp33_ASAP7_75t_L g7677 ( 
.A(n_7676),
.B(n_7674),
.Y(n_7677)
);

INVx2_ASAP7_75t_SL g7678 ( 
.A(n_7676),
.Y(n_7678)
);

AOI22xp5_ASAP7_75t_L g7679 ( 
.A1(n_7677),
.A2(n_1606),
.B1(n_1604),
.B2(n_1605),
.Y(n_7679)
);

XNOR2x1_ASAP7_75t_L g7680 ( 
.A(n_7678),
.B(n_1607),
.Y(n_7680)
);

AOI21xp5_ASAP7_75t_L g7681 ( 
.A1(n_7680),
.A2(n_1608),
.B(n_1609),
.Y(n_7681)
);

NOR2xp67_ASAP7_75t_L g7682 ( 
.A(n_7679),
.B(n_1608),
.Y(n_7682)
);

INVx1_ASAP7_75t_L g7683 ( 
.A(n_7682),
.Y(n_7683)
);

INVx2_ASAP7_75t_L g7684 ( 
.A(n_7681),
.Y(n_7684)
);

OR2x6_ASAP7_75t_L g7685 ( 
.A(n_7684),
.B(n_1609),
.Y(n_7685)
);

AOI21xp33_ASAP7_75t_L g7686 ( 
.A1(n_7685),
.A2(n_7683),
.B(n_1611),
.Y(n_7686)
);

AOI211xp5_ASAP7_75t_L g7687 ( 
.A1(n_7686),
.A2(n_1614),
.B(n_1612),
.C(n_1613),
.Y(n_7687)
);


endmodule