module real_aes_6962_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_119;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_729;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g184 ( .A1(n_0), .A2(n_185), .B(n_186), .C(n_190), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_1), .B(n_179), .Y(n_192) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g129 ( .A(n_2), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_3), .B(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_4), .A2(n_173), .B(n_479), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_5), .A2(n_153), .B(n_170), .C(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_6), .A2(n_173), .B(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_7), .B(n_179), .Y(n_485) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_8), .A2(n_145), .B(n_267), .Y(n_266) );
AND2x6_ASAP7_75t_L g170 ( .A(n_9), .B(n_171), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_10), .A2(n_153), .B(n_170), .C(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g576 ( .A(n_11), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_12), .B(n_41), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_13), .B(n_189), .Y(n_525) );
INVx1_ASAP7_75t_L g150 ( .A(n_14), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_15), .B(n_164), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_16), .A2(n_165), .B(n_534), .C(n_536), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_17), .B(n_179), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_18), .B(n_207), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_19), .A2(n_153), .B(n_199), .C(n_206), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_20), .A2(n_188), .B(n_241), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_21), .B(n_189), .Y(n_507) );
AOI222xp33_ASAP7_75t_L g454 ( .A1(n_22), .A2(n_455), .B1(n_724), .B2(n_725), .C1(n_734), .C2(n_738), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_23), .B(n_189), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_24), .Y(n_503) );
INVx1_ASAP7_75t_L g473 ( .A(n_25), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_26), .A2(n_153), .B(n_206), .C(n_270), .Y(n_269) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_27), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_28), .A2(n_105), .B1(n_116), .B2(n_741), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_29), .Y(n_521) );
INVx1_ASAP7_75t_L g497 ( .A(n_30), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_31), .A2(n_173), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_32), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g155 ( .A(n_33), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_34), .A2(n_168), .B(n_222), .C(n_223), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_35), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_36), .A2(n_188), .B(n_482), .C(n_484), .Y(n_481) );
INVxp67_ASAP7_75t_L g498 ( .A(n_37), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_38), .B(n_272), .Y(n_271) );
CKINVDCx14_ASAP7_75t_R g480 ( .A(n_39), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_40), .A2(n_153), .B(n_206), .C(n_472), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_42), .A2(n_190), .B(n_574), .C(n_575), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_43), .B(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_44), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_45), .B(n_164), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_46), .B(n_173), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_47), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_48), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_49), .A2(n_168), .B(n_222), .C(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g187 ( .A(n_50), .Y(n_187) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_51), .A2(n_67), .B1(n_132), .B2(n_133), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_51), .Y(n_133) );
INVx1_ASAP7_75t_L g251 ( .A(n_52), .Y(n_251) );
INVx1_ASAP7_75t_L g541 ( .A(n_53), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_54), .B(n_173), .Y(n_248) );
OAI22xp5_ASAP7_75t_SL g135 ( .A1(n_55), .A2(n_72), .B1(n_136), .B2(n_137), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_55), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_56), .Y(n_211) );
CKINVDCx14_ASAP7_75t_R g572 ( .A(n_57), .Y(n_572) );
INVx1_ASAP7_75t_L g171 ( .A(n_58), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_59), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_60), .B(n_179), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_61), .A2(n_160), .B(n_205), .C(n_262), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_62), .A2(n_71), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_62), .Y(n_731) );
INVx1_ASAP7_75t_L g149 ( .A(n_63), .Y(n_149) );
INVx1_ASAP7_75t_SL g483 ( .A(n_64), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_65), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_66), .B(n_164), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_67), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_67), .B(n_179), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_68), .B(n_165), .Y(n_238) );
INVx1_ASAP7_75t_L g506 ( .A(n_69), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_70), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_71), .Y(n_732) );
INVx1_ASAP7_75t_L g137 ( .A(n_72), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_73), .B(n_201), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_74), .A2(n_153), .B(n_158), .C(n_168), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_75), .Y(n_260) );
INVx1_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_77), .A2(n_173), .B(n_571), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_78), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_79), .A2(n_173), .B(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_80), .A2(n_197), .B(n_493), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_81), .Y(n_470) );
INVx1_ASAP7_75t_L g532 ( .A(n_82), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_83), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_83), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_84), .B(n_203), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_85), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_86), .A2(n_173), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g535 ( .A(n_87), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_88), .A2(n_726), .B1(n_727), .B2(n_733), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_88), .Y(n_726) );
INVx2_ASAP7_75t_L g147 ( .A(n_89), .Y(n_147) );
INVx1_ASAP7_75t_L g524 ( .A(n_90), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_91), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_92), .B(n_189), .Y(n_239) );
INVx2_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
OR2x2_ASAP7_75t_L g126 ( .A(n_93), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g459 ( .A(n_93), .B(n_128), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_94), .A2(n_153), .B(n_168), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_95), .B(n_173), .Y(n_220) );
INVx1_ASAP7_75t_L g224 ( .A(n_96), .Y(n_224) );
INVxp67_ASAP7_75t_L g263 ( .A(n_97), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_98), .B(n_145), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_99), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g159 ( .A(n_100), .Y(n_159) );
INVx1_ASAP7_75t_L g234 ( .A(n_101), .Y(n_234) );
INVx2_ASAP7_75t_L g544 ( .A(n_102), .Y(n_544) );
AND2x2_ASAP7_75t_L g253 ( .A(n_103), .B(n_209), .Y(n_253) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g741 ( .A(n_106), .Y(n_741) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_114), .Y(n_108) );
OR2x2_ASAP7_75t_L g723 ( .A(n_110), .B(n_128), .Y(n_723) );
NOR2x2_ASAP7_75t_L g740 ( .A(n_110), .B(n_127), .Y(n_740) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g128 ( .A(n_115), .B(n_129), .Y(n_128) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_453), .Y(n_116) );
BUFx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_118), .B(n_450), .C(n_454), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_130), .B(n_450), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_126), .Y(n_452) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_134), .B1(n_448), .B2(n_449), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_131), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_134), .Y(n_449) );
XNOR2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_138), .Y(n_134) );
INVx1_ASAP7_75t_L g456 ( .A(n_138), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_138), .A2(n_461), .B1(n_735), .B2(n_736), .Y(n_734) );
OR3x1_ASAP7_75t_L g138 ( .A(n_139), .B(n_356), .C(n_405), .Y(n_138) );
NAND5xp2_ASAP7_75t_L g139 ( .A(n_140), .B(n_290), .C(n_319), .D(n_327), .E(n_342), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_213), .B(n_229), .C(n_274), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_193), .Y(n_141) );
AND2x2_ASAP7_75t_L g285 ( .A(n_142), .B(n_282), .Y(n_285) );
AND2x2_ASAP7_75t_L g318 ( .A(n_142), .B(n_194), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_142), .B(n_217), .Y(n_411) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_178), .Y(n_142) );
INVx2_ASAP7_75t_L g216 ( .A(n_143), .Y(n_216) );
BUFx2_ASAP7_75t_L g385 ( .A(n_143), .Y(n_385) );
AO21x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_151), .B(n_176), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_144), .B(n_177), .Y(n_176) );
INVx3_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_144), .B(n_228), .Y(n_227) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_144), .A2(n_233), .B(n_243), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_144), .B(n_476), .Y(n_475) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_144), .A2(n_502), .B(n_509), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_144), .B(n_527), .Y(n_526) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_145), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_145), .A2(n_268), .B(n_269), .Y(n_267) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g245 ( .A(n_146), .Y(n_245) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x2_ASAP7_75t_SL g209 ( .A(n_147), .B(n_148), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_172), .Y(n_151) );
INVx5_ASAP7_75t_L g183 ( .A(n_153), .Y(n_183) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
BUFx3_ASAP7_75t_L g191 ( .A(n_154), .Y(n_191) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
INVx1_ASAP7_75t_L g242 ( .A(n_155), .Y(n_242) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_157), .Y(n_162) );
INVx3_ASAP7_75t_L g165 ( .A(n_157), .Y(n_165) );
AND2x2_ASAP7_75t_L g174 ( .A(n_157), .B(n_175), .Y(n_174) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
INVx1_ASAP7_75t_L g272 ( .A(n_157), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_163), .C(n_166), .Y(n_158) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_161), .A2(n_164), .B1(n_497), .B2(n_498), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_161), .B(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_161), .B(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g201 ( .A(n_162), .Y(n_201) );
INVx2_ASAP7_75t_L g185 ( .A(n_164), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_164), .B(n_263), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_164), .A2(n_204), .B(n_473), .C(n_474), .Y(n_472) );
INVx5_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_165), .B(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx3_ASAP7_75t_L g484 ( .A(n_167), .Y(n_484) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_SL g181 ( .A1(n_169), .A2(n_182), .B(n_183), .C(n_184), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_169), .A2(n_183), .B(n_260), .C(n_261), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_169), .A2(n_183), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_169), .A2(n_183), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_169), .A2(n_183), .B(n_532), .C(n_533), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_SL g540 ( .A1(n_169), .A2(n_183), .B(n_541), .C(n_542), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_SL g571 ( .A1(n_169), .A2(n_183), .B(n_572), .C(n_573), .Y(n_571) );
INVx4_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
AND2x4_ASAP7_75t_L g173 ( .A(n_170), .B(n_174), .Y(n_173) );
BUFx3_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g235 ( .A(n_170), .B(n_174), .Y(n_235) );
BUFx2_ASAP7_75t_L g197 ( .A(n_173), .Y(n_197) );
INVx1_ASAP7_75t_L g205 ( .A(n_175), .Y(n_205) );
AND2x2_ASAP7_75t_L g193 ( .A(n_178), .B(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g283 ( .A(n_178), .Y(n_283) );
AND2x2_ASAP7_75t_L g369 ( .A(n_178), .B(n_282), .Y(n_369) );
AND2x2_ASAP7_75t_L g424 ( .A(n_178), .B(n_216), .Y(n_424) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_192), .Y(n_178) );
INVx2_ASAP7_75t_L g222 ( .A(n_183), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_188), .B(n_483), .Y(n_482) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g574 ( .A(n_189), .Y(n_574) );
INVx2_ASAP7_75t_L g508 ( .A(n_190), .Y(n_508) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_191), .Y(n_226) );
INVx1_ASAP7_75t_L g536 ( .A(n_191), .Y(n_536) );
INVx1_ASAP7_75t_L g341 ( .A(n_193), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_193), .B(n_217), .Y(n_388) );
INVx5_ASAP7_75t_L g282 ( .A(n_194), .Y(n_282) );
AND2x4_ASAP7_75t_L g303 ( .A(n_194), .B(n_283), .Y(n_303) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_194), .Y(n_325) );
AND2x2_ASAP7_75t_L g400 ( .A(n_194), .B(n_385), .Y(n_400) );
AND2x2_ASAP7_75t_L g403 ( .A(n_194), .B(n_218), .Y(n_403) );
OR2x6_ASAP7_75t_L g194 ( .A(n_195), .B(n_210), .Y(n_194) );
AOI21xp5_ASAP7_75t_SL g195 ( .A1(n_196), .A2(n_198), .B(n_207), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_202), .B(n_204), .Y(n_199) );
INVx2_ASAP7_75t_L g203 ( .A(n_201), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_203), .A2(n_224), .B(n_225), .C(n_226), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_203), .A2(n_226), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_203), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
O2A1O1Ixp5_ASAP7_75t_L g523 ( .A1(n_203), .A2(n_508), .B(n_524), .C(n_525), .Y(n_523) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_205), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_208), .B(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g212 ( .A(n_209), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_209), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_209), .A2(n_248), .B(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_209), .A2(n_235), .B(n_470), .C(n_471), .Y(n_469) );
OA21x2_ASAP7_75t_L g569 ( .A1(n_209), .A2(n_570), .B(n_577), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_212), .A2(n_520), .B(n_526), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_213), .B(n_283), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_213), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
AND2x2_ASAP7_75t_L g308 ( .A(n_215), .B(n_283), .Y(n_308) );
AND2x2_ASAP7_75t_L g326 ( .A(n_215), .B(n_218), .Y(n_326) );
INVx1_ASAP7_75t_L g346 ( .A(n_215), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_215), .B(n_282), .Y(n_391) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_215), .Y(n_433) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_216), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_217), .B(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_217), .Y(n_335) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_217), .A2(n_278), .B(n_339), .C(n_341), .Y(n_338) );
AND2x2_ASAP7_75t_L g345 ( .A(n_217), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g354 ( .A(n_217), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g358 ( .A(n_217), .B(n_282), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_217), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g373 ( .A(n_217), .B(n_283), .Y(n_373) );
AND2x2_ASAP7_75t_L g423 ( .A(n_217), .B(n_424), .Y(n_423) );
INVx5_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx2_ASAP7_75t_L g287 ( .A(n_218), .Y(n_287) );
AND2x2_ASAP7_75t_L g328 ( .A(n_218), .B(n_281), .Y(n_328) );
AND2x2_ASAP7_75t_L g340 ( .A(n_218), .B(n_315), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_218), .B(n_369), .Y(n_387) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_227), .Y(n_218) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_254), .Y(n_229) );
INVx1_ASAP7_75t_L g276 ( .A(n_230), .Y(n_276) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_246), .Y(n_230) );
OR2x2_ASAP7_75t_L g278 ( .A(n_231), .B(n_246), .Y(n_278) );
NAND3xp33_ASAP7_75t_L g284 ( .A(n_231), .B(n_285), .C(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_231), .B(n_256), .Y(n_295) );
OR2x2_ASAP7_75t_L g310 ( .A(n_231), .B(n_298), .Y(n_310) );
AND2x2_ASAP7_75t_L g316 ( .A(n_231), .B(n_265), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_231), .B(n_447), .Y(n_446) );
INVx5_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_232), .B(n_256), .Y(n_313) );
AND2x2_ASAP7_75t_L g352 ( .A(n_232), .B(n_266), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_232), .B(n_265), .Y(n_380) );
OR2x2_ASAP7_75t_L g383 ( .A(n_232), .B(n_265), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_236), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_235), .A2(n_503), .B(n_504), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_235), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_240), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_240), .A2(n_271), .B(n_273), .Y(n_270) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx2_ASAP7_75t_L g491 ( .A(n_245), .Y(n_491) );
INVx5_ASAP7_75t_SL g298 ( .A(n_246), .Y(n_298) );
OR2x2_ASAP7_75t_L g304 ( .A(n_246), .B(n_255), .Y(n_304) );
AND2x2_ASAP7_75t_L g320 ( .A(n_246), .B(n_321), .Y(n_320) );
AOI321xp33_ASAP7_75t_L g327 ( .A1(n_246), .A2(n_328), .A3(n_329), .B1(n_330), .B2(n_336), .C(n_338), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_246), .B(n_254), .Y(n_337) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_246), .Y(n_350) );
OR2x2_ASAP7_75t_L g397 ( .A(n_246), .B(n_295), .Y(n_397) );
AND2x2_ASAP7_75t_L g419 ( .A(n_246), .B(n_316), .Y(n_419) );
AND2x2_ASAP7_75t_L g438 ( .A(n_246), .B(n_256), .Y(n_438) );
OR2x6_ASAP7_75t_L g246 ( .A(n_247), .B(n_253), .Y(n_246) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_265), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_256), .B(n_265), .Y(n_279) );
AND2x2_ASAP7_75t_L g288 ( .A(n_256), .B(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g315 ( .A(n_256), .Y(n_315) );
AND2x2_ASAP7_75t_L g321 ( .A(n_256), .B(n_316), .Y(n_321) );
INVxp67_ASAP7_75t_L g351 ( .A(n_256), .Y(n_351) );
OR2x2_ASAP7_75t_L g393 ( .A(n_256), .B(n_298), .Y(n_393) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_264), .Y(n_256) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_257), .A2(n_478), .B(n_485), .Y(n_477) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_257), .A2(n_530), .B(n_537), .Y(n_529) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_257), .A2(n_539), .B(n_545), .Y(n_538) );
OR2x2_ASAP7_75t_L g275 ( .A(n_265), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_SL g289 ( .A(n_265), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_265), .B(n_278), .Y(n_322) );
AND2x2_ASAP7_75t_L g371 ( .A(n_265), .B(n_315), .Y(n_371) );
AND2x2_ASAP7_75t_L g409 ( .A(n_265), .B(n_298), .Y(n_409) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_266), .B(n_298), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_277), .B(n_280), .C(n_284), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_275), .A2(n_277), .B1(n_402), .B2(n_404), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_277), .A2(n_300), .B1(n_355), .B2(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_SL g429 ( .A(n_278), .Y(n_429) );
INVx1_ASAP7_75t_SL g329 ( .A(n_279), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_281), .B(n_301), .Y(n_331) );
AOI222xp33_ASAP7_75t_L g342 ( .A1(n_281), .A2(n_322), .B1(n_329), .B2(n_343), .C1(n_347), .C2(n_353), .Y(n_342) );
AND2x2_ASAP7_75t_L g432 ( .A(n_281), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_282), .B(n_302), .Y(n_377) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_282), .Y(n_414) );
AND2x2_ASAP7_75t_L g417 ( .A(n_282), .B(n_326), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_282), .B(n_433), .Y(n_443) );
INVx1_ASAP7_75t_L g334 ( .A(n_283), .Y(n_334) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_283), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_L g425 ( .A1(n_285), .A2(n_426), .B(n_427), .C(n_430), .Y(n_425) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND3xp33_ASAP7_75t_L g348 ( .A(n_287), .B(n_349), .C(n_352), .Y(n_348) );
OR2x2_ASAP7_75t_L g376 ( .A(n_287), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_287), .B(n_303), .Y(n_404) );
OR2x2_ASAP7_75t_L g309 ( .A(n_289), .B(n_310), .Y(n_309) );
AOI211xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_293), .B(n_299), .C(n_311), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_292), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g398 ( .A(n_293), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_294), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g312 ( .A(n_297), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_298), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g366 ( .A(n_298), .B(n_316), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_298), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_298), .B(n_315), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_304), .B1(n_305), .B2(n_309), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_301), .B(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_303), .B(n_345), .Y(n_344) );
OAI221xp5_ASAP7_75t_SL g367 ( .A1(n_304), .A2(n_368), .B1(n_370), .B2(n_372), .C(n_374), .Y(n_367) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AND2x2_ASAP7_75t_L g422 ( .A(n_307), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g435 ( .A(n_307), .B(n_424), .Y(n_435) );
INVx1_ASAP7_75t_L g355 ( .A(n_308), .Y(n_355) );
INVx1_ASAP7_75t_L g426 ( .A(n_309), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_310), .A2(n_393), .B(n_416), .Y(n_415) );
AOI21xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_314), .B(n_317), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI21xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_322), .B(n_323), .Y(n_319) );
INVx1_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_321), .A2(n_407), .B1(n_410), .B2(n_412), .C(n_415), .Y(n_406) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_329), .A2(n_419), .B1(n_420), .B2(n_422), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g395 ( .A(n_331), .Y(n_395) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR2xp67_ASAP7_75t_SL g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g399 ( .A(n_335), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g364 ( .A(n_340), .Y(n_364) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_345), .B(n_369), .Y(n_421) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_351), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g437 ( .A(n_352), .B(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g444 ( .A(n_352), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI211xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_359), .B(n_360), .C(n_394), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI211xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B(n_367), .C(n_386), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g447 ( .A(n_371), .Y(n_447) );
AND2x2_ASAP7_75t_L g384 ( .A(n_373), .B(n_385), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_382), .B2(n_384), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
OR2x2_ASAP7_75t_L g392 ( .A(n_380), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g445 ( .A(n_381), .Y(n_445) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI31xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .A3(n_389), .B(n_392), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI211xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_398), .C(n_401), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_403), .Y(n_402) );
NAND5xp2_ASAP7_75t_L g405 ( .A(n_406), .B(n_418), .C(n_425), .D(n_439), .E(n_442), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_417), .A2(n_443), .B1(n_444), .B2(n_446), .Y(n_442) );
INVx1_ASAP7_75t_SL g441 ( .A(n_419), .Y(n_441) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_434), .B(n_436), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_457), .B1(n_460), .B2(n_723), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g735 ( .A(n_458), .Y(n_735) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR3x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_634), .C(n_681), .Y(n_461) );
NAND3xp33_ASAP7_75t_SL g462 ( .A(n_463), .B(n_580), .C(n_605), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_518), .B1(n_546), .B2(n_549), .C(n_557), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_486), .B(n_511), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_466), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_466), .B(n_562), .Y(n_678) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .Y(n_466) );
AND2x2_ASAP7_75t_L g548 ( .A(n_467), .B(n_517), .Y(n_548) );
AND2x2_ASAP7_75t_L g598 ( .A(n_467), .B(n_516), .Y(n_598) );
AND2x2_ASAP7_75t_L g619 ( .A(n_467), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g624 ( .A(n_467), .B(n_591), .Y(n_624) );
OR2x2_ASAP7_75t_L g632 ( .A(n_467), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g704 ( .A(n_467), .B(n_500), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_467), .B(n_653), .Y(n_718) );
INVx3_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g563 ( .A(n_468), .B(n_477), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_468), .B(n_500), .Y(n_564) );
AND2x4_ASAP7_75t_L g586 ( .A(n_468), .B(n_517), .Y(n_586) );
AND2x2_ASAP7_75t_L g616 ( .A(n_468), .B(n_488), .Y(n_616) );
AND2x2_ASAP7_75t_L g625 ( .A(n_468), .B(n_615), .Y(n_625) );
AND2x2_ASAP7_75t_L g641 ( .A(n_468), .B(n_501), .Y(n_641) );
OR2x2_ASAP7_75t_L g650 ( .A(n_468), .B(n_633), .Y(n_650) );
AND2x2_ASAP7_75t_L g656 ( .A(n_468), .B(n_591), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_468), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g670 ( .A(n_468), .B(n_513), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_468), .B(n_559), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_468), .B(n_620), .Y(n_709) );
OR2x6_ASAP7_75t_L g468 ( .A(n_469), .B(n_475), .Y(n_468) );
INVx2_ASAP7_75t_L g517 ( .A(n_477), .Y(n_517) );
AND2x2_ASAP7_75t_L g615 ( .A(n_477), .B(n_500), .Y(n_615) );
AND2x2_ASAP7_75t_L g620 ( .A(n_477), .B(n_501), .Y(n_620) );
INVx1_ASAP7_75t_L g676 ( .A(n_477), .Y(n_676) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g585 ( .A(n_487), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_500), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_488), .B(n_548), .Y(n_547) );
BUFx3_ASAP7_75t_L g562 ( .A(n_488), .Y(n_562) );
OR2x2_ASAP7_75t_L g633 ( .A(n_488), .B(n_500), .Y(n_633) );
OR2x2_ASAP7_75t_L g694 ( .A(n_488), .B(n_601), .Y(n_694) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_492), .B(n_499), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_490), .A2(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g514 ( .A(n_492), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_499), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_500), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g653 ( .A(n_500), .B(n_513), .Y(n_653) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g592 ( .A(n_501), .Y(n_592) );
INVx1_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_512), .A2(n_698), .B1(n_702), .B2(n_705), .C(n_706), .Y(n_697) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_516), .Y(n_512) );
INVx1_ASAP7_75t_SL g560 ( .A(n_513), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_513), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g692 ( .A(n_513), .B(n_548), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_516), .B(n_562), .Y(n_684) );
AND2x2_ASAP7_75t_L g591 ( .A(n_517), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g595 ( .A(n_518), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_518), .B(n_601), .Y(n_631) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
AND2x2_ASAP7_75t_L g556 ( .A(n_519), .B(n_529), .Y(n_556) );
INVx4_ASAP7_75t_L g568 ( .A(n_519), .Y(n_568) );
BUFx3_ASAP7_75t_L g611 ( .A(n_519), .Y(n_611) );
AND3x2_ASAP7_75t_L g626 ( .A(n_519), .B(n_627), .C(n_628), .Y(n_626) );
AND2x2_ASAP7_75t_L g708 ( .A(n_528), .B(n_622), .Y(n_708) );
AND2x2_ASAP7_75t_L g716 ( .A(n_528), .B(n_601), .Y(n_716) );
INVx1_ASAP7_75t_SL g721 ( .A(n_528), .Y(n_721) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .Y(n_528) );
INVx1_ASAP7_75t_SL g579 ( .A(n_529), .Y(n_579) );
AND2x2_ASAP7_75t_L g602 ( .A(n_529), .B(n_568), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_529), .B(n_552), .Y(n_604) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_529), .Y(n_644) );
OR2x2_ASAP7_75t_L g649 ( .A(n_529), .B(n_568), .Y(n_649) );
INVx2_ASAP7_75t_L g554 ( .A(n_538), .Y(n_554) );
AND2x2_ASAP7_75t_L g589 ( .A(n_538), .B(n_569), .Y(n_589) );
OR2x2_ASAP7_75t_L g609 ( .A(n_538), .B(n_569), .Y(n_609) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_538), .Y(n_629) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AOI21xp33_ASAP7_75t_L g679 ( .A1(n_547), .A2(n_588), .B(n_680), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g715 ( .A1(n_549), .A2(n_559), .A3(n_586), .B1(n_716), .B2(n_717), .C1(n_719), .C2(n_722), .Y(n_715) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_555), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_551), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_552), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g578 ( .A(n_553), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g646 ( .A(n_554), .B(n_568), .Y(n_646) );
AND2x2_ASAP7_75t_L g713 ( .A(n_554), .B(n_569), .Y(n_713) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g654 ( .A(n_556), .B(n_608), .Y(n_654) );
AOI31xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .A3(n_564), .B(n_565), .Y(n_557) );
AND2x2_ASAP7_75t_L g613 ( .A(n_559), .B(n_591), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_559), .B(n_583), .Y(n_695) );
AND2x2_ASAP7_75t_L g714 ( .A(n_559), .B(n_619), .Y(n_714) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_562), .B(n_591), .Y(n_603) );
NAND2x1p5_ASAP7_75t_L g637 ( .A(n_562), .B(n_620), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_562), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_562), .B(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_563), .B(n_620), .Y(n_652) );
INVx1_ASAP7_75t_L g696 ( .A(n_563), .Y(n_696) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_578), .Y(n_566) );
INVxp67_ASAP7_75t_L g648 ( .A(n_567), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_568), .B(n_579), .Y(n_584) );
INVx1_ASAP7_75t_L g690 ( .A(n_568), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_568), .B(n_667), .Y(n_701) );
BUFx3_ASAP7_75t_L g601 ( .A(n_569), .Y(n_601) );
AND2x2_ASAP7_75t_L g627 ( .A(n_569), .B(n_579), .Y(n_627) );
INVx2_ASAP7_75t_L g667 ( .A(n_569), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_578), .B(n_700), .Y(n_699) );
AOI211xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_585), .B(n_587), .C(n_596), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI21xp33_ASAP7_75t_L g630 ( .A1(n_582), .A2(n_631), .B(n_632), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_583), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_583), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g663 ( .A(n_584), .B(n_609), .Y(n_663) );
INVx3_ASAP7_75t_L g594 ( .A(n_586), .Y(n_594) );
OAI22xp5_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_590), .B1(n_593), .B2(n_595), .Y(n_587) );
OAI21xp5_ASAP7_75t_SL g612 ( .A1(n_589), .A2(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g638 ( .A(n_589), .B(n_602), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_589), .B(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g593 ( .A(n_592), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g662 ( .A(n_592), .Y(n_662) );
OAI21xp5_ASAP7_75t_SL g606 ( .A1(n_593), .A2(n_607), .B(n_612), .Y(n_606) );
OAI22xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_599), .B1(n_603), .B2(n_604), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_598), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g622 ( .A(n_601), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_601), .B(n_644), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_617), .C(n_630), .Y(n_605) );
OAI22xp5_ASAP7_75t_SL g672 ( .A1(n_607), .A2(n_673), .B1(n_677), .B2(n_678), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g677 ( .A(n_609), .B(n_610), .Y(n_677) );
AND2x2_ASAP7_75t_L g685 ( .A(n_610), .B(n_666), .Y(n_685) );
CKINVDCx16_ASAP7_75t_R g610 ( .A(n_611), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_SL g693 ( .A1(n_611), .A2(n_694), .B(n_695), .C(n_696), .Y(n_693) );
OR2x2_ASAP7_75t_L g720 ( .A(n_611), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B(n_623), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_619), .A2(n_656), .B(n_657), .C(n_660), .Y(n_655) );
OAI21xp33_ASAP7_75t_SL g623 ( .A1(n_624), .A2(n_625), .B(n_626), .Y(n_623) );
AND2x2_ASAP7_75t_L g688 ( .A(n_627), .B(n_646), .Y(n_688) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g666 ( .A(n_629), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g671 ( .A(n_631), .Y(n_671) );
NAND3xp33_ASAP7_75t_SL g634 ( .A(n_635), .B(n_655), .C(n_668), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B(n_639), .C(n_647), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g705 ( .A(n_642), .Y(n_705) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g665 ( .A(n_644), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_644), .B(n_713), .Y(n_712) );
INVxp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B(n_650), .C(n_651), .Y(n_647) );
INVx2_ASAP7_75t_SL g659 ( .A(n_649), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_650), .A2(n_661), .B1(n_663), .B2(n_664), .Y(n_660) );
OAI21xp33_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_653), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_672), .C(n_679), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVxp33_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g722 ( .A(n_676), .Y(n_722) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_682), .B(n_697), .C(n_710), .D(n_715), .Y(n_681) );
AOI211xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_685), .B(n_686), .C(n_693), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_691), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_687), .A2(n_707), .B(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_694), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .Y(n_710) );
INVxp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g737 ( .A(n_723), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
CKINVDCx16_ASAP7_75t_R g733 ( .A(n_727), .Y(n_733) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
endmodule