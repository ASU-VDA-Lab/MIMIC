module fake_jpeg_10646_n_87 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_87);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_87;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_27),
.Y(n_32)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_10),
.B(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_10),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_30),
.C(n_17),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_22),
.C(n_26),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_18),
.B(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_56),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_18),
.B(n_13),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_19),
.B(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_9),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_19),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_60),
.Y(n_70)
);

OAI22x1_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_26),
.B1(n_21),
.B2(n_24),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_21),
.B1(n_19),
.B2(n_12),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_48),
.B(n_57),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_68),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_56),
.B(n_2),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_70),
.B1(n_64),
.B2(n_58),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_58),
.C(n_59),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_50),
.C(n_24),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_76),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_75),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_50),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_27),
.C(n_24),
.Y(n_76)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_69),
.B(n_24),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_72),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_79),
.B(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_81),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_27),
.C(n_9),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_80),
.C(n_5),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_3),
.B(n_6),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_7),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_84),
.Y(n_87)
);


endmodule