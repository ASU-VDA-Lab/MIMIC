module fake_aes_9830_n_948 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_948);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_948;
wire n_117;
wire n_663;
wire n_791;
wire n_707;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_858;
wire n_604;
wire n_603;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_228;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_568;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_805;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_889;
wire n_635;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_926;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_666;
wire n_799;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_899;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_723;
wire n_597;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g111 ( .A(n_87), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_25), .Y(n_112) );
BUFx5_ASAP7_75t_L g113 ( .A(n_110), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_22), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_85), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_41), .Y(n_116) );
BUFx10_ASAP7_75t_L g117 ( .A(n_20), .Y(n_117) );
BUFx2_ASAP7_75t_SL g118 ( .A(n_103), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_54), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_3), .Y(n_120) );
BUFx10_ASAP7_75t_L g121 ( .A(n_78), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_19), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_101), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_95), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_59), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_37), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_97), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_105), .Y(n_128) );
CKINVDCx14_ASAP7_75t_R g129 ( .A(n_96), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_93), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_84), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_7), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_38), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_102), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_56), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_14), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_98), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_24), .Y(n_139) );
INVxp67_ASAP7_75t_L g140 ( .A(n_14), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_90), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_76), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_5), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_92), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_40), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_36), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_42), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_61), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_49), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_55), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_45), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_31), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_18), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_113), .B(n_0), .Y(n_154) );
BUFx12f_ASAP7_75t_L g155 ( .A(n_121), .Y(n_155) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_111), .A2(n_0), .B(n_1), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_123), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g158 ( .A(n_129), .Y(n_158) );
NOR2x1_ASAP7_75t_L g159 ( .A(n_139), .B(n_1), .Y(n_159) );
BUFx12f_ASAP7_75t_L g160 ( .A(n_121), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_139), .B(n_2), .Y(n_161) );
INVxp33_ASAP7_75t_SL g162 ( .A(n_145), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_123), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_139), .Y(n_164) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_112), .A2(n_50), .B(n_108), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_113), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_140), .B(n_2), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_120), .B(n_3), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_143), .B(n_4), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_113), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_113), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_127), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_123), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_115), .A2(n_4), .B(n_5), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_133), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_122), .B(n_6), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_166), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_155), .B(n_117), .Y(n_179) );
OR2x6_ASAP7_75t_L g180 ( .A(n_155), .B(n_118), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_172), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_158), .B(n_133), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_169), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_155), .B(n_117), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_164), .B(n_116), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_164), .B(n_119), .Y(n_187) );
AND3x2_ASAP7_75t_L g188 ( .A(n_169), .B(n_114), .C(n_152), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_166), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_172), .B(n_125), .Y(n_191) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_161), .B(n_113), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_166), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_172), .B(n_126), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_172), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_158), .B(n_121), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_170), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_162), .A2(n_153), .B1(n_137), .B2(n_150), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_160), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_170), .Y(n_200) );
AOI21x1_ASAP7_75t_L g201 ( .A1(n_170), .A2(n_136), .B(n_131), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_170), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_169), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_171), .Y(n_204) );
NAND2xp33_ASAP7_75t_SL g205 ( .A(n_161), .B(n_137), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_157), .Y(n_206) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_160), .Y(n_207) );
OR2x6_ASAP7_75t_L g208 ( .A(n_160), .B(n_130), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_171), .Y(n_209) );
BUFx8_ASAP7_75t_SL g210 ( .A(n_160), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_162), .B(n_135), .Y(n_211) );
OAI22x1_ASAP7_75t_L g212 ( .A1(n_156), .A2(n_153), .B1(n_151), .B2(n_150), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_171), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_169), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_169), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_156), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_156), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_174), .B(n_142), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_154), .A2(n_149), .B(n_147), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_157), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
AOI22xp33_ASAP7_75t_SL g224 ( .A1(n_176), .A2(n_117), .B1(n_132), .B2(n_128), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_156), .Y(n_225) );
INVxp33_ASAP7_75t_SL g226 ( .A(n_167), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_216), .A2(n_156), .B1(n_175), .B2(n_154), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_211), .B(n_167), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_211), .B(n_128), .Y(n_230) );
NAND2xp33_ASAP7_75t_L g231 ( .A(n_199), .B(n_113), .Y(n_231) );
OR2x6_ASAP7_75t_L g232 ( .A(n_180), .B(n_176), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_203), .B(n_132), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_203), .B(n_134), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_203), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_217), .B(n_146), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_180), .B(n_168), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_226), .B(n_168), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_216), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_203), .B(n_134), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_199), .B(n_138), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_208), .A2(n_177), .B1(n_159), .B2(n_175), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_184), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_217), .B(n_113), .Y(n_244) );
NOR3xp33_ASAP7_75t_L g245 ( .A(n_224), .B(n_198), .C(n_205), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_179), .B(n_177), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_184), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_179), .B(n_138), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_184), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_185), .B(n_141), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_184), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_185), .B(n_141), .Y(n_252) );
NOR3x1_ASAP7_75t_L g253 ( .A(n_198), .B(n_165), .C(n_174), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_180), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_215), .Y(n_255) );
NAND3xp33_ASAP7_75t_L g256 ( .A(n_217), .B(n_175), .C(n_159), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_180), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_180), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_210), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_189), .B(n_144), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_195), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_195), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_225), .A2(n_165), .B(n_175), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_215), .B(n_144), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_189), .B(n_151), .Y(n_265) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_215), .B(n_175), .Y(n_266) );
AND2x6_ASAP7_75t_L g267 ( .A(n_215), .B(n_127), .Y(n_267) );
INVxp33_ASAP7_75t_L g268 ( .A(n_207), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_195), .Y(n_269) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_178), .Y(n_270) );
NOR2xp67_ASAP7_75t_L g271 ( .A(n_212), .B(n_8), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_188), .B(n_124), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_186), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_188), .B(n_175), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_217), .B(n_165), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_218), .B(n_123), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_186), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_182), .B(n_9), .Y(n_278) );
INVx8_ASAP7_75t_L g279 ( .A(n_180), .Y(n_279) );
NOR2x1p5_ASAP7_75t_L g280 ( .A(n_182), .B(n_148), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_187), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_187), .B(n_148), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_218), .B(n_148), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_227), .B(n_148), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_196), .B(n_26), .Y(n_285) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_208), .B(n_157), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_208), .B(n_157), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_191), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_181), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_208), .B(n_27), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_208), .B(n_157), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_237), .A2(n_208), .B1(n_225), .B2(n_224), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_286), .B(n_227), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_235), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_245), .A2(n_212), .B1(n_192), .B2(n_221), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_236), .A2(n_225), .B(n_181), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_238), .B(n_191), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_238), .B(n_219), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_273), .A2(n_281), .B1(n_277), .B2(n_288), .Y(n_299) );
AOI21x1_ASAP7_75t_L g300 ( .A1(n_275), .A2(n_201), .B(n_194), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_246), .B(n_194), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_236), .A2(n_181), .B(n_190), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_263), .A2(n_190), .B(n_197), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_243), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_246), .B(n_178), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_237), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_276), .A2(n_200), .B(n_197), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_279), .B(n_201), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_235), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_229), .B(n_221), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_247), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_230), .B(n_221), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_248), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_276), .A2(n_200), .B(n_221), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_249), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_270), .B(n_183), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_250), .B(n_183), .Y(n_317) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_239), .A2(n_204), .B(n_183), .C(n_193), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_274), .A2(n_213), .B(n_202), .C(n_204), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_254), .B(n_193), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_279), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_252), .B(n_193), .Y(n_322) );
BUFx8_ASAP7_75t_L g323 ( .A(n_259), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_283), .A2(n_213), .B(n_202), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_237), .A2(n_209), .B1(n_202), .B2(n_204), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_264), .B(n_209), .Y(n_326) );
INVx4_ASAP7_75t_L g327 ( .A(n_279), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_257), .B(n_209), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_251), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_268), .B(n_213), .Y(n_330) );
OAI21xp5_ASAP7_75t_L g331 ( .A1(n_256), .A2(n_214), .B(n_222), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_232), .A2(n_214), .B1(n_163), .B2(n_173), .Y(n_332) );
A2O1A1Ixp33_ASAP7_75t_SL g333 ( .A1(n_290), .A2(n_214), .B(n_222), .C(n_220), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_283), .A2(n_223), .B(n_222), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_264), .B(n_9), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_232), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_260), .B(n_10), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_265), .B(n_10), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_261), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_241), .B(n_11), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_244), .A2(n_223), .B(n_220), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_233), .B(n_11), .Y(n_342) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_271), .A2(n_173), .B(n_163), .C(n_157), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_330), .Y(n_344) );
BUFx8_ASAP7_75t_L g345 ( .A(n_336), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_312), .A2(n_284), .B(n_275), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_298), .A2(n_290), .B(n_242), .C(n_285), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_321), .B(n_258), .Y(n_348) );
AOI21x1_ASAP7_75t_L g349 ( .A1(n_300), .A2(n_282), .B(n_284), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_303), .A2(n_291), .B(n_287), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_321), .B(n_268), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_299), .B(n_278), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_296), .A2(n_244), .B(n_255), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_343), .B(n_295), .C(n_332), .Y(n_354) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_331), .A2(n_266), .B(n_289), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_299), .B(n_232), .Y(n_356) );
AO31x2_ASAP7_75t_L g357 ( .A1(n_343), .A2(n_285), .A3(n_253), .B(n_269), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_305), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_297), .B(n_280), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_293), .A2(n_240), .B(n_234), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_293), .A2(n_228), .B(n_266), .Y(n_361) );
AOI21x1_ASAP7_75t_L g362 ( .A1(n_335), .A2(n_262), .B(n_223), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_292), .A2(n_267), .B1(n_272), .B2(n_231), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_304), .Y(n_364) );
O2A1O1Ixp33_ASAP7_75t_SL g365 ( .A1(n_333), .A2(n_267), .B(n_220), .C(n_228), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_314), .A2(n_267), .B(n_173), .Y(n_366) );
OA22x2_ASAP7_75t_L g367 ( .A1(n_306), .A2(n_267), .B1(n_13), .B2(n_15), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_327), .Y(n_368) );
BUFx12f_ASAP7_75t_L g369 ( .A(n_323), .Y(n_369) );
OR2x6_ASAP7_75t_L g370 ( .A(n_327), .B(n_308), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_310), .A2(n_206), .B(n_267), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_313), .B(n_12), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_298), .A2(n_173), .B1(n_163), .B2(n_206), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g374 ( .A1(n_310), .A2(n_173), .B(n_163), .C(n_206), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_301), .B(n_12), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_366), .A2(n_341), .B(n_319), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_356), .B(n_337), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_350), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_349), .A2(n_324), .B(n_334), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_364), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_370), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_358), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_344), .Y(n_383) );
INVx3_ASAP7_75t_L g384 ( .A(n_370), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_356), .A2(n_322), .B1(n_338), .B2(n_340), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_362), .A2(n_342), .B(n_325), .Y(n_386) );
AOI22x1_ASAP7_75t_L g387 ( .A1(n_371), .A2(n_302), .B1(n_339), .B2(n_307), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_369), .Y(n_388) );
AOI22x1_ASAP7_75t_L g389 ( .A1(n_360), .A2(n_339), .B1(n_329), .B2(n_315), .Y(n_389) );
OAI21x1_ASAP7_75t_L g390 ( .A1(n_361), .A2(n_326), .B(n_328), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_352), .Y(n_391) );
AO21x2_ASAP7_75t_L g392 ( .A1(n_354), .A2(n_333), .B(n_318), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_348), .Y(n_393) );
OAI21x1_ASAP7_75t_L g394 ( .A1(n_346), .A2(n_328), .B(n_320), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_355), .Y(n_395) );
AOI21x1_ASAP7_75t_L g396 ( .A1(n_354), .A2(n_308), .B(n_320), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_353), .A2(n_317), .B(n_311), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_345), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_367), .A2(n_316), .B(n_322), .Y(n_399) );
NOR2x1_ASAP7_75t_R g400 ( .A(n_351), .B(n_323), .Y(n_400) );
AO21x1_ASAP7_75t_L g401 ( .A1(n_375), .A2(n_309), .B(n_294), .Y(n_401) );
OAI21x1_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_308), .B(n_318), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_363), .B(n_339), .Y(n_403) );
OAI21x1_ASAP7_75t_L g404 ( .A1(n_373), .A2(n_339), .B(n_173), .Y(n_404) );
OAI21x1_ASAP7_75t_L g405 ( .A1(n_365), .A2(n_173), .B(n_163), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_380), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_380), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_380), .B(n_357), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_377), .B(n_347), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_382), .A2(n_372), .B1(n_359), .B2(n_368), .C(n_374), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_383), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_378), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_393), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_381), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_383), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_384), .B(n_370), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_382), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_378), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_384), .B(n_357), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_393), .B(n_377), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_393), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_378), .Y(n_422) );
BUFx2_ASAP7_75t_L g423 ( .A(n_381), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_391), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_400), .B(n_345), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_377), .B(n_357), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_384), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_402), .Y(n_428) );
AO21x2_ASAP7_75t_L g429 ( .A1(n_401), .A2(n_173), .B(n_163), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_391), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_395), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_397), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_384), .B(n_63), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_395), .Y(n_434) );
OAI21x1_ASAP7_75t_L g435 ( .A1(n_405), .A2(n_348), .B(n_163), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_397), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_385), .B(n_13), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_403), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_398), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_397), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_402), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_402), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_400), .Y(n_443) );
OAI21x1_ASAP7_75t_L g444 ( .A1(n_405), .A2(n_163), .B(n_206), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_385), .B(n_15), .Y(n_445) );
OR2x6_ASAP7_75t_L g446 ( .A(n_403), .B(n_16), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_401), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_399), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_394), .B(n_396), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_403), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_401), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_388), .B(n_16), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_426), .B(n_392), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_406), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_419), .B(n_396), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_407), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_426), .B(n_392), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_424), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_424), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_437), .B(n_399), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_420), .B(n_392), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_430), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_420), .B(n_392), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_430), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
AND2x2_ASAP7_75t_SL g468 ( .A(n_438), .B(n_437), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_409), .B(n_399), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_446), .B(n_395), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_411), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_415), .B(n_394), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_412), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_425), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_421), .Y(n_476) );
BUFx3_ASAP7_75t_L g477 ( .A(n_421), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_415), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_409), .B(n_403), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_408), .B(n_390), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_417), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_421), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_413), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_413), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_408), .B(n_390), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_419), .B(n_405), .Y(n_486) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_418), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_417), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_432), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_419), .B(n_390), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_419), .B(n_394), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_441), .B(n_404), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_441), .B(n_442), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_443), .A2(n_387), .B1(n_389), .B2(n_386), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_450), .B(n_404), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_432), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_436), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_442), .B(n_404), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_436), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_440), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_443), .A2(n_387), .B1(n_389), .B2(n_386), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_445), .A2(n_386), .B1(n_376), .B2(n_379), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_428), .B(n_376), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_414), .B(n_376), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_445), .B(n_17), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_440), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_413), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_412), .Y(n_508) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_418), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_414), .B(n_17), .Y(n_510) );
INVx4_ASAP7_75t_R g511 ( .A(n_427), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_428), .B(n_379), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_422), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_447), .B(n_451), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_422), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_422), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_431), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_423), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_450), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_447), .B(n_379), .Y(n_520) );
INVxp67_ASAP7_75t_SL g521 ( .A(n_423), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_431), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_416), .B(n_18), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_431), .Y(n_524) );
INVx4_ASAP7_75t_L g525 ( .A(n_446), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_434), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_451), .B(n_19), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_450), .B(n_20), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_450), .B(n_21), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_434), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_438), .B(n_66), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_463), .B(n_448), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_463), .B(n_449), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_467), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_459), .B(n_434), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_469), .B(n_416), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_525), .B(n_449), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_469), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_467), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_472), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_525), .B(n_449), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_465), .B(n_449), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_459), .B(n_427), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_518), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_472), .B(n_416), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_478), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_465), .B(n_429), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_477), .Y(n_548) );
INVx4_ASAP7_75t_L g549 ( .A(n_525), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_453), .B(n_429), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_474), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_525), .B(n_446), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_478), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_453), .B(n_429), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_474), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_481), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_481), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_480), .B(n_429), .Y(n_558) );
NAND4xp25_ASAP7_75t_L g559 ( .A(n_523), .B(n_452), .C(n_410), .D(n_416), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_480), .B(n_446), .Y(n_560) );
BUFx2_ASAP7_75t_SL g561 ( .A(n_477), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_485), .B(n_446), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_476), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_485), .B(n_433), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_479), .B(n_433), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_488), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_468), .A2(n_410), .B1(n_433), .B2(n_439), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_508), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_488), .B(n_433), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_456), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_479), .B(n_435), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_460), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_470), .B(n_435), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_482), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_491), .B(n_514), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_456), .Y(n_576) );
NOR2xp33_ASAP7_75t_R g577 ( .A(n_468), .B(n_21), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_491), .B(n_435), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_514), .B(n_444), .Y(n_579) );
INVxp67_ASAP7_75t_SL g580 ( .A(n_487), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_457), .B(n_444), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_460), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_484), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_461), .Y(n_584) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_495), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_461), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_527), .B(n_22), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_468), .B(n_477), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_490), .B(n_444), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_470), .B(n_23), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_490), .B(n_23), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_464), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_509), .B(n_24), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_493), .B(n_28), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_464), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_527), .B(n_29), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_466), .B(n_30), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_483), .B(n_206), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_457), .B(n_32), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_508), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_458), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_493), .B(n_33), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_462), .B(n_34), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_457), .B(n_35), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_524), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_524), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_483), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_466), .B(n_39), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_458), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_520), .B(n_43), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_457), .B(n_44), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_507), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_454), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_520), .B(n_46), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_475), .B(n_47), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_521), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_454), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_455), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_512), .B(n_48), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_512), .B(n_51), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_455), .B(n_52), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_503), .B(n_53), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_503), .B(n_57), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_483), .B(n_206), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_492), .B(n_58), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_492), .B(n_60), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_498), .B(n_62), .Y(n_627) );
BUFx2_ASAP7_75t_L g628 ( .A(n_471), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_489), .Y(n_629) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_510), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_498), .B(n_64), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_526), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_489), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_526), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_530), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_530), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_496), .B(n_65), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_538), .Y(n_638) );
AND2x4_ASAP7_75t_L g639 ( .A(n_549), .B(n_471), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_630), .B(n_497), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_629), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_544), .B(n_497), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_538), .Y(n_643) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_580), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_559), .B(n_505), .Y(n_645) );
INVx3_ASAP7_75t_SL g646 ( .A(n_549), .Y(n_646) );
AND2x4_ASAP7_75t_SL g647 ( .A(n_549), .B(n_531), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_629), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_575), .B(n_519), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_575), .B(n_513), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_546), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_546), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_590), .B(n_506), .Y(n_653) );
INVxp33_ASAP7_75t_L g654 ( .A(n_577), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_564), .B(n_519), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_548), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_633), .Y(n_657) );
NAND2xp33_ASAP7_75t_SL g658 ( .A(n_588), .B(n_511), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_564), .B(n_519), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_533), .B(n_519), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_616), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_533), .B(n_495), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_563), .Y(n_663) );
AND3x2_ASAP7_75t_L g664 ( .A(n_552), .B(n_529), .C(n_528), .Y(n_664) );
NOR2xp67_ASAP7_75t_R g665 ( .A(n_628), .B(n_511), .Y(n_665) );
INVxp67_ASAP7_75t_SL g666 ( .A(n_574), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g667 ( .A1(n_567), .A2(n_510), .B(n_529), .Y(n_667) );
BUFx3_ASAP7_75t_L g668 ( .A(n_583), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_542), .B(n_495), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_612), .B(n_522), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_542), .B(n_495), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_560), .B(n_486), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_552), .B(n_531), .Y(n_673) );
NOR2xp67_ASAP7_75t_L g674 ( .A(n_552), .B(n_531), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_553), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_553), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_633), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_534), .Y(n_678) );
NAND2x1p5_ASAP7_75t_L g679 ( .A(n_599), .B(n_531), .Y(n_679) );
OR2x2_ASAP7_75t_L g680 ( .A(n_573), .B(n_513), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_590), .B(n_496), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_570), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_560), .B(n_486), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_562), .B(n_486), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_562), .B(n_486), .Y(n_685) );
AND2x4_ASAP7_75t_L g686 ( .A(n_537), .B(n_500), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_591), .B(n_500), .Y(n_687) );
INVx2_ASAP7_75t_SL g688 ( .A(n_607), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_591), .B(n_506), .Y(n_689) );
INVx4_ASAP7_75t_L g690 ( .A(n_599), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_556), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_532), .B(n_499), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_570), .Y(n_693) );
NAND2x1p5_ASAP7_75t_L g694 ( .A(n_599), .B(n_528), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_572), .B(n_499), .Y(n_695) );
AND2x4_ASAP7_75t_L g696 ( .A(n_537), .B(n_504), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_556), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_582), .B(n_473), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_576), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_584), .B(n_522), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_576), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_586), .B(n_517), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_532), .B(n_517), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_561), .Y(n_704) );
INVx4_ASAP7_75t_L g705 ( .A(n_604), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_578), .B(n_516), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_592), .B(n_516), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_573), .B(n_515), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_535), .B(n_515), .Y(n_709) );
INVxp33_ASAP7_75t_L g710 ( .A(n_604), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_578), .B(n_504), .Y(n_711) );
BUFx2_ASAP7_75t_L g712 ( .A(n_604), .Y(n_712) );
INVx2_ASAP7_75t_SL g713 ( .A(n_585), .Y(n_713) );
INVxp67_ASAP7_75t_SL g714 ( .A(n_593), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_619), .B(n_502), .Y(n_715) );
INVx2_ASAP7_75t_SL g716 ( .A(n_585), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_535), .B(n_502), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_595), .B(n_501), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_601), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_601), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_619), .B(n_494), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_620), .B(n_67), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_620), .B(n_68), .Y(n_723) );
NAND2x1_ASAP7_75t_SL g724 ( .A(n_611), .B(n_69), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_540), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_557), .B(n_70), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_566), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_534), .Y(n_728) );
AND2x6_ASAP7_75t_SL g729 ( .A(n_615), .B(n_71), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_611), .B(n_72), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_539), .Y(n_731) );
BUFx2_ASAP7_75t_L g732 ( .A(n_611), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_539), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_622), .B(n_73), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_571), .B(n_74), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_622), .B(n_75), .Y(n_736) );
OR2x2_ASAP7_75t_L g737 ( .A(n_571), .B(n_77), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_609), .Y(n_738) );
AND2x4_ASAP7_75t_L g739 ( .A(n_537), .B(n_541), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_613), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_541), .B(n_79), .Y(n_741) );
NAND2x1_ASAP7_75t_L g742 ( .A(n_541), .B(n_80), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_623), .B(n_81), .Y(n_743) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_593), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_661), .Y(n_745) );
NOR2x1_ASAP7_75t_L g746 ( .A(n_730), .B(n_561), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_661), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_662), .B(n_547), .Y(n_748) );
INVxp67_ASAP7_75t_SL g749 ( .A(n_644), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_669), .B(n_547), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_671), .B(n_554), .Y(n_751) );
AND2x2_ASAP7_75t_SL g752 ( .A(n_705), .B(n_690), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_678), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_644), .B(n_554), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_672), .B(n_550), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_683), .B(n_550), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_650), .B(n_543), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_646), .B(n_628), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_666), .B(n_617), .Y(n_759) );
AND3x1_ASAP7_75t_L g760 ( .A(n_667), .B(n_587), .C(n_594), .Y(n_760) );
OR2x2_ASAP7_75t_L g761 ( .A(n_680), .B(n_543), .Y(n_761) );
INVxp67_ASAP7_75t_SL g762 ( .A(n_678), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_666), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_642), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_725), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_727), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_692), .B(n_618), .Y(n_767) );
INVxp67_ASAP7_75t_L g768 ( .A(n_668), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_738), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_668), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_684), .B(n_558), .Y(n_771) );
OR2x2_ASAP7_75t_L g772 ( .A(n_708), .B(n_558), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_640), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_641), .B(n_600), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_641), .B(n_600), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_638), .Y(n_776) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_663), .Y(n_777) );
INVx2_ASAP7_75t_SL g778 ( .A(n_656), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_685), .B(n_585), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_648), .B(n_606), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_649), .B(n_585), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_648), .B(n_606), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_643), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_651), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_654), .B(n_545), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_660), .B(n_585), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_652), .Y(n_787) );
OR2x2_ASAP7_75t_L g788 ( .A(n_703), .B(n_565), .Y(n_788) );
INVx2_ASAP7_75t_SL g789 ( .A(n_688), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_711), .B(n_589), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_663), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_675), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_657), .B(n_605), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_717), .B(n_565), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_676), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_688), .B(n_589), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_691), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_697), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_699), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_657), .B(n_555), .Y(n_800) );
OR2x2_ASAP7_75t_L g801 ( .A(n_709), .B(n_536), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_701), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_655), .B(n_659), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_719), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_677), .B(n_551), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_677), .B(n_551), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_696), .B(n_579), .Y(n_807) );
INVxp67_ASAP7_75t_L g808 ( .A(n_714), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g809 ( .A(n_646), .B(n_581), .Y(n_809) );
INVx1_ASAP7_75t_SL g810 ( .A(n_704), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_670), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_682), .Y(n_812) );
OR2x2_ASAP7_75t_L g813 ( .A(n_706), .B(n_687), .Y(n_813) );
OR2x2_ASAP7_75t_L g814 ( .A(n_689), .B(n_579), .Y(n_814) );
OR2x2_ASAP7_75t_L g815 ( .A(n_653), .B(n_632), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_728), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_682), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_654), .B(n_569), .Y(n_818) );
INVx2_ASAP7_75t_SL g819 ( .A(n_647), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_696), .B(n_581), .Y(n_820) );
OR2x2_ASAP7_75t_L g821 ( .A(n_681), .B(n_696), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_714), .B(n_632), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_693), .B(n_555), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_693), .B(n_605), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_730), .A2(n_598), .B(n_624), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_720), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_720), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_645), .B(n_596), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_753), .Y(n_829) );
AOI32xp33_ASAP7_75t_L g830 ( .A1(n_760), .A2(n_658), .A3(n_710), .B1(n_647), .B2(n_705), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_745), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_808), .B(n_744), .Y(n_832) );
OAI21xp33_ASAP7_75t_L g833 ( .A1(n_808), .A2(n_645), .B(n_744), .Y(n_833) );
INVxp67_ASAP7_75t_L g834 ( .A(n_749), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_747), .B(n_718), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_759), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_752), .A2(n_705), .B1(n_690), .B2(n_679), .Y(n_837) );
O2A1O1Ixp33_ASAP7_75t_L g838 ( .A1(n_749), .A2(n_742), .B(n_673), .C(n_608), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_759), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_763), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_764), .B(n_715), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_777), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_791), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_815), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_816), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_765), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_822), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_766), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_769), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_820), .B(n_807), .Y(n_850) );
OAI21xp33_ASAP7_75t_L g851 ( .A1(n_754), .A2(n_768), .B(n_828), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_767), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_785), .A2(n_721), .B1(n_673), .B2(n_710), .Y(n_853) );
INVx1_ASAP7_75t_SL g854 ( .A(n_810), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_773), .B(n_740), .Y(n_855) );
OAI211xp5_ASAP7_75t_L g856 ( .A1(n_746), .A2(n_724), .B(n_658), .C(n_674), .Y(n_856) );
AND2x2_ASAP7_75t_L g857 ( .A(n_796), .B(n_739), .Y(n_857) );
NOR2x1_ASAP7_75t_L g858 ( .A(n_758), .B(n_741), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_767), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_790), .B(n_739), .Y(n_860) );
NAND2xp33_ASAP7_75t_SL g861 ( .A(n_819), .B(n_712), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_762), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_776), .Y(n_863) );
OR2x2_ASAP7_75t_L g864 ( .A(n_754), .B(n_698), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_783), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_784), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_779), .B(n_739), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_787), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_792), .Y(n_869) );
O2A1O1Ixp33_ASAP7_75t_L g870 ( .A1(n_768), .A2(n_608), .B(n_737), .C(n_735), .Y(n_870) );
OAI222xp33_ASAP7_75t_L g871 ( .A1(n_809), .A2(n_694), .B1(n_679), .B2(n_732), .C1(n_686), .C2(n_639), .Y(n_871) );
INVx1_ASAP7_75t_SL g872 ( .A(n_778), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_811), .B(n_686), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_818), .A2(n_686), .B1(n_664), .B2(n_694), .Y(n_874) );
OAI21xp33_ASAP7_75t_L g875 ( .A1(n_821), .A2(n_639), .B(n_713), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_813), .A2(n_639), .B1(n_741), .B2(n_736), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_762), .Y(n_877) );
OAI21xp33_ASAP7_75t_L g878 ( .A1(n_770), .A2(n_716), .B(n_713), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g879 ( .A1(n_833), .A2(n_795), .B1(n_798), .B2(n_797), .C(n_802), .Y(n_879) );
OAI211xp5_ASAP7_75t_L g880 ( .A1(n_830), .A2(n_789), .B(n_825), .C(n_794), .Y(n_880) );
NAND4xp25_ASAP7_75t_L g881 ( .A(n_838), .B(n_825), .C(n_741), .D(n_743), .Y(n_881) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_854), .B(n_757), .Y(n_882) );
AOI222xp33_ASAP7_75t_L g883 ( .A1(n_851), .A2(n_799), .B1(n_804), .B2(n_827), .C1(n_826), .C2(n_817), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_861), .A2(n_781), .B1(n_786), .B2(n_664), .Y(n_884) );
AOI221xp5_ASAP7_75t_L g885 ( .A1(n_861), .A2(n_748), .B1(n_750), .B2(n_751), .C(n_755), .Y(n_885) );
AOI322xp5_ASAP7_75t_L g886 ( .A1(n_853), .A2(n_756), .A3(n_771), .B1(n_803), .B2(n_812), .C1(n_824), .C2(n_805), .Y(n_886) );
AOI221xp5_ASAP7_75t_L g887 ( .A1(n_834), .A2(n_801), .B1(n_814), .B2(n_761), .C(n_772), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_853), .A2(n_788), .B1(n_723), .B2(n_734), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_874), .A2(n_722), .B1(n_716), .B2(n_806), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_836), .B(n_824), .Y(n_890) );
AOI221xp5_ASAP7_75t_L g891 ( .A1(n_834), .A2(n_823), .B1(n_806), .B2(n_805), .C(n_800), .Y(n_891) );
BUFx2_ASAP7_75t_L g892 ( .A(n_858), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_876), .A2(n_581), .B1(n_623), .B2(n_626), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_839), .B(n_823), .Y(n_894) );
OAI221xp5_ASAP7_75t_L g895 ( .A1(n_875), .A2(n_800), .B1(n_793), .B2(n_782), .C(n_780), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_842), .A2(n_793), .B1(n_782), .B2(n_780), .C(n_775), .Y(n_896) );
NOR2xp33_ASAP7_75t_L g897 ( .A(n_872), .B(n_729), .Y(n_897) );
AOI222xp33_ASAP7_75t_L g898 ( .A1(n_843), .A2(n_665), .B1(n_774), .B2(n_775), .C1(n_695), .C2(n_594), .Y(n_898) );
OAI221xp5_ASAP7_75t_L g899 ( .A1(n_838), .A2(n_774), .B1(n_707), .B2(n_702), .C(n_700), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_852), .A2(n_626), .B1(n_631), .B2(n_627), .Y(n_900) );
OAI221xp5_ASAP7_75t_SL g901 ( .A1(n_856), .A2(n_603), .B1(n_602), .B2(n_631), .C(n_627), .Y(n_901) );
OR2x2_ASAP7_75t_L g902 ( .A(n_864), .B(n_733), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_859), .A2(n_625), .B1(n_614), .B2(n_610), .Y(n_903) );
AOI31xp33_ASAP7_75t_L g904 ( .A1(n_856), .A2(n_602), .A3(n_625), .B(n_610), .Y(n_904) );
OAI31xp33_ASAP7_75t_SL g905 ( .A1(n_837), .A2(n_614), .A3(n_637), .B(n_621), .Y(n_905) );
A2O1A1Ixp33_ASAP7_75t_L g906 ( .A1(n_870), .A2(n_603), .B(n_637), .C(n_621), .Y(n_906) );
OAI221xp5_ASAP7_75t_L g907 ( .A1(n_880), .A2(n_832), .B1(n_878), .B2(n_835), .C(n_855), .Y(n_907) );
OAI211xp5_ASAP7_75t_L g908 ( .A1(n_881), .A2(n_870), .B(n_877), .C(n_862), .Y(n_908) );
NAND4xp75_ASAP7_75t_L g909 ( .A(n_897), .B(n_877), .C(n_873), .D(n_831), .Y(n_909) );
AOI21xp5_ASAP7_75t_L g910 ( .A1(n_904), .A2(n_871), .B(n_840), .Y(n_910) );
NOR3xp33_ASAP7_75t_L g911 ( .A(n_899), .B(n_871), .C(n_726), .Y(n_911) );
OAI22xp33_ASAP7_75t_L g912 ( .A1(n_884), .A2(n_847), .B1(n_841), .B2(n_844), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_895), .A2(n_849), .B1(n_848), .B2(n_846), .C(n_866), .Y(n_913) );
AOI221xp5_ASAP7_75t_L g914 ( .A1(n_879), .A2(n_869), .B1(n_868), .B2(n_865), .C(n_863), .Y(n_914) );
AOI211xp5_ASAP7_75t_L g915 ( .A1(n_901), .A2(n_857), .B(n_867), .C(n_847), .Y(n_915) );
NOR2xp67_ASAP7_75t_L g916 ( .A(n_889), .B(n_829), .Y(n_916) );
AOI21xp5_ASAP7_75t_L g917 ( .A1(n_901), .A2(n_885), .B(n_892), .Y(n_917) );
NAND3xp33_ASAP7_75t_L g918 ( .A(n_886), .B(n_845), .C(n_597), .Y(n_918) );
OAI211xp5_ASAP7_75t_SL g919 ( .A1(n_898), .A2(n_845), .B(n_731), .C(n_728), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_896), .B(n_850), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_891), .B(n_860), .Y(n_921) );
OAI21x1_ASAP7_75t_SL g922 ( .A1(n_910), .A2(n_888), .B(n_887), .Y(n_922) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_917), .A2(n_882), .B1(n_890), .B2(n_894), .C(n_906), .Y(n_923) );
NOR4xp25_ASAP7_75t_L g924 ( .A(n_908), .B(n_893), .C(n_902), .D(n_903), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_914), .B(n_883), .Y(n_925) );
AND4x1_ASAP7_75t_L g926 ( .A(n_915), .B(n_905), .C(n_900), .D(n_88), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_920), .B(n_733), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_913), .B(n_731), .Y(n_928) );
OAI21xp33_ASAP7_75t_L g929 ( .A1(n_919), .A2(n_636), .B(n_635), .Y(n_929) );
OR2x2_ASAP7_75t_L g930 ( .A(n_927), .B(n_921), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_924), .B(n_909), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_928), .Y(n_932) );
OA22x2_ASAP7_75t_L g933 ( .A1(n_922), .A2(n_907), .B1(n_912), .B2(n_911), .Y(n_933) );
INVx3_ASAP7_75t_L g934 ( .A(n_926), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g935 ( .A1(n_931), .A2(n_925), .B1(n_923), .B2(n_918), .C(n_929), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_930), .Y(n_936) );
NOR3xp33_ASAP7_75t_L g937 ( .A(n_934), .B(n_916), .C(n_636), .Y(n_937) );
XNOR2x1_ASAP7_75t_L g938 ( .A(n_936), .B(n_933), .Y(n_938) );
XNOR2x1_ASAP7_75t_L g939 ( .A(n_935), .B(n_934), .Y(n_939) );
INVx2_ASAP7_75t_L g940 ( .A(n_939), .Y(n_940) );
AOI21xp5_ASAP7_75t_L g941 ( .A1(n_938), .A2(n_932), .B(n_937), .Y(n_941) );
OR3x1_ASAP7_75t_L g942 ( .A(n_941), .B(n_932), .C(n_83), .Y(n_942) );
BUFx2_ASAP7_75t_L g943 ( .A(n_940), .Y(n_943) );
OAI22xp33_ASAP7_75t_L g944 ( .A1(n_943), .A2(n_635), .B1(n_634), .B2(n_568), .Y(n_944) );
AOI222xp33_ASAP7_75t_L g945 ( .A1(n_944), .A2(n_942), .B1(n_634), .B2(n_568), .C1(n_94), .C2(n_99), .Y(n_945) );
OAI221xp5_ASAP7_75t_SL g946 ( .A1(n_945), .A2(n_82), .B1(n_89), .B2(n_91), .C(n_100), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_946), .B(n_104), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g948 ( .A1(n_947), .A2(n_109), .B1(n_106), .B2(n_107), .Y(n_948) );
endmodule