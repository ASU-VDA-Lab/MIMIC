module fake_jpeg_1928_n_115 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_115);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_SL g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_3),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_12),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_15),
.B1(n_20),
.B2(n_18),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_27),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_21),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_39),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_29),
.B1(n_18),
.B2(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_53),
.B1(n_57),
.B2(n_38),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_30),
.B1(n_14),
.B2(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_14),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_31),
.B1(n_23),
.B2(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_39),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_65),
.B1(n_67),
.B2(n_50),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_69),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_38),
.B1(n_23),
.B2(n_42),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

XOR2x2_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_31),
.Y(n_70)
);

AO22x1_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_57),
.B1(n_34),
.B2(n_31),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_47),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_70),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_87),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_68),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.C(n_75),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_57),
.C(n_68),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_57),
.B(n_4),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_79),
.B(n_71),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_77),
.B(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_97),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.C(n_34),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_95),
.C(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_106),
.Y(n_109)
);

AOI321xp33_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_97),
.A3(n_84),
.B1(n_89),
.B2(n_8),
.C(n_9),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_3),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_105),
.B(n_101),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_107),
.Y(n_111)
);

OAI21x1_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_4),
.B(n_7),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_108),
.B(n_111),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_10),
.Y(n_115)
);


endmodule