module fake_jpeg_9194_n_234 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_0),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_1),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_34),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_31),
.B1(n_24),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_50),
.B1(n_60),
.B2(n_62),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_31),
.B1(n_24),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_57),
.B1(n_59),
.B2(n_30),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_31),
.B1(n_28),
.B2(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_64),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_24),
.B1(n_32),
.B2(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_21),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_30),
.B1(n_19),
.B2(n_27),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_21),
.B1(n_34),
.B2(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_73),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_83),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_72),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_18),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_40),
.B1(n_36),
.B2(n_44),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_75),
.B1(n_68),
.B2(n_67),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_17),
.B1(n_25),
.B2(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_78),
.Y(n_99)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_88),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_22),
.B(n_25),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_52),
.C(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_15),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_29),
.B(n_23),
.C(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_89),
.B1(n_54),
.B2(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_14),
.Y(n_89)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_103),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_1),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_93),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_100),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_52),
.C(n_44),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_65),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_83),
.B(n_70),
.Y(n_128)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_108),
.Y(n_132)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_109),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_13),
.C(n_3),
.Y(n_108)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_61),
.B1(n_49),
.B2(n_30),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_75),
.B1(n_74),
.B2(n_66),
.Y(n_122)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_66),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_82),
.B1(n_30),
.B2(n_27),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_29),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_101),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_115),
.B(n_92),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_131),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_67),
.B(n_74),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_119),
.B(n_128),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_74),
.B(n_77),
.C(n_68),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_88),
.B1(n_76),
.B2(n_74),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_134),
.B1(n_113),
.B2(n_103),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_130),
.B1(n_2),
.B2(n_3),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_89),
.Y(n_126)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_66),
.B1(n_49),
.B2(n_19),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_102),
.Y(n_139)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g133 ( 
.A(n_111),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_91),
.A2(n_27),
.B1(n_19),
.B2(n_63),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_136),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_18),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_94),
.B1(n_106),
.B2(n_93),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_129),
.A2(n_96),
.B1(n_95),
.B2(n_94),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_138),
.A2(n_143),
.B1(n_152),
.B2(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_100),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_148),
.B(n_149),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_96),
.B(n_98),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_97),
.B(n_23),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_97),
.B(n_27),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_155),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_102),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_156),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_2),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_114),
.B(n_122),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_119),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_167),
.B1(n_146),
.B2(n_119),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_124),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_170),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_119),
.B1(n_124),
.B2(n_127),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_143),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_144),
.B(n_150),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_175),
.B(n_176),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_124),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_147),
.C(n_133),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_145),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_179),
.Y(n_195)
);

OAI322xp33_ASAP7_75t_L g179 ( 
.A1(n_163),
.A2(n_151),
.A3(n_146),
.B1(n_138),
.B2(n_149),
.C1(n_145),
.C2(n_137),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_187),
.C(n_189),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_186),
.B1(n_166),
.B2(n_160),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g185 ( 
.A(n_164),
.B(n_119),
.CI(n_127),
.CON(n_185),
.SN(n_185)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_168),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_147),
.B1(n_156),
.B2(n_134),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_2),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_3),
.C(n_5),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_192),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_6),
.C(n_7),
.Y(n_192)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_194),
.B(n_198),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_183),
.B1(n_185),
.B2(n_188),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_166),
.B1(n_160),
.B2(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_200),
.B1(n_180),
.B2(n_189),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_161),
.B(n_162),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_178),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_169),
.B(n_174),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_173),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_192),
.C(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_206),
.B(n_196),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_208),
.C(n_210),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_173),
.C(n_7),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_6),
.C(n_7),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_212),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_6),
.C(n_8),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_216),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_204),
.A2(n_199),
.B(n_193),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_212),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_217),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_195),
.B(n_202),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_9),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_195),
.C(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_213),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_217),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_221),
.A2(n_214),
.B1(n_9),
.B2(n_12),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_12),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_228),
.C(n_221),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_227),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_12),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_223),
.C(n_220),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_228),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_229),
.Y(n_234)
);


endmodule