module fake_jpeg_13721_n_171 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_15),
.B(n_47),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_49),
.C(n_48),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_0),
.Y(n_79)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_52),
.Y(n_80)
);

AO22x1_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_71),
.B1(n_67),
.B2(n_69),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_61),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_43),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_70),
.B1(n_65),
.B2(n_73),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_94),
.B1(n_99),
.B2(n_72),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_70),
.B(n_65),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_78),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2x1_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_71),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_57),
.B(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_1),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_59),
.B1(n_68),
.B2(n_54),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_28),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_75),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_53),
.B1(n_54),
.B2(n_60),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_109),
.B(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_62),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_64),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_19),
.C(n_40),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_50),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_110),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_53),
.B1(n_75),
.B2(n_67),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_112),
.B1(n_5),
.B2(n_6),
.Y(n_123)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_115),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_58),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_56),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_2),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_118),
.B(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_4),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_120),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_102),
.C(n_100),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_131),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_152)
);

XNOR2x1_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_42),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_104),
.B(n_119),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_128),
.B(n_136),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_116),
.B(n_103),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_21),
.C(n_35),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_135),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_8),
.B(n_9),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_10),
.B(n_11),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_12),
.Y(n_144)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_138),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_154),
.C(n_155),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_12),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_150),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_129),
.A2(n_26),
.B1(n_33),
.B2(n_32),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_29),
.B(n_30),
.Y(n_161)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_152),
.B1(n_144),
.B2(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_18),
.Y(n_153)
);

NOR4xp25_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_131),
.C(n_137),
.D(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_24),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_161),
.B1(n_145),
.B2(n_149),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_146),
.C(n_124),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_164),
.C(n_158),
.Y(n_165)
);

AO221x1_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_136),
.B1(n_127),
.B2(n_145),
.C(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_147),
.Y(n_168)
);

NOR4xp25_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_160),
.C(n_166),
.D(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_146),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_154),
.Y(n_171)
);


endmodule