module fake_jpeg_11877_n_421 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_421);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_421;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_44),
.B(n_45),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_49),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_0),
.Y(n_48)
);

NAND2x1_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_89),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_51),
.B(n_87),
.Y(n_115)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_60),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_59),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_12),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_19),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_65),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_12),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_28),
.Y(n_69)
);

NAND2x1_ASAP7_75t_SL g141 ( 
.A(n_69),
.B(n_83),
.Y(n_141)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_28),
.B(n_7),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_78),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_32),
.B(n_7),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_81),
.Y(n_143)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_91),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_29),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_93),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g94 ( 
.A(n_31),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_37),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_37),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_48),
.A2(n_18),
.B1(n_39),
.B2(n_21),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_100),
.B(n_148),
.C(n_0),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_40),
.B1(n_33),
.B2(n_18),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_105),
.A2(n_119),
.B1(n_120),
.B2(n_75),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_39),
.B1(n_21),
.B2(n_31),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_131),
.B1(n_144),
.B2(n_145),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_39),
.B1(n_21),
.B2(n_14),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_14),
.B1(n_24),
.B2(n_37),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_89),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_80),
.A2(n_37),
.B1(n_31),
.B2(n_34),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_69),
.B(n_33),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_24),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_84),
.A2(n_37),
.B1(n_31),
.B2(n_34),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_55),
.A2(n_27),
.B1(n_23),
.B2(n_8),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_48),
.A2(n_27),
.B1(n_23),
.B2(n_2),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_150),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_SL g193 ( 
.A(n_151),
.B(n_160),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_67),
.B1(n_59),
.B2(n_63),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_158),
.B1(n_162),
.B2(n_176),
.Y(n_192)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_101),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_71),
.B1(n_57),
.B2(n_74),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g209 ( 
.A1(n_159),
.A2(n_123),
.B1(n_127),
.B2(n_124),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_89),
.B(n_85),
.C(n_73),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_107),
.B(n_52),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_171),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_106),
.A2(n_68),
.B1(n_77),
.B2(n_50),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_94),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_98),
.B(n_94),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_110),
.B(n_70),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_177),
.Y(n_202)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

BUFx4f_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_100),
.A2(n_83),
.B1(n_54),
.B2(n_46),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_122),
.B1(n_109),
.B2(n_113),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_126),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_178),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_112),
.A2(n_56),
.B1(n_95),
.B2(n_72),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_104),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_117),
.B(n_53),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_180),
.Y(n_217)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_181),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_182),
.A2(n_141),
.B1(n_133),
.B2(n_137),
.Y(n_208)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_183),
.Y(n_205)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_141),
.A2(n_93),
.B1(n_81),
.B2(n_8),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_97),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_139),
.A2(n_43),
.B1(n_7),
.B2(n_9),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_191),
.A2(n_145),
.B1(n_122),
.B2(n_109),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_140),
.C(n_147),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_195),
.B(n_211),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_149),
.B1(n_113),
.B2(n_129),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_200),
.A2(n_201),
.B1(n_220),
.B2(n_191),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_108),
.B1(n_131),
.B2(n_144),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_209),
.B1(n_173),
.B2(n_149),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_161),
.B(n_103),
.CI(n_148),
.CON(n_207),
.SN(n_207)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_207),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_137),
.B(n_187),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_118),
.Y(n_211)
);

NAND2xp33_ASAP7_75t_SL g213 ( 
.A(n_160),
.B(n_167),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_133),
.B(n_143),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_151),
.B1(n_154),
.B2(n_134),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_151),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_229),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_225),
.A2(n_209),
.B1(n_215),
.B2(n_198),
.Y(n_264)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_171),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_230),
.A2(n_234),
.B1(n_245),
.B2(n_205),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_218),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_239),
.Y(n_269)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_157),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_152),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_236),
.B(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_132),
.B1(n_124),
.B2(n_121),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_238),
.A2(n_201),
.B1(n_209),
.B2(n_192),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_185),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_242),
.B(n_219),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_208),
.B(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_155),
.Y(n_244)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_132),
.B1(n_116),
.B2(n_127),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_180),
.Y(n_246)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_163),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_248),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_213),
.B(n_193),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_250),
.A2(n_251),
.B(n_254),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_193),
.B(n_219),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_258),
.A2(n_259),
.B1(n_264),
.B2(n_266),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_225),
.A2(n_207),
.B1(n_209),
.B2(n_192),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_242),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_263),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_223),
.B1(n_245),
.B2(n_234),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_184),
.B1(n_198),
.B2(n_190),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_265),
.Y(n_273)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_235),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_275),
.C(n_281),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_235),
.C(n_246),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_277),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_269),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_228),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_282),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_246),
.C(n_237),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_237),
.C(n_244),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_230),
.B1(n_245),
.B2(n_239),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_284),
.A2(n_292),
.B1(n_263),
.B2(n_251),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_224),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_286),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_224),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_233),
.C(n_229),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_289),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_SL g288 ( 
.A1(n_250),
.A2(n_240),
.B(n_229),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_295),
.B(n_257),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_233),
.C(n_248),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_258),
.A2(n_232),
.B1(n_227),
.B2(n_238),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_231),
.C(n_236),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_294),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_238),
.C(n_247),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_241),
.C(n_214),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_261),
.Y(n_301)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_305),
.Y(n_318)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_313),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_282),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_317),
.B1(n_252),
.B2(n_271),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_291),
.A2(n_256),
.B1(n_253),
.B2(n_252),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_312),
.A2(n_301),
.B1(n_299),
.B2(n_296),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_279),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_285),
.A2(n_256),
.B(n_253),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_249),
.Y(n_326)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_275),
.C(n_274),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_324),
.C(n_330),
.Y(n_344)
);

FAx1_ASAP7_75t_SL g320 ( 
.A(n_316),
.B(n_287),
.CI(n_281),
.CON(n_320),
.SN(n_320)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_320),
.B(n_297),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_323),
.A2(n_188),
.B1(n_221),
.B2(n_186),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_271),
.C(n_197),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_306),
.A2(n_249),
.B1(n_226),
.B2(n_194),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_325),
.A2(n_328),
.B1(n_329),
.B2(n_335),
.Y(n_343)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_326),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_301),
.A2(n_315),
.B1(n_305),
.B2(n_313),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_197),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_SL g331 ( 
.A(n_314),
.B(n_150),
.C(n_221),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_331),
.A2(n_334),
.B(n_316),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_317),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_332),
.B(n_310),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_308),
.A2(n_312),
.B(n_303),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_311),
.A2(n_226),
.B1(n_214),
.B2(n_183),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_307),
.C(n_309),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_316),
.C(n_297),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_333),
.A2(n_304),
.B1(n_298),
.B2(n_296),
.Y(n_341)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_341),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_346),
.B(n_327),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_354),
.Y(n_362)
);

NOR2x1_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_179),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_206),
.C(n_128),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_353),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_335),
.A2(n_150),
.B1(n_168),
.B2(n_221),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_350),
.A2(n_327),
.B1(n_339),
.B2(n_334),
.Y(n_361)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_337),
.Y(n_351)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_351),
.Y(n_371)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_352),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_206),
.C(n_102),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_L g354 ( 
.A1(n_318),
.A2(n_221),
.B(n_150),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_356),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_328),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_325),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_357),
.B(n_320),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_364),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_361),
.A2(n_365),
.B1(n_340),
.B2(n_357),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_346),
.C(n_336),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_363),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_330),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_343),
.A2(n_338),
.B1(n_320),
.B2(n_322),
.Y(n_365)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_366),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_353),
.B(n_342),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_367),
.A2(n_137),
.B(n_179),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_331),
.C(n_102),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_368),
.B(n_351),
.Y(n_378)
);

AOI21x1_ASAP7_75t_L g375 ( 
.A1(n_370),
.A2(n_352),
.B(n_348),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_347),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_381),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_375),
.A2(n_385),
.B1(n_373),
.B2(n_359),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_370),
.A2(n_356),
.B(n_340),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_382),
.B(n_383),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_372),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_379),
.B(n_386),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_343),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_365),
.A2(n_355),
.B(n_349),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_360),
.A2(n_169),
.B(n_166),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_384),
.B(n_368),
.Y(n_392)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_371),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_181),
.Y(n_386)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_389),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_391),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_393),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_380),
.A2(n_377),
.B1(n_374),
.B2(n_382),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_381),
.C(n_376),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_394),
.A2(n_396),
.B(n_123),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_364),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_395),
.B(n_398),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_386),
.B(n_369),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_380),
.B(n_362),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_369),
.Y(n_402)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_402),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_403),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_5),
.C(n_10),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_404),
.B(n_406),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_390),
.C(n_397),
.Y(n_407)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_407),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_390),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_409),
.A2(n_412),
.B(n_9),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_5),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_402),
.C(n_400),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_413),
.B(n_414),
.C(n_416),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_7),
.Y(n_414)
);

AOI321xp33_ASAP7_75t_L g417 ( 
.A1(n_415),
.A2(n_408),
.A3(n_411),
.B1(n_10),
.B2(n_11),
.C(n_2),
.Y(n_417)
);

AO21x1_ASAP7_75t_L g419 ( 
.A1(n_417),
.A2(n_414),
.B(n_1),
.Y(n_419)
);

AO221x1_ASAP7_75t_L g420 ( 
.A1(n_419),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.C(n_418),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_1),
.Y(n_421)
);


endmodule