module fake_jpeg_1393_n_74 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_32),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_39),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_23),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_29),
.B1(n_23),
.B2(n_21),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_0),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_31),
.C(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_47),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_49),
.B1(n_52),
.B2(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_4),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_41),
.B1(n_2),
.B2(n_3),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_1),
.B(n_4),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_61),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_60),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_15),
.C(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_66),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_59),
.C(n_56),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_69),
.B(n_63),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_68),
.C(n_62),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_65),
.C(n_7),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_5),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_63),
.C2(n_60),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_10),
.Y(n_74)
);


endmodule