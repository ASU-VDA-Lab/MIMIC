module fake_netlist_6_2671_n_773 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_773);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_773;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_148;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_153;
wire n_758;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_515;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_8),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_76),
.Y(n_148)
);

BUFx2_ASAP7_75t_SL g149 ( 
.A(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_1),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_31),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_34),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_48),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_41),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_140),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_49),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_105),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_38),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_4),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_71),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_47),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_93),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_81),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_68),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_39),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_18),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_138),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_91),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_62),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_51),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_86),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_12),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_0),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_4),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_19),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_60),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_14),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_102),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_61),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_40),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_25),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_32),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_0),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_172),
.B(n_1),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_2),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_153),
.B(n_2),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_150),
.B(n_3),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_165),
.B(n_173),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_3),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

AND2x6_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_145),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_5),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_5),
.Y(n_228)
);

AND2x4_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_144),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_151),
.B(n_6),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_154),
.B(n_26),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_155),
.B(n_141),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_157),
.B(n_158),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_221),
.B1(n_207),
.B2(n_216),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_152),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_152),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_L g243 ( 
.A1(n_231),
.A2(n_184),
.B1(n_156),
.B2(n_181),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_231),
.B1(n_212),
.B2(n_214),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

OR2x6_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_230),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_220),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_148),
.B1(n_156),
.B2(n_181),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_205),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_184),
.B1(n_148),
.B2(n_183),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_220),
.Y(n_252)
);

AO22x2_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_149),
.B1(n_7),
.B2(n_9),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_183),
.B1(n_192),
.B2(n_190),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_203),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_169),
.B1(n_177),
.B2(n_175),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g257 ( 
.A1(n_230),
.A2(n_182),
.B1(n_170),
.B2(n_168),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_160),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_R g259 ( 
.A1(n_202),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_163),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_167),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_215),
.Y(n_262)
);

NAND3x1_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_10),
.C(n_11),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_226),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_230),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_230),
.B(n_13),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_235),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_230),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g273 ( 
.A1(n_232),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_235),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_232),
.A2(n_234),
.B1(n_205),
.B2(n_210),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_232),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_204),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_L g278 ( 
.A1(n_232),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_206),
.B(n_20),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_235),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_233),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_204),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_205),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_232),
.B(n_29),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_232),
.A2(n_234),
.B1(n_210),
.B2(n_211),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_276),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_234),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_249),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_252),
.B(n_242),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_247),
.B(n_205),
.Y(n_296)
);

BUFx6f_ASAP7_75t_SL g297 ( 
.A(n_247),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_200),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

INVxp33_ASAP7_75t_SL g300 ( 
.A(n_239),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_205),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_244),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_200),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_258),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_254),
.B(n_234),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_200),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_277),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_261),
.B(n_229),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_275),
.A2(n_229),
.B(n_238),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_205),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_275),
.A2(n_229),
.B(n_224),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_206),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_257),
.B(n_200),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_254),
.B(n_234),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_206),
.Y(n_325)
);

NAND2x1p5_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_235),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_253),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_253),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_253),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_209),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_250),
.B(n_236),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_243),
.B(n_234),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_243),
.B(n_210),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_267),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_263),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_285),
.B(n_236),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_281),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_267),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_251),
.B(n_210),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_273),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_273),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_278),
.Y(n_345)
);

OR2x6_ASAP7_75t_L g346 ( 
.A(n_259),
.B(n_236),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_278),
.B(n_236),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_276),
.B(n_200),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_210),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_316),
.B(n_317),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_292),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_294),
.B(n_210),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_314),
.Y(n_355)
);

AND2x2_ASAP7_75t_SL g356 ( 
.A(n_307),
.B(n_217),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_320),
.A2(n_224),
.B(n_225),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_286),
.B(n_200),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_288),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_316),
.B(n_219),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_312),
.B(n_219),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_312),
.B(n_219),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_201),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_289),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_201),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_321),
.Y(n_370)
);

BUFx4f_ASAP7_75t_L g371 ( 
.A(n_319),
.Y(n_371)
);

AND2x2_ASAP7_75t_SL g372 ( 
.A(n_307),
.B(n_225),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_201),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_290),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_301),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_305),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_308),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_309),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_324),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_321),
.B(n_224),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_313),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_324),
.B(n_211),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_287),
.B(n_201),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_287),
.B(n_201),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_312),
.B(n_209),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_331),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_331),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_336),
.B(n_209),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_315),
.B(n_201),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_325),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_306),
.B(n_227),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_328),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_306),
.B(n_211),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_325),
.B(n_224),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_342),
.B(n_215),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_311),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_339),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_297),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_347),
.A2(n_224),
.B(n_215),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_333),
.B(n_224),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_339),
.B(n_211),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_318),
.B(n_211),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_329),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_335),
.B(n_202),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_334),
.B(n_211),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_300),
.B(n_204),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_326),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_347),
.A2(n_224),
.B(n_222),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_348),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_338),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_364),
.Y(n_417)
);

OR2x6_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_326),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_332),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_349),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_330),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_346),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_337),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_332),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_381),
.B(n_300),
.Y(n_426)
);

BUFx12f_ASAP7_75t_L g427 ( 
.A(n_403),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_356),
.B(n_341),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_349),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_371),
.B(n_343),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_349),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_364),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_351),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_351),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_351),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_360),
.B(n_346),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_356),
.B(n_344),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_346),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_377),
.B(n_296),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_377),
.B(n_302),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_356),
.B(n_297),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_394),
.B(n_346),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_377),
.B(n_345),
.Y(n_444)
);

BUFx12f_ASAP7_75t_L g445 ( 
.A(n_364),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_293),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_387),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_372),
.B(n_297),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_375),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_372),
.B(n_322),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_375),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_392),
.B(n_303),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_395),
.Y(n_454)
);

OR2x6_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_223),
.Y(n_455)
);

BUFx4f_ASAP7_75t_L g456 ( 
.A(n_392),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

AND2x6_ASAP7_75t_L g458 ( 
.A(n_382),
.B(n_304),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_380),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_352),
.B(n_303),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_372),
.B(n_204),
.Y(n_461)
);

NAND2x1_ASAP7_75t_L g462 ( 
.A(n_364),
.B(n_298),
.Y(n_462)
);

OR2x6_ASAP7_75t_L g463 ( 
.A(n_412),
.B(n_223),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_380),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_363),
.B(n_204),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_388),
.B(n_310),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_352),
.B(n_30),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_388),
.B(n_222),
.Y(n_468)
);

AND2x2_ASAP7_75t_SL g469 ( 
.A(n_412),
.B(n_204),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_389),
.B(n_222),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_392),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_454),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_452),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_427),
.Y(n_476)
);

BUFx8_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_428),
.B(n_409),
.Y(n_478)
);

INVx8_ASAP7_75t_L g479 ( 
.A(n_418),
.Y(n_479)
);

BUFx5_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_417),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_437),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_420),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_439),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_428),
.A2(n_389),
.B1(n_357),
.B2(n_392),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_416),
.Y(n_486)
);

BUFx4_ASAP7_75t_SL g487 ( 
.A(n_443),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_416),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_444),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_444),
.Y(n_490)
);

BUFx2_ASAP7_75t_R g491 ( 
.A(n_446),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_426),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_417),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_426),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_442),
.Y(n_495)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_456),
.B(n_371),
.Y(n_496)
);

BUFx2_ASAP7_75t_SL g497 ( 
.A(n_452),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_459),
.Y(n_498)
);

BUFx12f_ASAP7_75t_L g499 ( 
.A(n_467),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

INVx3_ASAP7_75t_SL g501 ( 
.A(n_419),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_417),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_438),
.B(n_392),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_467),
.Y(n_504)
);

BUFx2_ASAP7_75t_SL g505 ( 
.A(n_459),
.Y(n_505)
);

INVx6_ASAP7_75t_SL g506 ( 
.A(n_455),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_449),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_424),
.B(n_409),
.Y(n_509)
);

CKINVDCx8_ASAP7_75t_R g510 ( 
.A(n_419),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_425),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_425),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_453),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_453),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_455),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_451),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_424),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_474),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_478),
.B(n_438),
.Y(n_520)
);

BUFx8_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_494),
.A2(n_442),
.B1(n_448),
.B2(n_461),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_473),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_483),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_514),
.A2(n_392),
.B1(n_448),
.B2(n_340),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_515),
.A2(n_512),
.B1(n_511),
.B2(n_478),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_508),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_507),
.Y(n_529)
);

CKINVDCx6p67_ASAP7_75t_R g530 ( 
.A(n_476),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_481),
.Y(n_531)
);

BUFx8_ASAP7_75t_L g532 ( 
.A(n_472),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_502),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_489),
.A2(n_340),
.B1(n_450),
.B2(n_423),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_494),
.A2(n_461),
.B1(n_357),
.B2(n_469),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_498),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_499),
.A2(n_450),
.B1(n_447),
.B2(n_441),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_499),
.A2(n_501),
.B1(n_504),
.B2(n_486),
.Y(n_538)
);

INVx6_ASAP7_75t_L g539 ( 
.A(n_477),
.Y(n_539)
);

INVx6_ASAP7_75t_L g540 ( 
.A(n_477),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_501),
.A2(n_441),
.B1(n_440),
.B2(n_430),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_SL g542 ( 
.A1(n_492),
.A2(n_495),
.B1(n_518),
.B2(n_477),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_498),
.Y(n_543)
);

INVx8_ASAP7_75t_L g544 ( 
.A(n_479),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_481),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_509),
.A2(n_371),
.B1(n_418),
.B2(n_469),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_479),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_517),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_503),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_485),
.A2(n_371),
.B1(n_418),
.B2(n_421),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_488),
.B(n_363),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_503),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_SL g553 ( 
.A1(n_492),
.A2(n_456),
.B1(n_404),
.B2(n_413),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_486),
.A2(n_440),
.B1(n_430),
.B2(n_399),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_490),
.A2(n_399),
.B1(n_365),
.B2(n_366),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_510),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_502),
.Y(n_557)
);

NAND2x1p5_ASAP7_75t_L g558 ( 
.A(n_502),
.B(n_435),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_481),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_481),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_485),
.B(n_421),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_475),
.B(n_395),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_535),
.A2(n_482),
.B1(n_484),
.B2(n_490),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_523),
.A2(n_516),
.B1(n_350),
.B2(n_354),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_552),
.B(n_390),
.Y(n_565)
);

NOR2x1_ASAP7_75t_L g566 ( 
.A(n_561),
.B(n_500),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_526),
.A2(n_510),
.B1(n_491),
.B2(n_455),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_522),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_549),
.B(n_390),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_539),
.A2(n_479),
.B1(n_404),
.B2(n_413),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_534),
.A2(n_365),
.B1(n_366),
.B2(n_410),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_521),
.Y(n_572)
);

OAI222xp33_ASAP7_75t_L g573 ( 
.A1(n_553),
.A2(n_463),
.B1(n_358),
.B2(n_496),
.C1(n_471),
.C2(n_466),
.Y(n_573)
);

OAI222xp33_ASAP7_75t_L g574 ( 
.A1(n_527),
.A2(n_463),
.B1(n_358),
.B2(n_496),
.C1(n_466),
.C2(n_384),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_520),
.B(n_395),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_525),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_SL g577 ( 
.A1(n_539),
.A2(n_479),
.B1(n_391),
.B2(n_505),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_L g578 ( 
.A1(n_556),
.A2(n_463),
.B1(n_506),
.B2(n_374),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_519),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_529),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_521),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_520),
.B(n_396),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_524),
.A2(n_374),
.B1(n_368),
.B2(n_362),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_396),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_542),
.A2(n_397),
.B(n_382),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_548),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_528),
.B(n_396),
.Y(n_587)
);

AND2x2_ASAP7_75t_SL g588 ( 
.A(n_561),
.B(n_432),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_537),
.A2(n_497),
.B1(n_506),
.B2(n_475),
.Y(n_589)
);

AOI222xp33_ASAP7_75t_L g590 ( 
.A1(n_555),
.A2(n_368),
.B1(n_362),
.B2(n_408),
.C1(n_355),
.C2(n_470),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_538),
.A2(n_398),
.B(n_382),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_536),
.B(n_472),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_SL g594 ( 
.A1(n_540),
.A2(n_480),
.B1(n_458),
.B2(n_500),
.Y(n_594)
);

BUFx4f_ASAP7_75t_SL g595 ( 
.A(n_530),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_554),
.A2(n_546),
.B1(n_550),
.B2(n_540),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_562),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_558),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_536),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_546),
.A2(n_506),
.B1(n_458),
.B2(n_383),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_541),
.A2(n_398),
.B(n_382),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_550),
.A2(n_398),
.B(n_405),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_532),
.A2(n_480),
.B1(n_458),
.B2(n_500),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_536),
.Y(n_604)
);

BUFx12f_ASAP7_75t_L g605 ( 
.A(n_532),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_547),
.A2(n_458),
.B1(n_383),
.B2(n_355),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_543),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_547),
.A2(n_465),
.B1(n_414),
.B2(n_480),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_544),
.A2(n_480),
.B1(n_468),
.B2(n_470),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_531),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_596),
.A2(n_480),
.B1(n_544),
.B2(n_543),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_L g612 ( 
.A1(n_567),
.A2(n_544),
.B1(n_543),
.B2(n_468),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_564),
.A2(n_480),
.B1(n_407),
.B2(n_376),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_563),
.A2(n_480),
.B1(n_379),
.B2(n_376),
.Y(n_614)
);

OAI221xp5_ASAP7_75t_L g615 ( 
.A1(n_585),
.A2(n_408),
.B1(n_462),
.B2(n_406),
.C(n_487),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_588),
.A2(n_375),
.B1(n_379),
.B2(n_376),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_588),
.A2(n_379),
.B1(n_361),
.B2(n_378),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_SL g618 ( 
.A1(n_589),
.A2(n_531),
.B1(n_533),
.B2(n_557),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_578),
.A2(n_378),
.B1(n_353),
.B2(n_361),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_583),
.A2(n_531),
.B1(n_558),
.B2(n_533),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_600),
.A2(n_353),
.B1(n_361),
.B2(n_378),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_571),
.A2(n_353),
.B1(n_361),
.B2(n_378),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_565),
.A2(n_353),
.B1(n_398),
.B2(n_401),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_565),
.A2(n_401),
.B1(n_222),
.B2(n_559),
.Y(n_624)
);

OAI221xp5_ASAP7_75t_L g625 ( 
.A1(n_591),
.A2(n_373),
.B1(n_401),
.B2(n_557),
.C(n_493),
.Y(n_625)
);

OAI222xp33_ASAP7_75t_L g626 ( 
.A1(n_570),
.A2(n_431),
.B1(n_436),
.B2(n_434),
.C1(n_433),
.C2(n_429),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_SL g627 ( 
.A1(n_569),
.A2(n_432),
.B(n_457),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_586),
.B(n_575),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_590),
.A2(n_559),
.B1(n_405),
.B2(n_457),
.Y(n_629)
);

OAI221xp5_ASAP7_75t_L g630 ( 
.A1(n_601),
.A2(n_493),
.B1(n_457),
.B2(n_213),
.C(n_367),
.Y(n_630)
);

OAI22x1_ASAP7_75t_L g631 ( 
.A1(n_566),
.A2(n_493),
.B1(n_502),
.B2(n_545),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_577),
.A2(n_502),
.B1(n_559),
.B2(n_513),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_605),
.A2(n_405),
.B1(n_213),
.B2(n_513),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_605),
.A2(n_405),
.B1(n_213),
.B2(n_513),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_602),
.A2(n_213),
.B1(n_359),
.B2(n_369),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_SL g636 ( 
.A1(n_607),
.A2(n_513),
.B1(n_545),
.B2(n_560),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_609),
.A2(n_213),
.B1(n_560),
.B2(n_385),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_608),
.A2(n_213),
.B1(n_386),
.B2(n_36),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_L g639 ( 
.A(n_566),
.B(n_33),
.C(n_35),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_586),
.A2(n_594),
.B1(n_606),
.B2(n_579),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_579),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_603),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_575),
.B(n_50),
.Y(n_643)
);

NOR2xp67_ASAP7_75t_L g644 ( 
.A(n_576),
.B(n_52),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_SL g645 ( 
.A1(n_607),
.A2(n_572),
.B1(n_595),
.B2(n_581),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_604),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_646)
);

OAI21xp33_ASAP7_75t_L g647 ( 
.A1(n_584),
.A2(n_56),
.B(n_57),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_628),
.B(n_580),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_643),
.B(n_580),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_640),
.B(n_593),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_635),
.B(n_568),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_635),
.B(n_568),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_611),
.B(n_576),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_612),
.B(n_598),
.Y(n_654)
);

NAND4xp25_ASAP7_75t_SL g655 ( 
.A(n_645),
.B(n_572),
.C(n_610),
.D(n_587),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_644),
.B(n_593),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_615),
.A2(n_581),
.B1(n_592),
.B2(n_599),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_644),
.B(n_597),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_614),
.A2(n_599),
.B1(n_610),
.B2(n_582),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_613),
.B(n_597),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_SL g661 ( 
.A1(n_630),
.A2(n_598),
.B(n_573),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_618),
.B(n_58),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_647),
.B(n_574),
.C(n_63),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_616),
.B(n_59),
.Y(n_664)
);

OAI221xp5_ASAP7_75t_SL g665 ( 
.A1(n_642),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.C(n_67),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_636),
.B(n_625),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_631),
.B(n_69),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_623),
.B(n_70),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_631),
.B(n_72),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_617),
.B(n_73),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_637),
.B(n_74),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_629),
.B(n_75),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_641),
.B(n_78),
.C(n_79),
.Y(n_673)
);

OAI21xp33_ASAP7_75t_L g674 ( 
.A1(n_646),
.A2(n_80),
.B(n_82),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_632),
.B(n_83),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_627),
.B(n_84),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_648),
.B(n_639),
.Y(n_677)
);

NOR3xp33_ASAP7_75t_L g678 ( 
.A(n_657),
.B(n_620),
.C(n_626),
.Y(n_678)
);

NOR2x1_ASAP7_75t_SL g679 ( 
.A(n_656),
.B(n_627),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_L g680 ( 
.A(n_666),
.B(n_638),
.C(n_634),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_653),
.Y(n_681)
);

OAI221xp5_ASAP7_75t_SL g682 ( 
.A1(n_674),
.A2(n_633),
.B1(n_619),
.B2(n_624),
.C(n_622),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_649),
.B(n_621),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_651),
.B(n_85),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_651),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_658),
.B(n_87),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_653),
.B(n_88),
.Y(n_687)
);

AOI211x1_ASAP7_75t_L g688 ( 
.A1(n_655),
.A2(n_89),
.B(n_90),
.C(n_92),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_650),
.B(n_94),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_652),
.B(n_95),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_652),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_660),
.B(n_96),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_660),
.B(n_667),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_693),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_693),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_685),
.Y(n_696)
);

XNOR2xp5_ASAP7_75t_L g697 ( 
.A(n_688),
.B(n_662),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_685),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_686),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_691),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_691),
.B(n_667),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_681),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_679),
.Y(n_703)
);

XNOR2x2_ASAP7_75t_L g704 ( 
.A(n_680),
.B(n_663),
.Y(n_704)
);

XOR2x2_ASAP7_75t_L g705 ( 
.A(n_697),
.B(n_689),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_702),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_696),
.Y(n_707)
);

XNOR2xp5_ASAP7_75t_L g708 ( 
.A(n_697),
.B(n_692),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_698),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_706),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_705),
.A2(n_703),
.B1(n_678),
.B2(n_699),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_707),
.Y(n_712)
);

AO22x2_ASAP7_75t_L g713 ( 
.A1(n_707),
.A2(n_695),
.B1(n_696),
.B2(n_701),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_709),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_714),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_710),
.Y(n_716)
);

OA22x2_ASAP7_75t_L g717 ( 
.A1(n_711),
.A2(n_708),
.B1(n_705),
.B2(n_701),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_712),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_715),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_717),
.A2(n_708),
.B1(n_694),
.B2(n_699),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_SL g721 ( 
.A1(n_716),
.A2(n_704),
.B1(n_699),
.B2(n_713),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_721),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_720),
.A2(n_718),
.B1(n_713),
.B2(n_694),
.Y(n_723)
);

OAI22x1_ASAP7_75t_L g724 ( 
.A1(n_719),
.A2(n_704),
.B1(n_689),
.B2(n_701),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_720),
.A2(n_699),
.B1(n_692),
.B2(n_687),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_724),
.B(n_699),
.Y(n_726)
);

AO22x2_ASAP7_75t_L g727 ( 
.A1(n_722),
.A2(n_686),
.B1(n_663),
.B2(n_690),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_725),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_723),
.A2(n_662),
.B1(n_677),
.B2(n_669),
.Y(n_729)
);

AOI221xp5_ASAP7_75t_L g730 ( 
.A1(n_722),
.A2(n_661),
.B1(n_665),
.B2(n_684),
.C(n_674),
.Y(n_730)
);

NOR4xp25_ASAP7_75t_L g731 ( 
.A(n_722),
.B(n_669),
.C(n_675),
.D(n_676),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_722),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_732),
.B(n_700),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_728),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_726),
.B(n_700),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_727),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_729),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_731),
.B(n_683),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_730),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_736),
.Y(n_740)
);

NAND4xp25_ASAP7_75t_L g741 ( 
.A(n_734),
.B(n_676),
.C(n_673),
.D(n_682),
.Y(n_741)
);

AO22x2_ASAP7_75t_L g742 ( 
.A1(n_737),
.A2(n_671),
.B1(n_664),
.B2(n_654),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_738),
.A2(n_671),
.B1(n_670),
.B2(n_664),
.Y(n_743)
);

NOR3xp33_ASAP7_75t_L g744 ( 
.A(n_739),
.B(n_733),
.C(n_735),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_735),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_735),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_734),
.A2(n_670),
.B1(n_659),
.B2(n_672),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_734),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_745),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_740),
.B(n_661),
.Y(n_750)
);

INVxp33_ASAP7_75t_SL g751 ( 
.A(n_744),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_746),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_743),
.A2(n_668),
.B1(n_100),
.B2(n_101),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_748),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_742),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_747),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_751),
.A2(n_754),
.B1(n_750),
.B2(n_752),
.Y(n_757)
);

OAI22x1_ASAP7_75t_L g758 ( 
.A1(n_755),
.A2(n_741),
.B1(n_104),
.B2(n_106),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_756),
.A2(n_99),
.B1(n_108),
.B2(n_109),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_749),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_SL g761 ( 
.A1(n_749),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_753),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_760),
.B(n_114),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_757),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_758),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_L g766 ( 
.A1(n_765),
.A2(n_762),
.B1(n_759),
.B2(n_761),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_764),
.A2(n_115),
.B1(n_117),
.B2(n_119),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_763),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_766),
.Y(n_769)
);

OAI22xp33_ASAP7_75t_L g770 ( 
.A1(n_769),
.A2(n_768),
.B1(n_767),
.B2(n_126),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_770),
.B(n_124),
.Y(n_771)
);

AOI221xp5_ASAP7_75t_L g772 ( 
.A1(n_771),
.A2(n_125),
.B1(n_127),
.B2(n_129),
.C(n_130),
.Y(n_772)
);

AOI211xp5_ASAP7_75t_L g773 ( 
.A1(n_772),
.A2(n_131),
.B(n_132),
.C(n_134),
.Y(n_773)
);


endmodule