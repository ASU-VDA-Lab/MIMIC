module real_jpeg_4780_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_525;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_0),
.A2(n_179),
.B1(n_183),
.B2(n_186),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_0),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_0),
.B(n_199),
.C(n_203),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_0),
.B(n_73),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_0),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_0),
.B(n_125),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_0),
.B(n_293),
.Y(n_292)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_1),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_1),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_1),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_1),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_1),
.Y(n_312)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_1),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_55),
.B1(n_59),
.B2(n_62),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_2),
.A2(n_62),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_2),
.A2(n_62),
.B1(n_231),
.B2(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_2),
.A2(n_62),
.B1(n_81),
.B2(n_239),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_3),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_3),
.A2(n_98),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_3),
.A2(n_98),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_4),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g358 ( 
.A(n_4),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_4),
.Y(n_387)
);

INVx6_ASAP7_75t_L g390 ( 
.A(n_4),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_4),
.Y(n_432)
);

BUFx5_ASAP7_75t_L g456 ( 
.A(n_4),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_5),
.A2(n_51),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_5),
.A2(n_51),
.B1(n_239),
.B2(n_418),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_5),
.A2(n_51),
.B1(n_314),
.B2(n_428),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_6),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_8),
.A2(n_210),
.B1(n_215),
.B2(n_216),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_8),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_8),
.A2(n_179),
.B1(n_215),
.B2(n_284),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_8),
.A2(n_162),
.B1(n_215),
.B2(n_394),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_8),
.A2(n_215),
.B1(n_431),
.B2(n_433),
.Y(n_430)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_9),
.Y(n_537)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_12),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_12),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_12),
.A2(n_190),
.B1(n_231),
.B2(n_234),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_12),
.A2(n_190),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_12),
.A2(n_190),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_13),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_13),
.Y(n_233)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_15),
.A2(n_86),
.B1(n_88),
.B2(n_92),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_15),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_15),
.A2(n_92),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g407 ( 
.A1(n_15),
.A2(n_92),
.B1(n_261),
.B2(n_408),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_15),
.A2(n_92),
.B1(n_397),
.B2(n_438),
.Y(n_437)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_17),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_17),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_17),
.A2(n_241),
.B1(n_260),
.B2(n_263),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_17),
.A2(n_241),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_17),
.A2(n_241),
.B1(n_455),
.B2(n_457),
.Y(n_454)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_18),
.A2(n_150),
.B1(n_151),
.B2(n_154),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_18),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_18),
.A2(n_150),
.B1(n_303),
.B2(n_307),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_18),
.A2(n_105),
.B1(n_150),
.B2(n_397),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_18),
.A2(n_150),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_535),
.B(n_538),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_168),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_166),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_141),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_23),
.B(n_141),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_130),
.B2(n_131),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_63),
.C(n_99),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_26),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_27),
.A2(n_52),
.B1(n_54),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_27),
.A2(n_50),
.B1(n_52),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_27),
.A2(n_385),
.B(n_430),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_27),
.A2(n_40),
.B1(n_430),
.B2(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_28),
.A2(n_383),
.B(n_384),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_28),
.B(n_386),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_40),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_39),
.Y(n_362)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_40),
.B(n_186),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_40)
);

INVx6_ASAP7_75t_L g360 ( 
.A(n_41),
.Y(n_360)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g298 ( 
.A(n_43),
.Y(n_298)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_44),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_45),
.Y(n_334)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_46),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_46),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_46),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_46),
.Y(n_365)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_47),
.Y(n_297)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_52),
.A2(n_454),
.B(n_480),
.Y(n_490)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_53),
.B(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_53),
.B(n_149),
.Y(n_479)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_57),
.Y(n_458)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_58),
.Y(n_369)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_63),
.A2(n_99),
.B1(n_100),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_85),
.B1(n_93),
.B2(n_94),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_64),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_64),
.A2(n_85),
.B1(n_93),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_64),
.A2(n_93),
.B1(n_332),
.B2(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_64),
.A2(n_93),
.B1(n_424),
.B2(n_427),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_73),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_67),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_69),
.Y(n_425)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_70),
.Y(n_321)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_73),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

AOI22x1_ASAP7_75t_L g459 ( 
.A1(n_73),
.A2(n_133),
.B1(n_336),
.B2(n_460),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_73),
.A2(n_133),
.B1(n_160),
.B2(n_468),
.Y(n_467)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_81),
.B2(n_83),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_79),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_80),
.Y(n_315)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_80),
.Y(n_420)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_86),
.Y(n_290)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_93),
.B(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_93),
.A2(n_332),
.B(n_335),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_95),
.Y(n_426)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_99),
.B(n_147),
.C(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_99),
.A2(n_100),
.B1(n_157),
.B2(n_158),
.Y(n_524)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_124),
.B(n_126),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_101),
.A2(n_178),
.B(n_187),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_101),
.A2(n_124),
.B1(n_238),
.B2(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_101),
.A2(n_187),
.B(n_283),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_101),
.A2(n_124),
.B1(n_396),
.B2(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_102),
.B(n_188),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_102),
.A2(n_125),
.B1(n_417),
.B2(n_421),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_102),
.A2(n_125),
.B1(n_421),
.B2(n_437),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_102),
.A2(n_125),
.B1(n_437),
.B2(n_471),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_106),
.Y(n_240)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_106),
.Y(n_243)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_113),
.A2(n_238),
.B(n_244),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_120),
.B2(n_122),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_118),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_121),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_121),
.Y(n_262)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_121),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_121),
.Y(n_413)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_124),
.A2(n_244),
.B(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_125),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_126),
.Y(n_471)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_133),
.A2(n_289),
.B(n_295),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_133),
.B(n_336),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_133),
.A2(n_295),
.B(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.C(n_155),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_530)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_146),
.A2(n_147),
.B1(n_524),
.B2(n_525),
.Y(n_523)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_SL g383 ( 
.A1(n_151),
.A2(n_186),
.B(n_366),
.Y(n_383)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_155),
.A2(n_156),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_164),
.Y(n_394)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_519),
.B(n_532),
.Y(n_169)
);

OAI311xp33_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_401),
.A3(n_495),
.B1(n_513),
.C1(n_514),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_350),
.B(n_400),
.Y(n_171)
);

AO21x1_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_323),
.B(n_349),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_277),
.B(n_322),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_247),
.B(n_276),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_207),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_176),
.B(n_207),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_193),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_177),
.A2(n_193),
.B1(n_194),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_177),
.Y(n_274)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

INVx5_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_185),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_186),
.A2(n_219),
.B(n_227),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_SL g289 ( 
.A1(n_186),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_186),
.B(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_206),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_235),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_208),
.B(n_236),
.C(n_246),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_219),
.B(n_227),
.Y(n_208)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_214),
.Y(n_410)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_218),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_219),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_219),
.A2(n_407),
.B1(n_411),
.B2(n_412),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_219),
.A2(n_412),
.B(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_220),
.B(n_230),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_220),
.A2(n_228),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_220),
.A2(n_302),
.B1(n_340),
.B2(n_346),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_220),
.A2(n_375),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_223),
.Y(n_347)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_223),
.Y(n_451)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_233),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_245),
.B2(n_246),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp33_ASAP7_75t_SL g319 ( 
.A(n_242),
.B(n_320),
.Y(n_319)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_269),
.B(n_275),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_257),
.B(n_268),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_256),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_253),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_255),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_267),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_267),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_265),
.B(n_266),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_301),
.B(n_310),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_273),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_279),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_299),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_287),
.B2(n_288),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_287),
.C(n_299),
.Y(n_324)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI32xp33_ASAP7_75t_L g313 ( 
.A1(n_292),
.A2(n_314),
.A3(n_315),
.B1(n_316),
.B2(n_319),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_313),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_313),
.Y(n_329)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_324),
.B(n_325),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_330),
.B2(n_348),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_329),
.C(n_348),
.Y(n_351)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_330),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_337),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_331),
.B(n_338),
.C(n_339),
.Y(n_377)
);

OAI32xp33_ASAP7_75t_L g356 ( 
.A1(n_334),
.A2(n_357),
.A3(n_359),
.B1(n_361),
.B2(n_366),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_351),
.B(n_352),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_380),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_353)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_370),
.B2(n_371),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_356),
.B(n_370),
.Y(n_491)
);

INVx8_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

INVx6_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_377),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_377),
.B(n_378),
.C(n_380),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_382),
.B1(n_391),
.B2(n_399),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_381),
.B(n_392),
.C(n_395),
.Y(n_504)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx8_ASAP7_75t_L g433 ( 
.A(n_390),
.Y(n_433)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_391),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_393),
.Y(n_493)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NAND2xp33_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_481),
.Y(n_401)
);

A2O1A1Ixp33_ASAP7_75t_SL g514 ( 
.A1(n_402),
.A2(n_481),
.B(n_515),
.C(n_518),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_461),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_403),
.B(n_461),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_434),
.C(n_444),
.Y(n_403)
);

FAx1_ASAP7_75t_SL g494 ( 
.A(n_404),
.B(n_434),
.CI(n_444),
.CON(n_494),
.SN(n_494)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_422),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_405),
.B(n_423),
.C(n_429),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_416),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_406),
.B(n_416),
.Y(n_487)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_407),
.Y(n_449)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_417),
.Y(n_447)
);

INVx4_ASAP7_75t_SL g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_420),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_429),
.Y(n_422)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_424),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_427),
.Y(n_468)
);

INVx8_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_435),
.A2(n_436),
.B1(n_440),
.B2(n_443),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_440),
.Y(n_475)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_440),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_440),
.A2(n_443),
.B1(n_477),
.B2(n_478),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_440),
.A2(n_475),
.B(n_478),
.Y(n_522)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_452),
.C(n_459),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_445),
.B(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_446),
.B(n_448),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_446),
.B(n_448),
.Y(n_503)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_452),
.A2(n_453),
.B1(n_459),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_459),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_462),
.B(n_465),
.C(n_473),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_464),
.A2(n_465),
.B1(n_473),
.B2(n_474),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_466),
.A2(n_469),
.B(n_472),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_467),
.B(n_470),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

FAx1_ASAP7_75t_SL g521 ( 
.A(n_472),
.B(n_522),
.CI(n_523),
.CON(n_521),
.SN(n_521)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_472),
.B(n_522),
.C(n_523),
.Y(n_531)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_494),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_482),
.B(n_494),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_487),
.C(n_488),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_483),
.A2(n_484),
.B1(n_487),
.B2(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_487),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_506),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_491),
.C(n_492),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_489),
.A2(n_490),
.B1(n_492),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_492),
.Y(n_501)
);

BUFx24_ASAP7_75t_SL g542 ( 
.A(n_494),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_508),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_497),
.A2(n_516),
.B(n_517),
.Y(n_515)
);

NOR2x1_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_505),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_498),
.B(n_505),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_502),
.C(n_504),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_511),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_502),
.A2(n_503),
.B1(n_504),
.B2(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_504),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_510),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_510),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_527),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_526),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_526),
.Y(n_533)
);

BUFx24_ASAP7_75t_SL g543 ( 
.A(n_521),
.Y(n_543)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_524),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_527),
.A2(n_533),
.B(n_534),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_528),
.B(n_531),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_528),
.B(n_531),
.Y(n_534)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

BUFx4f_ASAP7_75t_SL g535 ( 
.A(n_536),
.Y(n_535)
);

BUFx12f_ASAP7_75t_L g539 ( 
.A(n_536),
.Y(n_539)
);

INVx13_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_540),
.Y(n_538)
);


endmodule