module real_jpeg_29203_n_31 (n_17, n_8, n_0, n_157, n_21, n_2, n_29, n_10, n_9, n_12, n_154, n_156, n_152, n_24, n_6, n_28, n_153, n_151, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_150, n_1, n_26, n_27, n_20, n_19, n_30, n_158, n_149, n_16, n_15, n_13, n_155, n_31);

input n_17;
input n_8;
input n_0;
input n_157;
input n_21;
input n_2;
input n_29;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_24;
input n_6;
input n_28;
input n_153;
input n_151;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_150;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_30;
input n_158;
input n_149;
input n_16;
input n_15;
input n_13;
input n_155;

output n_31;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_0),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_1),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_3),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_4),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_4),
.B(n_56),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_6),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_6),
.B(n_121),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_7),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_8),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_8),
.B(n_112),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_9),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_11),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_49),
.C(n_133),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_13),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_13),
.B(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_14),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_15),
.B(n_60),
.C(n_124),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_16),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_16),
.B(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_17),
.B(n_70),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_18),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_20),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_20),
.B(n_51),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_22),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_23),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_23),
.B(n_46),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_23),
.B(n_138),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_23),
.B(n_141),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_23),
.B(n_41),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_24),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_25),
.B(n_95),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_26),
.B(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_27),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_28),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_29),
.B(n_64),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_29),
.B(n_64),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_30),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_39),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_35),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_35),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_35),
.B(n_113),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_35),
.B(n_117),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_35),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_35),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_35),
.B(n_139),
.Y(n_138)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_36),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_37),
.A2(n_137),
.B(n_140),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B(n_147),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_136),
.B(n_144),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B(n_135),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_132),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_127),
.B(n_131),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B(n_126),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_58),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_120),
.B(n_123),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_115),
.B(n_119),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_67),
.B(n_111),
.C(n_114),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_65),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_110),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B(n_109),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_104),
.B(n_108),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B(n_103),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_98),
.B(n_102),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_94),
.B(n_97),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_93),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_85),
.B(n_88),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_96),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_91),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_99),
.B(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_106),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_118),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_130),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_149),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_150),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_151),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_152),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_153),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_154),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_155),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_156),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_157),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_158),
.Y(n_113)
);


endmodule