module fake_jpeg_20076_n_175 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_38),
.Y(n_43)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_25),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_23),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_25),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_17),
.B1(n_16),
.B2(n_18),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_18),
.Y(n_71)
);

OAI32xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_32),
.A3(n_38),
.B1(n_19),
.B2(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_77),
.Y(n_78)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_36),
.B1(n_39),
.B2(n_38),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_63),
.B1(n_67),
.B2(n_72),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_39),
.B1(n_35),
.B2(n_32),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_39),
.B1(n_35),
.B2(n_33),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_56),
.B(n_31),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_73),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_39),
.B1(n_34),
.B2(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_20),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_93),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_20),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_28),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_94),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_56),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_19),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_50),
.B1(n_16),
.B2(n_44),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_97),
.B1(n_27),
.B2(n_24),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_28),
.B1(n_22),
.B2(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_103),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_69),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_86),
.B(n_82),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_62),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_67),
.B1(n_59),
.B2(n_60),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_67),
.B1(n_66),
.B2(n_65),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_27),
.B1(n_15),
.B2(n_64),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_84),
.B(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_72),
.B1(n_50),
.B2(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_114),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_72),
.C(n_56),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_26),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_42),
.B1(n_45),
.B2(n_21),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_121),
.B(n_126),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_95),
.B(n_87),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_125),
.B(n_130),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_87),
.B(n_79),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_85),
.C(n_15),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_81),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_31),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_79),
.B(n_81),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_113),
.B1(n_109),
.B2(n_98),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_133),
.B1(n_141),
.B2(n_142),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_120),
.A2(n_101),
.B1(n_42),
.B2(n_45),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_101),
.C(n_51),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_140),
.C(n_127),
.Y(n_145)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_122),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_21),
.B1(n_26),
.B2(n_3),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_51),
.B1(n_26),
.B2(n_13),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_119),
.C(n_123),
.Y(n_150)
);

AOI31xp67_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_142),
.A3(n_133),
.B(n_115),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_116),
.C(n_130),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_155),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_146),
.B(n_147),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_4),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_154),
.A2(n_150),
.B1(n_151),
.B2(n_117),
.Y(n_161)
);

NAND4xp25_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_51),
.C(n_2),
.D(n_3),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_162),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_12),
.B(n_11),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_168),
.C(n_162),
.Y(n_169)
);

NOR4xp25_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_152),
.C(n_158),
.D(n_10),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_167),
.B(n_7),
.Y(n_170)
);

AOI31xp33_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_11),
.A3(n_5),
.B(n_6),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_5),
.B(n_6),
.Y(n_171)
);

INVxp33_ASAP7_75t_SL g173 ( 
.A(n_170),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_5),
.B(n_6),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_172),
.Y(n_175)
);


endmodule