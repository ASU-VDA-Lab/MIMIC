module fake_aes_2633_n_42 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_42);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_30;
wire n_16;
wire n_25;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
INVx1_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
OA21x2_ASAP7_75t_L g17 ( .A1(n_8), .A2(n_10), .B(n_2), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_15), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_1), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_9), .Y(n_21) );
NOR2x1_ASAP7_75t_L g22 ( .A(n_13), .B(n_4), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_3), .B(n_0), .Y(n_23) );
BUFx6f_ASAP7_75t_L g24 ( .A(n_11), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g25 ( .A1(n_19), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_21), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_19), .A2(n_6), .B1(n_7), .B2(n_18), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_18), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_23), .A2(n_22), .B1(n_20), .B2(n_16), .Y(n_29) );
AOI21xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_21), .B(n_17), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_28), .B(n_17), .Y(n_31) );
INVx4_ASAP7_75t_L g32 ( .A(n_27), .Y(n_32) );
INVx5_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_30), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
AND2x2_ASAP7_75t_L g36 ( .A(n_33), .B(n_32), .Y(n_36) );
NOR2xp33_ASAP7_75t_L g37 ( .A(n_36), .B(n_32), .Y(n_37) );
AOI221xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_34), .B1(n_35), .B2(n_25), .C(n_26), .Y(n_38) );
AND3x4_ASAP7_75t_L g39 ( .A(n_38), .B(n_33), .C(n_24), .Y(n_39) );
HB1xp67_ASAP7_75t_L g40 ( .A(n_39), .Y(n_40) );
INVx2_ASAP7_75t_L g41 ( .A(n_40), .Y(n_41) );
INVxp67_ASAP7_75t_L g42 ( .A(n_41), .Y(n_42) );
endmodule