module real_jpeg_15777_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_1),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_1),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_2),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_2),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_3),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_3),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_3),
.A2(n_114),
.B1(n_250),
.B2(n_253),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_3),
.A2(n_114),
.B1(n_374),
.B2(n_376),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_3),
.A2(n_114),
.B1(n_340),
.B2(n_447),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_4),
.A2(n_267),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_4),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_4),
.A2(n_321),
.B1(n_420),
.B2(n_432),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_5),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_5),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_6),
.A2(n_196),
.B1(n_199),
.B2(n_202),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_6),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_6),
.A2(n_202),
.B1(n_416),
.B2(n_419),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_6),
.A2(n_202),
.B1(n_474),
.B2(n_476),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_7),
.Y(n_109)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_7),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g383 ( 
.A(n_7),
.Y(n_383)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_7),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_8),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_8),
.A2(n_63),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_8),
.A2(n_41),
.B1(n_63),
.B2(n_375),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_8),
.A2(n_63),
.B1(n_483),
.B2(n_485),
.Y(n_482)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_9),
.Y(n_343)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_9),
.Y(n_350)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_25),
.A3(n_31),
.B1(n_34),
.B2(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_10),
.A2(n_38),
.B1(n_143),
.B2(n_147),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_10),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_10),
.B(n_117),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_10),
.B(n_282),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_10),
.B(n_237),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_10),
.A2(n_323),
.A3(n_326),
.B1(n_331),
.B2(n_338),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_10),
.A2(n_38),
.B1(n_359),
.B2(n_361),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_154),
.B1(n_159),
.B2(n_161),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_11),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_11),
.A2(n_161),
.B1(n_239),
.B2(n_245),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_11),
.A2(n_161),
.B1(n_284),
.B2(n_288),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_11),
.A2(n_161),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_12),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_13),
.A2(n_67),
.B1(n_72),
.B2(n_73),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_13),
.A2(n_72),
.B1(n_382),
.B2(n_384),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_13),
.A2(n_72),
.B1(n_441),
.B2(n_443),
.Y(n_440)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_15),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_15),
.Y(n_352)
);

BUFx8_ASAP7_75t_L g354 ( 
.A(n_15),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_458),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_391),
.B(n_454),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_309),
.B(n_390),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_214),
.B(n_308),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_163),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_22),
.B(n_163),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_78),
.C(n_115),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_23),
.B(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_24),
.B(n_48),
.Y(n_165)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_29),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_29),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_30),
.Y(n_134)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_30),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_30),
.Y(n_184)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_32),
.Y(n_174)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_38),
.B(n_91),
.Y(n_225)
);

OAI21xp33_ASAP7_75t_SL g234 ( 
.A1(n_38),
.A2(n_225),
.B(n_235),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_38),
.A2(n_50),
.B1(n_281),
.B2(n_283),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_38),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_43),
.Y(n_158)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_43),
.Y(n_325)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_58),
.B(n_65),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_49),
.A2(n_265),
.B1(n_274),
.B2(n_275),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_49),
.A2(n_195),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_49),
.A2(n_65),
.B(n_319),
.Y(n_412)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_50),
.B(n_66),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_50),
.A2(n_249),
.B(n_255),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_50),
.A2(n_266),
.B1(n_283),
.B2(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_50),
.A2(n_59),
.B(n_464),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_53),
.Y(n_201)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_56),
.Y(n_298)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_59),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_60),
.Y(n_320)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_61),
.Y(n_254)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_61),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_62),
.Y(n_271)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_64),
.Y(n_221)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_71),
.Y(n_198)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_71),
.Y(n_252)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_71),
.Y(n_287)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_77),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_78),
.B(n_115),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_92),
.B1(n_99),
.B2(n_110),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_79),
.A2(n_169),
.B(n_380),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_79),
.A2(n_92),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g467 ( 
.A1(n_79),
.A2(n_380),
.B(n_431),
.Y(n_467)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_80),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_80),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_80),
.A2(n_100),
.B1(n_237),
.B2(n_238),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_80),
.B(n_381),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_92),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_87),
.B2(n_91),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_83),
.Y(n_220)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_84),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_86),
.Y(n_224)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_92),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_92),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_103),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_103),
.Y(n_433)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_104),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_105),
.A2(n_106),
.B1(n_208),
.B2(n_212),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_105),
.A2(n_106),
.B1(n_267),
.B2(n_272),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_105),
.A2(n_106),
.B1(n_369),
.B2(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_142),
.B1(n_153),
.B2(n_162),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_116),
.A2(n_162),
.B1(n_207),
.B2(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_116),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_116),
.A2(n_408),
.B(n_439),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_116),
.A2(n_162),
.B1(n_472),
.B2(n_473),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_127),
.Y(n_116)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_117),
.B(n_440),
.Y(n_439)
);

AO22x2_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_132),
.B1(n_135),
.B2(n_138),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_134),
.Y(n_444)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_141),
.Y(n_337)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_141),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_144),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AO22x2_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_153),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_204)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_158),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_162),
.B(n_408),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_175),
.B1(n_176),
.B2(n_213),
.Y(n_163)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_165),
.B(n_166),
.C(n_175),
.Y(n_389)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_204),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_187),
.B2(n_188),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_178),
.B(n_188),
.C(n_204),
.Y(n_313)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_180),
.B(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_180),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_180),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_180),
.B(n_482),
.Y(n_481)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g357 ( 
.A(n_183),
.Y(n_357)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_184),
.Y(n_442)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_195),
.B(n_203),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_SL g258 ( 
.A(n_192),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_192),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_194),
.Y(n_318)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_198),
.Y(n_288)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_203),
.B(n_256),
.Y(n_428)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_303),
.B(n_307),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_262),
.B(n_302),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_247),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_217),
.B(n_247),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_232),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_218),
.A2(n_232),
.B1(n_233),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_221),
.A3(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_237),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_237),
.B(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_259),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_248),
.B(n_260),
.C(n_261),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

OAI21x1_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_278),
.B(n_301),
.Y(n_262)
);

NOR2x1_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_276),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_276),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_269),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_294),
.B(n_300),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_289),
.Y(n_279)
);

INVx6_ASAP7_75t_L g465 ( 
.A(n_281),
.Y(n_465)
);

BUFx12f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_299),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_299),
.Y(n_300)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_389),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_310),
.B(n_389),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_344),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_313),
.B(n_314),
.C(n_344),
.Y(n_451)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_322),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_316),
.B(n_322),
.Y(n_409)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_329),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_329),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_337),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_371),
.Y(n_344)
);

MAJx2_ASAP7_75t_L g410 ( 
.A(n_345),
.B(n_372),
.C(n_379),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_358),
.B1(n_365),
.B2(n_370),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_346),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_346),
.A2(n_370),
.B1(n_401),
.B2(n_446),
.Y(n_445)
);

OAI21x1_ASAP7_75t_SL g480 ( 
.A1(n_346),
.A2(n_446),
.B(n_481),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_348),
.A2(n_351),
.B1(n_353),
.B2(n_355),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx12f_ASAP7_75t_L g360 ( 
.A(n_352),
.Y(n_360)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_354),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_363),
.Y(n_367)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_364),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_379),
.Y(n_371)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_450),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_424),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_394),
.B(n_424),
.C(n_457),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_410),
.C(n_411),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_395),
.B(n_453),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_409),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_404),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_404),
.C(n_409),
.Y(n_425)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_406),
.B(n_407),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_410),
.B(n_411),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_413),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_423),
.Y(n_413)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_415),
.Y(n_430)
);

BUFx2_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx5_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_425),
.B(n_434),
.C(n_449),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_434),
.B1(n_435),
.B2(n_449),
.Y(n_426)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_427),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_428),
.B(n_429),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_435),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_436),
.B(n_491),
.C(n_492),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_445),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_438),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_445),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_452),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_455),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_R g458 ( 
.A(n_459),
.B(n_495),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_494),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_494),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_461),
.A2(n_489),
.B1(n_490),
.B2(n_493),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_461),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_469),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_466),
.B1(n_467),
.B2(n_468),
.Y(n_462)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_463),
.Y(n_468)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

XNOR2x1_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_488),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_480),
.Y(n_470)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);


endmodule