module fake_jpeg_2455_n_586 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_586);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_586;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_1),
.B(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_59),
.Y(n_171)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_62),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_64),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_65),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_66),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_67),
.Y(n_209)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_31),
.B(n_9),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_83),
.Y(n_129)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_25),
.B(n_9),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_76),
.B(n_117),
.Y(n_183)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_81),
.Y(n_182)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g211 ( 
.A(n_82),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_8),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_84),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_86),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_8),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_41),
.B(n_18),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_87),
.B(n_89),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_88),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_8),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_90),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_22),
.B(n_8),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_102),
.Y(n_142)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_93),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_94),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_95),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_25),
.A2(n_7),
.B1(n_16),
.B2(n_14),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_96),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_203)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

BUFx4f_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_101),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_29),
.B(n_7),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_45),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_107),
.B(n_108),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_29),
.B(n_7),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_42),
.B(n_10),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_118),
.Y(n_134)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

INVx6_ASAP7_75t_SL g180 ( 
.A(n_117),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_44),
.B(n_10),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_33),
.Y(n_121)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_19),
.Y(n_122)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_35),
.Y(n_125)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_128),
.B(n_163),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_59),
.A2(n_45),
.B1(n_36),
.B2(n_47),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_131),
.A2(n_137),
.B1(n_140),
.B2(n_156),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_59),
.A2(n_36),
.B1(n_47),
.B2(n_35),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_36),
.B1(n_47),
.B2(n_35),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_82),
.A2(n_47),
.B1(n_42),
.B2(n_55),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_144),
.A2(n_154),
.B1(n_174),
.B2(n_177),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_97),
.A2(n_47),
.B1(n_55),
.B2(n_48),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_90),
.A2(n_44),
.B1(n_46),
.B2(n_19),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_79),
.A2(n_46),
.B1(n_24),
.B2(n_53),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_158),
.A2(n_168),
.B(n_203),
.C(n_132),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_101),
.B(n_48),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_159),
.B(n_132),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_125),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_SL g165 ( 
.A1(n_119),
.A2(n_53),
.B(n_24),
.Y(n_165)
);

AOI32xp33_ASAP7_75t_L g258 ( 
.A1(n_165),
.A2(n_188),
.A3(n_11),
.B1(n_16),
.B2(n_17),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_64),
.A2(n_57),
.B1(n_54),
.B2(n_39),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_74),
.B(n_13),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_169),
.B(n_173),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_99),
.B(n_13),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_123),
.A2(n_67),
.B1(n_120),
.B2(n_111),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_63),
.A2(n_56),
.B1(n_49),
.B2(n_54),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_210),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_72),
.B(n_121),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_184),
.B(n_204),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_80),
.A2(n_56),
.B(n_49),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

INVx6_ASAP7_75t_SL g191 ( 
.A(n_112),
.Y(n_191)
);

INVx4_ASAP7_75t_SL g245 ( 
.A(n_191),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_66),
.A2(n_109),
.B1(n_81),
.B2(n_103),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_198),
.A2(n_127),
.B1(n_152),
.B2(n_136),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_104),
.B(n_14),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_69),
.B(n_16),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_4),
.Y(n_251)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_93),
.B(n_56),
.C(n_49),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_94),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_134),
.B(n_2),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_214),
.B(n_217),
.Y(n_317)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_148),
.B(n_100),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_180),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_218),
.B(n_219),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_184),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_164),
.Y(n_221)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_221),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_181),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_222),
.B(n_235),
.Y(n_307)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_223),
.Y(n_291)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_224),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_175),
.A2(n_96),
.B1(n_98),
.B2(n_57),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_183),
.A2(n_56),
.B1(n_49),
.B2(n_39),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_228),
.A2(n_261),
.B1(n_280),
.B2(n_281),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_126),
.A2(n_49),
.B1(n_56),
.B2(n_5),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_229),
.Y(n_316)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_230),
.Y(n_300)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_231),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_126),
.A2(n_168),
.B1(n_204),
.B2(n_142),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_233),
.A2(n_242),
.B1(n_248),
.B2(n_283),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_3),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_234),
.B(n_254),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_238),
.B(n_243),
.Y(n_321)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_239),
.Y(n_326)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_240),
.Y(n_327)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_160),
.Y(n_241)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_167),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_133),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_169),
.B(n_3),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_244),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_201),
.A2(n_4),
.B1(n_5),
.B2(n_10),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_249),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_250),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_251),
.B(n_262),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_146),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_252),
.Y(n_292)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_135),
.B(n_5),
.Y(n_254)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_178),
.Y(n_257)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_267),
.Y(n_310)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_187),
.Y(n_259)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_138),
.B(n_11),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_260),
.B(n_278),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_130),
.A2(n_11),
.B1(n_129),
.B2(n_137),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_133),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_178),
.Y(n_263)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_263),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_193),
.Y(n_265)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_265),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_266),
.B(n_214),
.Y(n_342)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

OA22x2_ASAP7_75t_L g333 ( 
.A1(n_268),
.A2(n_272),
.B1(n_253),
.B2(n_267),
.Y(n_333)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_270),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_173),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_139),
.B(n_145),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_271),
.B(n_273),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_127),
.A2(n_152),
.B1(n_136),
.B2(n_196),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_157),
.B(n_153),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_147),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_274),
.B(n_275),
.Y(n_341)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_172),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_143),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

NOR2x1_ASAP7_75t_R g277 ( 
.A(n_176),
.B(n_189),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_277),
.B(n_244),
.C(n_232),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_149),
.B(n_151),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_207),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_279),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_140),
.A2(n_158),
.B1(n_131),
.B2(n_156),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_166),
.A2(n_182),
.B1(n_200),
.B2(n_195),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_143),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_282),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_155),
.B(n_162),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_284),
.B(n_286),
.Y(n_335)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_141),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_285),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_157),
.B(n_192),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_141),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_287),
.A2(n_263),
.B1(n_257),
.B2(n_245),
.Y(n_336)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_225),
.B(n_150),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_294),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_225),
.A2(n_196),
.B1(n_203),
.B2(n_209),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_297),
.A2(n_298),
.B1(n_309),
.B2(n_319),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_225),
.A2(n_203),
.B1(n_209),
.B2(n_199),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_255),
.A2(n_199),
.B1(n_166),
.B2(n_182),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_301),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_255),
.A2(n_217),
.B1(n_268),
.B2(n_246),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_306),
.A2(n_314),
.B1(n_283),
.B2(n_236),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_280),
.A2(n_200),
.B1(n_186),
.B2(n_197),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_283),
.A2(n_186),
.B1(n_197),
.B2(n_150),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_228),
.A2(n_197),
.B1(n_186),
.B2(n_150),
.Y(n_319)
);

AND2x2_ASAP7_75t_SL g320 ( 
.A(n_278),
.B(n_284),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_320),
.B(n_323),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_SL g323 ( 
.A(n_277),
.B(n_260),
.Y(n_323)
);

NOR3xp33_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_282),
.C(n_276),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_333),
.A2(n_283),
.B1(n_236),
.B2(n_245),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_254),
.A2(n_237),
.B1(n_220),
.B2(n_226),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_339),
.A2(n_241),
.B1(n_224),
.B2(n_231),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_342),
.B(n_279),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_344),
.A2(n_346),
.B1(n_353),
.B2(n_372),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_294),
.B(n_234),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_345),
.B(n_349),
.C(n_356),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_288),
.A2(n_320),
.B1(n_297),
.B2(n_306),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_341),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_347),
.B(n_371),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_348),
.A2(n_365),
.B(n_334),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_294),
.B(n_216),
.C(n_236),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_304),
.B(n_296),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_351),
.B(n_352),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_288),
.A2(n_236),
.B1(n_244),
.B2(n_240),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_295),
.A2(n_238),
.B(n_235),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_354),
.A2(n_340),
.B(n_328),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_303),
.B(n_275),
.C(n_285),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_332),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_327),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_215),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_360),
.B(n_361),
.Y(n_407)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_329),
.Y(n_362)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_329),
.Y(n_363)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_363),
.Y(n_400)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_364),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_316),
.A2(n_256),
.B1(n_265),
.B2(n_230),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_291),
.Y(n_366)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_341),
.Y(n_368)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_368),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_221),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_369),
.B(n_375),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_370),
.A2(n_376),
.B1(n_381),
.B2(n_384),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_341),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_298),
.A2(n_259),
.B1(n_264),
.B2(n_250),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_295),
.A2(n_223),
.B1(n_239),
.B2(n_314),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_373),
.A2(n_385),
.B1(n_313),
.B2(n_293),
.Y(n_412)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_343),
.Y(n_374)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_317),
.B(n_320),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_343),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_324),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_377),
.B(n_378),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_324),
.B(n_330),
.Y(n_378)
);

AOI21xp33_ASAP7_75t_L g379 ( 
.A1(n_310),
.A2(n_296),
.B(n_312),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_379),
.B(n_292),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_335),
.B(n_323),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_310),
.Y(n_391)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_335),
.A2(n_309),
.B1(n_310),
.B2(n_303),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_331),
.A2(n_316),
.B(n_321),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_386),
.A2(n_319),
.B(n_291),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_404),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_386),
.A2(n_307),
.B(n_312),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_392),
.A2(n_395),
.B(n_399),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_328),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_396),
.B(n_397),
.C(n_405),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_375),
.Y(n_397)
);

NAND2x1_ASAP7_75t_SL g402 ( 
.A(n_383),
.B(n_300),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_402),
.A2(n_403),
.B(n_411),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_380),
.A2(n_328),
.B(n_342),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_345),
.B(n_290),
.Y(n_405)
);

OA22x2_ASAP7_75t_L g409 ( 
.A1(n_344),
.A2(n_333),
.B1(n_302),
.B2(n_300),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_409),
.B(n_412),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_383),
.B(n_302),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_410),
.B(n_414),
.C(n_418),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_353),
.A2(n_346),
.B1(n_382),
.B2(n_355),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_360),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_299),
.C(n_292),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_385),
.A2(n_333),
.B1(n_322),
.B2(n_311),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_419),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_421),
.A2(n_350),
.B(n_354),
.Y(n_428)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_387),
.Y(n_426)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_426),
.Y(n_481)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_427),
.B(n_432),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_428),
.A2(n_418),
.B(n_402),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_393),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_429),
.B(n_434),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_411),
.A2(n_367),
.B1(n_369),
.B2(n_373),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_430),
.A2(n_442),
.B1(n_453),
.B2(n_410),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g431 ( 
.A(n_407),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_431),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_401),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_349),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_433),
.B(n_363),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_402),
.A2(n_350),
.B(n_355),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_356),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_439),
.C(n_445),
.Y(n_459)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_408),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_438),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_412),
.A2(n_372),
.B1(n_366),
.B2(n_364),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_437),
.A2(n_441),
.B1(n_446),
.B2(n_452),
.Y(n_475)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_368),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_394),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_443),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_420),
.A2(n_371),
.B1(n_347),
.B2(n_370),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_390),
.A2(n_333),
.B1(n_337),
.B2(n_311),
.Y(n_442)
);

INVxp33_ASAP7_75t_L g443 ( 
.A(n_389),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_401),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_450),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_396),
.B(n_376),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_407),
.A2(n_374),
.B1(n_358),
.B2(n_359),
.Y(n_446)
);

BUFx5_ASAP7_75t_L g448 ( 
.A(n_395),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_448),
.Y(n_456)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_400),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_416),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_390),
.A2(n_415),
.B1(n_399),
.B2(n_414),
.Y(n_453)
);

A2O1A1O1Ixp25_ASAP7_75t_L g457 ( 
.A1(n_423),
.A2(n_417),
.B(n_415),
.C(n_403),
.D(n_392),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_457),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_405),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_462),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_453),
.Y(n_460)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_460),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_449),
.A2(n_409),
.B1(n_419),
.B2(n_421),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_461),
.A2(n_476),
.B1(n_442),
.B2(n_438),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_391),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_463),
.A2(n_470),
.B1(n_441),
.B2(n_452),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_433),
.B(n_397),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_464),
.B(n_472),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_465),
.A2(n_422),
.B(n_425),
.Y(n_483)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_398),
.C(n_406),
.Y(n_467)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_467),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_409),
.C(n_340),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_482),
.C(n_425),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_431),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_469),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_449),
.A2(n_409),
.B1(n_398),
.B2(n_388),
.Y(n_470)
);

AND2x2_ASAP7_75t_SL g471 ( 
.A(n_447),
.B(n_362),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_471),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_447),
.A2(n_406),
.B1(n_357),
.B2(n_337),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_423),
.B(n_384),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_480),
.Y(n_491)
);

AO22x1_ASAP7_75t_L g479 ( 
.A1(n_447),
.A2(n_381),
.B1(n_357),
.B2(n_332),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_430),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_451),
.B(n_289),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_445),
.B(n_289),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_483),
.B(n_487),
.Y(n_523)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_485),
.Y(n_509)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_486),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_474),
.A2(n_422),
.B(n_434),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_488),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_424),
.C(n_444),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_489),
.B(n_490),
.C(n_497),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_424),
.C(n_432),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g494 ( 
.A(n_455),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_494),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_495),
.A2(n_499),
.B1(n_500),
.B2(n_471),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_427),
.Y(n_496)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_496),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_458),
.B(n_426),
.C(n_436),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_461),
.A2(n_448),
.B1(n_450),
.B2(n_440),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_456),
.A2(n_428),
.B1(n_293),
.B2(n_313),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_466),
.B(n_305),
.Y(n_503)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_503),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_326),
.C(n_318),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_464),
.C(n_462),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_473),
.A2(n_308),
.B(n_334),
.Y(n_505)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_505),
.Y(n_521)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_454),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_506),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_502),
.B(n_477),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_510),
.B(n_512),
.Y(n_534)
);

FAx1_ASAP7_75t_SL g512 ( 
.A(n_507),
.B(n_457),
.CI(n_468),
.CON(n_512),
.SN(n_512)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_514),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_519),
.B(n_520),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_489),
.B(n_472),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_496),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_522),
.B(n_525),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_465),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_524),
.B(n_492),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_506),
.B(n_478),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_490),
.B(n_484),
.C(n_491),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_526),
.B(n_487),
.C(n_497),
.Y(n_529)
);

INVx11_ASAP7_75t_L g527 ( 
.A(n_511),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_527),
.A2(n_528),
.B1(n_537),
.B2(n_517),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_521),
.A2(n_516),
.B1(n_509),
.B2(n_499),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_539),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_521),
.A2(n_495),
.B1(n_463),
.B2(n_486),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_530),
.A2(n_540),
.B1(n_514),
.B2(n_501),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_491),
.C(n_504),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_531),
.B(n_535),
.C(n_526),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_493),
.C(n_492),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_513),
.B(n_498),
.Y(n_536)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_536),
.Y(n_552)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_516),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_513),
.B(n_485),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_509),
.A2(n_471),
.B1(n_501),
.B2(n_488),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_541),
.B(n_519),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_542),
.B(n_543),
.Y(n_556)
);

BUFx24_ASAP7_75t_SL g544 ( 
.A(n_534),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_544),
.B(n_538),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_546),
.B(n_547),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_520),
.C(n_523),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_533),
.A2(n_517),
.B1(n_515),
.B2(n_483),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_548),
.A2(n_551),
.B1(n_530),
.B2(n_537),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_528),
.A2(n_515),
.B(n_508),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_549),
.B(n_550),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_540),
.A2(n_508),
.B(n_503),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_533),
.A2(n_470),
.B1(n_500),
.B2(n_512),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_553),
.B(n_532),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_529),
.B(n_523),
.C(n_524),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_554),
.B(n_532),
.C(n_535),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_558),
.B(n_559),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_543),
.A2(n_536),
.B1(n_534),
.B2(n_473),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_560),
.B(n_562),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_561),
.B(n_546),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_545),
.B(n_481),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_563),
.B(n_550),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_552),
.A2(n_512),
.B(n_505),
.Y(n_564)
);

AO21x1_ASAP7_75t_L g571 ( 
.A1(n_564),
.A2(n_541),
.B(n_551),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_565),
.A2(n_568),
.B(n_556),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_557),
.B(n_549),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_569),
.A2(n_571),
.B(n_572),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_555),
.A2(n_547),
.B(n_554),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_570),
.A2(n_553),
.B(n_556),
.Y(n_574)
);

A2O1A1Ixp33_ASAP7_75t_SL g572 ( 
.A1(n_557),
.A2(n_548),
.B(n_527),
.C(n_476),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_567),
.B(n_562),
.C(n_561),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_573),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_574),
.A2(n_569),
.B(n_572),
.Y(n_579)
);

NAND2x1_ASAP7_75t_SL g578 ( 
.A(n_576),
.B(n_577),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_566),
.B(n_475),
.C(n_482),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_579),
.A2(n_479),
.B(n_318),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_578),
.B(n_575),
.Y(n_581)
);

NOR3xp33_ASAP7_75t_L g583 ( 
.A(n_581),
.B(n_582),
.C(n_580),
.Y(n_583)
);

A2O1A1Ixp33_ASAP7_75t_L g584 ( 
.A1(n_583),
.A2(n_479),
.B(n_305),
.C(n_325),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_584),
.B(n_308),
.C(n_326),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_585),
.B(n_325),
.Y(n_586)
);


endmodule