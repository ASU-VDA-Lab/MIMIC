module fake_jpeg_30680_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_1),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx4f_ASAP7_75t_SL g12 ( 
.A(n_4),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_19),
.Y(n_24)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_15),
.B1(n_5),
.B2(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_8),
.B(n_0),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_13),
.B(n_17),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_12),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_27),
.C(n_28),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_12),
.C(n_9),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_12),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_24),
.B2(n_25),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_33),
.A2(n_32),
.B(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_34),
.B(n_5),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_9),
.Y(n_36)
);


endmodule