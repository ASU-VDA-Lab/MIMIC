module fake_netlist_5_2518_n_1201 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1201);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1201;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_1194;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_1178;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_523;
wire n_268;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_1191;
wire n_1198;
wire n_721;
wire n_998;
wire n_1157;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_501;
wire n_284;
wire n_245;
wire n_823;
wire n_983;
wire n_725;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_677;
wire n_244;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_1179;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_624;
wire n_252;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_1195;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_1090;
wire n_1200;
wire n_307;
wire n_633;
wire n_1192;
wire n_439;
wire n_530;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1185;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_1182;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_579;
wire n_250;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_1163;
wire n_519;
wire n_406;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_1172;
wire n_976;
wire n_1095;
wire n_1096;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_1045;
wire n_297;
wire n_833;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_995;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_1176;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_1149;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_962;
wire n_436;
wire n_930;
wire n_580;
wire n_290;
wire n_221;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1188;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_1165;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_1177;
wire n_680;
wire n_974;
wire n_395;
wire n_553;
wire n_432;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_1159;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_482;
wire n_517;
wire n_342;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_571;
wire n_477;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_1193;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_1197;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1187;
wire n_1015;
wire n_1000;
wire n_1140;
wire n_891;
wire n_466;
wire n_239;
wire n_1164;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_846;
wire n_586;
wire n_874;
wire n_465;
wire n_1058;
wire n_358;
wire n_838;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_1190;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_1052;
wire n_963;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_1175;
wire n_861;
wire n_534;
wire n_948;
wire n_1183;
wire n_1076;
wire n_884;
wire n_1091;
wire n_345;
wire n_210;
wire n_944;
wire n_899;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_679;
wire n_425;
wire n_513;
wire n_237;
wire n_407;
wire n_527;
wire n_647;
wire n_710;
wire n_707;
wire n_832;
wire n_695;
wire n_795;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_1072;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_1027;
wire n_490;
wire n_805;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_996;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_1037;
wire n_1160;
wire n_202;
wire n_1080;
wire n_266;
wire n_1162;
wire n_491;
wire n_272;
wire n_1074;
wire n_427;
wire n_1199;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_1181;
wire n_1196;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_1186;
wire n_242;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_200;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_1184;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_1189;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_1180;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_1170;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_155),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_85),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_83),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_91),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_48),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_127),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_37),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_56),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_39),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_122),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_77),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_180),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_3),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_43),
.Y(n_201)
);

BUFx8_ASAP7_75t_SL g202 ( 
.A(n_154),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_78),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_87),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_72),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_134),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_151),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_125),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_84),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_156),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_44),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_97),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_166),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_161),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_8),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_30),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_53),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_38),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_39),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_176),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_139),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_59),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_66),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_179),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_64),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_120),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_60),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_171),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_94),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_50),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_22),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_20),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_61),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_7),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_65),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_162),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_167),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_71),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_33),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_147),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_11),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_70),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_136),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_28),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_131),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_111),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_19),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_144),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_133),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_26),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_31),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_110),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_50),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_115),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_1),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_44),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_108),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_29),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_76),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_29),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_9),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_132),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_82),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_146),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_141),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_170),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_90),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_163),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_67),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_57),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_68),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_175),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_40),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_160),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_177),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_173),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_45),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_23),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_14),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_153),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_116),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_6),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_62),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_31),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_13),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_103),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_26),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_164),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_0),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_52),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_168),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_129),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_75),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_30),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_52),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_165),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_225),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_200),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_219),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_221),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_234),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_235),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_247),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_0),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_249),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_273),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_281),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_196),
.B(n_1),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_195),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_201),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_196),
.B(n_204),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_202),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_220),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_204),
.B(n_2),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_213),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_236),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_243),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_222),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_223),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_238),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_214),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_255),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_205),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_245),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_262),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_248),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_251),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_206),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_254),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_2),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_291),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_257),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_190),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_260),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_207),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_208),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_190),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_264),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_214),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_209),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_184),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_299),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_189),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_210),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_285),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_215),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_241),
.B(n_3),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_299),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_217),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_191),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_198),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_265),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_224),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_211),
.Y(n_365)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_193),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_193),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_246),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_258),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_271),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_275),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_218),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_227),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_282),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_276),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_278),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_241),
.B(n_55),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_228),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_282),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_229),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_283),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_218),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_233),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_183),
.B(n_4),
.Y(n_384)
);

XOR2x2_ASAP7_75t_SL g385 ( 
.A(n_283),
.B(n_4),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_279),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_287),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_288),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_314),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_320),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_387),
.B(n_183),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_182),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_305),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_197),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_306),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_307),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_319),
.B(n_216),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_330),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_333),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_377),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_182),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_350),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_377),
.B(n_218),
.Y(n_407)
);

OA21x2_ASAP7_75t_L g408 ( 
.A1(n_388),
.A2(n_212),
.B(n_197),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_352),
.B(n_185),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_379),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_353),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_359),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_317),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_302),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_354),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_361),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_318),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_362),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_322),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_365),
.B(n_212),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_368),
.B(n_185),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_311),
.B(n_288),
.Y(n_425)
);

OA21x2_ASAP7_75t_L g426 ( 
.A1(n_369),
.A2(n_295),
.B(n_231),
.Y(n_426)
);

OA21x2_ASAP7_75t_L g427 ( 
.A1(n_370),
.A2(n_295),
.B(n_231),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

AND2x2_ASAP7_75t_SL g429 ( 
.A(n_315),
.B(n_296),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_348),
.A2(n_298),
.B1(n_294),
.B2(n_293),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_327),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_328),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_324),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_386),
.B(n_186),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_329),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_331),
.B(n_296),
.Y(n_438)
);

AND2x6_ASAP7_75t_L g439 ( 
.A(n_323),
.B(n_218),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_367),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_332),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_335),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_358),
.B(n_226),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_340),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_384),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_321),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_321),
.B(n_300),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_343),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_346),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_346),
.B(n_218),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_303),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_389),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_302),
.B(n_230),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_303),
.B(n_186),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_304),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_304),
.B(n_230),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_403),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_397),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_397),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_403),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_429),
.A2(n_230),
.B1(n_348),
.B2(n_366),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_403),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_230),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_403),
.B(n_230),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_403),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_403),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_429),
.A2(n_366),
.B1(n_277),
.B2(n_289),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_403),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_396),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_429),
.A2(n_298),
.B1(n_289),
.B2(n_293),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_397),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_395),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_395),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_396),
.B(n_232),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_430),
.A2(n_294),
.B1(n_381),
.B2(n_374),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_396),
.A2(n_374),
.B1(n_381),
.B2(n_188),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_446),
.A2(n_187),
.B1(n_188),
.B2(n_192),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_408),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_338),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_408),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_398),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_446),
.B(n_308),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_435),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_408),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_446),
.B(n_308),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_398),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_435),
.Y(n_494)
);

AND3x1_ASAP7_75t_L g495 ( 
.A(n_425),
.B(n_385),
.C(n_356),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_393),
.B(n_341),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_408),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_439),
.A2(n_297),
.B1(n_192),
.B2(n_194),
.Y(n_500)
);

CKINVDCx11_ASAP7_75t_R g501 ( 
.A(n_417),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_444),
.B(n_345),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_435),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_425),
.B(n_347),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_398),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_455),
.B(n_351),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_455),
.B(n_355),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_435),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_419),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_445),
.B(n_309),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_405),
.B(n_309),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_399),
.B(n_325),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_390),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_419),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_439),
.A2(n_407),
.B1(n_445),
.B2(n_392),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_405),
.B(n_357),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_457),
.B(n_385),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_419),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_430),
.A2(n_349),
.B1(n_334),
.B2(n_336),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_456),
.B(n_360),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_398),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_402),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_398),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_428),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_456),
.B(n_364),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_518),
.A2(n_407),
.B1(n_439),
.B2(n_392),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_518),
.A2(n_439),
.B1(n_392),
.B2(n_457),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_485),
.B(n_452),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_518),
.A2(n_439),
.B1(n_457),
.B2(n_445),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_462),
.B(n_453),
.C(n_449),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_489),
.B(n_452),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_509),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_462),
.B(n_452),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_471),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_471),
.B(n_516),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_471),
.B(n_457),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_471),
.B(n_457),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_509),
.B(n_450),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_516),
.B(n_454),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_502),
.B(n_470),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_478),
.B(n_454),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_461),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_492),
.B(n_447),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_466),
.B(n_467),
.Y(n_546)
);

BUFx4_ASAP7_75t_L g547 ( 
.A(n_495),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_470),
.B(n_373),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_492),
.B(n_434),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_466),
.B(n_447),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_466),
.B(n_447),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_518),
.A2(n_383),
.B1(n_378),
.B2(n_380),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_467),
.B(n_473),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_467),
.B(n_439),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_492),
.B(n_434),
.Y(n_555)
);

AOI221xp5_ASAP7_75t_L g556 ( 
.A1(n_495),
.A2(n_443),
.B1(n_410),
.B2(n_453),
.C(n_449),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_458),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_461),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_467),
.B(n_439),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_L g560 ( 
.A(n_483),
.B(n_334),
.C(n_326),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_463),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_467),
.B(n_434),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_511),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_467),
.B(n_394),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_475),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_467),
.B(n_394),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_523),
.Y(n_567)
);

NOR2xp67_ASAP7_75t_SL g568 ( 
.A(n_481),
.B(n_426),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_458),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_511),
.B(n_443),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_473),
.B(n_514),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_513),
.B(n_440),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_458),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_512),
.B(n_434),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_469),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_473),
.B(n_434),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_514),
.B(n_434),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_469),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_514),
.B(n_434),
.Y(n_579)
);

NOR3xp33_ASAP7_75t_L g580 ( 
.A(n_504),
.B(n_417),
.C(n_336),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_511),
.B(n_450),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_469),
.B(n_451),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_480),
.B(n_450),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_496),
.B(n_326),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_469),
.B(n_451),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_459),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_463),
.B(n_451),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_481),
.B(n_418),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_481),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_484),
.B(n_486),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_510),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_510),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_464),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_484),
.B(n_418),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_515),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_518),
.B(n_391),
.Y(n_596)
);

OAI221xp5_ASAP7_75t_L g597 ( 
.A1(n_468),
.A2(n_409),
.B1(n_424),
.B2(n_436),
.C(n_422),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_480),
.B(n_337),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_515),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_484),
.B(n_418),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_459),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_486),
.B(n_418),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_475),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_486),
.B(n_418),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_476),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_500),
.B(n_518),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_506),
.B(n_337),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_491),
.B(n_426),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_507),
.B(n_339),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_476),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_482),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_482),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_588),
.A2(n_497),
.B(n_491),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_536),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_594),
.A2(n_497),
.B(n_491),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_600),
.A2(n_497),
.B(n_465),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_590),
.A2(n_465),
.B(n_490),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_542),
.B(n_517),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_602),
.A2(n_604),
.B(n_546),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_536),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_598),
.B(n_479),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_538),
.A2(n_464),
.B(n_498),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_529),
.A2(n_483),
.B1(n_312),
.B2(n_301),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_589),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_539),
.A2(n_464),
.B(n_498),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_553),
.A2(n_464),
.B(n_498),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_568),
.A2(n_494),
.B(n_490),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_530),
.B(n_521),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_571),
.A2(n_522),
.B(n_505),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_589),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_589),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_589),
.B(n_527),
.Y(n_632)
);

AO21x1_ASAP7_75t_L g633 ( 
.A1(n_606),
.A2(n_499),
.B(n_494),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_589),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_531),
.B(n_499),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_543),
.B(n_518),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_567),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_545),
.B(n_518),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_557),
.Y(n_639)
);

AND2x4_ASAP7_75t_SL g640 ( 
.A(n_570),
.B(n_310),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_591),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_545),
.B(n_488),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_550),
.A2(n_525),
.B(n_508),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_551),
.A2(n_585),
.B(n_582),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_563),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_563),
.B(n_488),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_584),
.B(n_520),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_591),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_528),
.B(n_503),
.Y(n_649)
);

BUFx12f_ASAP7_75t_L g650 ( 
.A(n_567),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_537),
.B(n_503),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_606),
.A2(n_472),
.B(n_520),
.C(n_479),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_592),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_607),
.B(n_313),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_570),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_547),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_533),
.B(n_565),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_603),
.B(n_519),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_541),
.B(n_524),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_557),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_592),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_605),
.B(n_524),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_595),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_610),
.B(n_526),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_544),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_572),
.B(n_472),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_608),
.A2(n_526),
.B(n_525),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_611),
.B(n_448),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_612),
.B(n_581),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_548),
.B(n_501),
.C(n_342),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_535),
.B(n_448),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_583),
.A2(n_448),
.B(n_422),
.C(n_432),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_593),
.A2(n_426),
.B1(n_427),
.B2(n_342),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_595),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_547),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_544),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_554),
.A2(n_493),
.B(n_487),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_559),
.A2(n_577),
.B(n_576),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_596),
.B(n_493),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_579),
.A2(n_493),
.B(n_487),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_598),
.B(n_339),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_558),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_593),
.A2(n_426),
.B1(n_427),
.B2(n_363),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_L g684 ( 
.A(n_558),
.B(n_237),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_534),
.B(n_448),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_569),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_569),
.B(n_477),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_561),
.Y(n_688)
);

O2A1O1Ixp33_ASAP7_75t_SL g689 ( 
.A1(n_549),
.A2(n_474),
.B(n_460),
.C(n_420),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_573),
.B(n_477),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_587),
.A2(n_487),
.B(n_477),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_540),
.B(n_416),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_561),
.B(n_344),
.Y(n_693)
);

AOI21x1_ASAP7_75t_L g694 ( 
.A1(n_555),
.A2(n_474),
.B(n_460),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_562),
.A2(n_487),
.B(n_477),
.Y(n_695)
);

AOI21x1_ASAP7_75t_L g696 ( 
.A1(n_574),
.A2(n_427),
.B(n_426),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_573),
.A2(n_487),
.B(n_477),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_692),
.B(n_540),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_613),
.A2(n_566),
.B(n_564),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_628),
.B(n_609),
.Y(n_700)
);

AOI21x1_ASAP7_75t_L g701 ( 
.A1(n_679),
.A2(n_599),
.B(n_586),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_640),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_628),
.B(n_552),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_641),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_618),
.A2(n_597),
.B(n_566),
.C(n_564),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_615),
.A2(n_540),
.B(n_575),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_640),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_641),
.Y(n_708)
);

A2O1A1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_618),
.A2(n_652),
.B(n_666),
.C(n_647),
.Y(n_709)
);

NOR2x1_ASAP7_75t_L g710 ( 
.A(n_637),
.B(n_532),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_648),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_652),
.A2(n_540),
.B1(n_578),
.B2(n_560),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_655),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_619),
.A2(n_578),
.B(n_599),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_623),
.B(n_556),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_648),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_636),
.B(n_601),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_653),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_642),
.B(n_580),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_653),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_638),
.A2(n_349),
.B1(n_363),
.B2(n_187),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_661),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_632),
.A2(n_297),
.B1(n_199),
.B2(n_203),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_654),
.B(n_194),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_667),
.A2(n_427),
.B(n_477),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_661),
.B(n_423),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_663),
.B(n_423),
.Y(n_727)
);

O2A1O1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_681),
.A2(n_632),
.B(n_693),
.C(n_621),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_654),
.B(n_203),
.C(n_199),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_692),
.B(n_280),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_650),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_616),
.A2(n_477),
.B(n_427),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_650),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_SL g734 ( 
.A1(n_678),
.A2(n_420),
.B(n_431),
.C(n_433),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_663),
.B(n_423),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_634),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_634),
.A2(n_290),
.B1(n_280),
.B2(n_284),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_674),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_657),
.A2(n_423),
.B(n_438),
.C(n_431),
.Y(n_739)
);

O2A1O1Ixp5_ASAP7_75t_L g740 ( 
.A1(n_679),
.A2(n_423),
.B(n_438),
.C(n_433),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_646),
.A2(n_433),
.B(n_428),
.C(n_437),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_645),
.A2(n_442),
.B(n_441),
.C(n_437),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_656),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_674),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_644),
.A2(n_421),
.B(n_418),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_R g746 ( 
.A(n_614),
.B(n_284),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_692),
.B(n_290),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_665),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_676),
.B(n_438),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_634),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_649),
.A2(n_421),
.B(n_418),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_682),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_688),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_620),
.B(n_437),
.Y(n_754)
);

O2A1O1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_685),
.A2(n_684),
.B(n_672),
.C(n_669),
.Y(n_755)
);

AO32x2_ASAP7_75t_L g756 ( 
.A1(n_673),
.A2(n_438),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_675),
.B(n_292),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_634),
.B(n_438),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_649),
.A2(n_421),
.B(n_401),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_624),
.B(n_292),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_748),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_705),
.A2(n_625),
.B(n_622),
.Y(n_762)
);

OAI22x1_ASAP7_75t_L g763 ( 
.A1(n_703),
.A2(n_651),
.B1(n_659),
.B2(n_635),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_736),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_699),
.A2(n_635),
.B(n_671),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_752),
.Y(n_766)
);

AO31x2_ASAP7_75t_L g767 ( 
.A1(n_712),
.A2(n_633),
.A3(n_683),
.B(n_629),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_755),
.A2(n_626),
.B(n_691),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_713),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_708),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_753),
.Y(n_771)
);

AOI221x1_ASAP7_75t_L g772 ( 
.A1(n_709),
.A2(n_700),
.B1(n_724),
.B2(n_745),
.C(n_732),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_719),
.B(n_668),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_736),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_704),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_711),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_736),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_719),
.B(n_659),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_715),
.A2(n_651),
.B(n_664),
.C(n_662),
.Y(n_779)
);

OA21x2_ASAP7_75t_L g780 ( 
.A1(n_725),
.A2(n_617),
.B(n_643),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_716),
.Y(n_781)
);

OAI21x1_ASAP7_75t_SL g782 ( 
.A1(n_728),
.A2(n_627),
.B(n_694),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_714),
.A2(n_695),
.B(n_680),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_710),
.A2(n_670),
.B1(n_658),
.B2(n_660),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_718),
.Y(n_785)
);

AOI31xp67_ASAP7_75t_L g786 ( 
.A1(n_717),
.A2(n_744),
.A3(n_720),
.B(n_687),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_698),
.B(n_630),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_729),
.A2(n_630),
.B(n_631),
.C(n_677),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_721),
.A2(n_689),
.B(n_442),
.C(n_441),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_706),
.A2(n_631),
.B(n_697),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_717),
.A2(n_689),
.B(n_687),
.Y(n_791)
);

AO32x2_ASAP7_75t_L g792 ( 
.A1(n_723),
.A2(n_696),
.A3(n_690),
.B1(n_686),
.B2(n_660),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_701),
.A2(n_751),
.B(n_759),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_750),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_740),
.A2(n_690),
.B(n_686),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_722),
.B(n_639),
.Y(n_796)
);

AO31x2_ASAP7_75t_L g797 ( 
.A1(n_739),
.A2(n_441),
.A3(n_442),
.B(n_413),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_726),
.A2(n_639),
.B(n_268),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_741),
.A2(n_412),
.B(n_415),
.Y(n_799)
);

OAI21x1_ASAP7_75t_L g800 ( 
.A1(n_726),
.A2(n_412),
.B(n_415),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_738),
.B(n_404),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_754),
.B(n_727),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_727),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_754),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_733),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_750),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_750),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_702),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_757),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_769),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_786),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_761),
.Y(n_812)
);

CKINVDCx11_ASAP7_75t_R g813 ( 
.A(n_809),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_773),
.A2(n_707),
.B1(n_743),
.B2(n_731),
.Y(n_814)
);

INVx6_ASAP7_75t_L g815 ( 
.A(n_777),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_787),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_766),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_808),
.Y(n_818)
);

BUFx4_ASAP7_75t_SL g819 ( 
.A(n_805),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_784),
.A2(n_747),
.B1(n_730),
.B2(n_760),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_SL g821 ( 
.A1(n_809),
.A2(n_746),
.B1(n_756),
.B2(n_749),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_786),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_778),
.A2(n_737),
.B1(n_749),
.B2(n_735),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_805),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_771),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_806),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_806),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_802),
.A2(n_735),
.B1(n_758),
.B2(n_269),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_777),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_802),
.A2(n_266),
.B1(n_240),
.B2(n_242),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_809),
.A2(n_270),
.B1(n_244),
.B2(n_250),
.Y(n_831)
);

INVx4_ASAP7_75t_SL g832 ( 
.A(n_797),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_777),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_804),
.B(n_58),
.Y(n_834)
);

BUFx4_ASAP7_75t_SL g835 ( 
.A(n_808),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_763),
.A2(n_272),
.B1(n_252),
.B2(n_253),
.Y(n_836)
);

OAI22xp33_ASAP7_75t_L g837 ( 
.A1(n_772),
.A2(n_239),
.B1(n_256),
.B2(n_261),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_777),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_803),
.A2(n_263),
.B1(n_267),
.B2(n_421),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_775),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_774),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_798),
.A2(n_414),
.B1(n_413),
.B2(n_411),
.Y(n_842)
);

OAI22xp33_ASAP7_75t_L g843 ( 
.A1(n_776),
.A2(n_756),
.B1(n_414),
.B2(n_411),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_796),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_770),
.Y(n_845)
);

BUFx4_ASAP7_75t_SL g846 ( 
.A(n_781),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_770),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_779),
.A2(n_742),
.B1(n_756),
.B2(n_734),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_785),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_785),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_764),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_764),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_801),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_801),
.A2(n_406),
.B1(n_9),
.B2(n_10),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_764),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_794),
.Y(n_856)
);

BUFx4f_ASAP7_75t_SL g857 ( 
.A(n_794),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_779),
.A2(n_406),
.B1(n_10),
.B2(n_11),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_762),
.A2(n_796),
.B1(n_765),
.B2(n_782),
.Y(n_859)
);

BUFx8_ASAP7_75t_L g860 ( 
.A(n_774),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_794),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_807),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_807),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_799),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_792),
.Y(n_865)
);

AO21x1_ASAP7_75t_L g866 ( 
.A1(n_843),
.A2(n_768),
.B(n_783),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_865),
.B(n_792),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_858),
.A2(n_788),
.B(n_789),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_811),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_832),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_811),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_865),
.B(n_792),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_822),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_832),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_822),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_865),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_865),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_820),
.A2(n_791),
.B1(n_780),
.B2(n_790),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_832),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_865),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_832),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_859),
.B(n_767),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_864),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_849),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_816),
.Y(n_885)
);

AO21x2_ASAP7_75t_L g886 ( 
.A1(n_848),
.A2(n_793),
.B(n_800),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_860),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_SL g888 ( 
.A1(n_834),
.A2(n_780),
.B1(n_795),
.B2(n_800),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_821),
.B(n_792),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_849),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_845),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_840),
.B(n_792),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_845),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_854),
.A2(n_780),
.B1(n_799),
.B2(n_14),
.Y(n_894)
);

INVxp67_ASAP7_75t_SL g895 ( 
.A(n_812),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_816),
.Y(n_896)
);

BUFx2_ASAP7_75t_SL g897 ( 
.A(n_817),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_850),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_850),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_844),
.B(n_767),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_853),
.B(n_767),
.Y(n_901)
);

NOR2x1_ASAP7_75t_SL g902 ( 
.A(n_897),
.B(n_825),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_884),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_897),
.B(n_826),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_SL g905 ( 
.A1(n_868),
.A2(n_814),
.B(n_837),
.C(n_818),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_884),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_887),
.Y(n_907)
);

OAI211xp5_ASAP7_75t_L g908 ( 
.A1(n_868),
.A2(n_836),
.B(n_831),
.C(n_813),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_878),
.A2(n_830),
.B(n_828),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_885),
.B(n_896),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_895),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_885),
.B(n_826),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_896),
.B(n_810),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_885),
.B(n_810),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_874),
.B(n_852),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_878),
.A2(n_834),
.B(n_823),
.C(n_839),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_SL g917 ( 
.A1(n_901),
.A2(n_895),
.B(n_882),
.C(n_881),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_900),
.B(n_827),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_884),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_887),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_898),
.B(n_847),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_874),
.B(n_852),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_900),
.B(n_851),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_897),
.B(n_834),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_883),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_887),
.B(n_856),
.Y(n_926)
);

NOR2x1_ASAP7_75t_SL g927 ( 
.A(n_874),
.B(n_900),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_900),
.B(n_767),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_901),
.B(n_813),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_878),
.A2(n_842),
.B(n_862),
.C(n_856),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_874),
.B(n_829),
.Y(n_931)
);

AOI211xp5_ASAP7_75t_SL g932 ( 
.A1(n_889),
.A2(n_841),
.B(n_857),
.C(n_861),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_882),
.B(n_797),
.Y(n_933)
);

NOR3xp33_ASAP7_75t_SL g934 ( 
.A(n_879),
.B(n_824),
.C(n_862),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_894),
.A2(n_855),
.B(n_861),
.C(n_841),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_887),
.B(n_829),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_898),
.B(n_855),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_894),
.A2(n_824),
.B1(n_846),
.B2(n_815),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_890),
.B(n_829),
.Y(n_939)
);

OAI21x1_ASAP7_75t_SL g940 ( 
.A1(n_874),
.A2(n_863),
.B(n_835),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_874),
.B(n_829),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_925),
.B(n_867),
.Y(n_942)
);

NAND4xp25_ASAP7_75t_SL g943 ( 
.A(n_908),
.B(n_889),
.C(n_882),
.D(n_866),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_903),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_925),
.B(n_867),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_927),
.B(n_876),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_903),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_906),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_909),
.A2(n_889),
.B1(n_866),
.B2(n_886),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_906),
.B(n_876),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_928),
.B(n_867),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_938),
.A2(n_889),
.B1(n_866),
.B2(n_886),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_911),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_933),
.B(n_867),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_904),
.B(n_876),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_919),
.Y(n_956)
);

NOR2xp67_ASAP7_75t_L g957 ( 
.A(n_920),
.B(n_929),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_941),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_937),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_939),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_910),
.B(n_872),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_910),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_918),
.B(n_872),
.Y(n_963)
);

AO22x1_ASAP7_75t_L g964 ( 
.A1(n_907),
.A2(n_870),
.B1(n_881),
.B2(n_879),
.Y(n_964)
);

NAND4xp25_ASAP7_75t_L g965 ( 
.A(n_905),
.B(n_890),
.C(n_892),
.D(n_888),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_923),
.B(n_872),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_946),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_947),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_962),
.B(n_872),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_947),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_947),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_943),
.A2(n_929),
.B1(n_866),
.B2(n_924),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_947),
.Y(n_973)
);

INVx5_ASAP7_75t_L g974 ( 
.A(n_958),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_943),
.A2(n_916),
.B(n_905),
.Y(n_975)
);

AOI33xp33_ASAP7_75t_L g976 ( 
.A1(n_949),
.A2(n_935),
.A3(n_914),
.B1(n_912),
.B2(n_917),
.B3(n_892),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_959),
.B(n_892),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_942),
.B(n_880),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_959),
.B(n_892),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_948),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_948),
.Y(n_981)
);

CKINVDCx6p67_ASAP7_75t_R g982 ( 
.A(n_958),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_959),
.B(n_913),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_946),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_959),
.B(n_953),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_948),
.Y(n_986)
);

NOR2x1_ASAP7_75t_L g987 ( 
.A(n_965),
.B(n_904),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_985),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_983),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_967),
.B(n_962),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_967),
.B(n_960),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_984),
.B(n_960),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_985),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_970),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_977),
.B(n_979),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_977),
.B(n_979),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_968),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_974),
.B(n_946),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_989),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_995),
.B(n_983),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_995),
.B(n_982),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_988),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_996),
.B(n_982),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_988),
.B(n_976),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_990),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_996),
.B(n_982),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_L g1007 ( 
.A(n_1004),
.B(n_975),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_1005),
.B(n_990),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_999),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_1000),
.B(n_993),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1001),
.B(n_993),
.Y(n_1011)
);

OAI322xp33_ASAP7_75t_L g1012 ( 
.A1(n_1009),
.A2(n_1006),
.A3(n_1003),
.B1(n_1002),
.B2(n_997),
.C1(n_913),
.C2(n_994),
.Y(n_1012)
);

AOI311xp33_ASAP7_75t_L g1013 ( 
.A1(n_1007),
.A2(n_975),
.A3(n_997),
.B(n_916),
.C(n_986),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1007),
.B(n_991),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_1011),
.A2(n_987),
.B(n_972),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1008),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_1010),
.B(n_974),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1007),
.B(n_991),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1008),
.Y(n_1019)
);

OAI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_1009),
.A2(n_965),
.B1(n_987),
.B2(n_974),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1009),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_1009),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1008),
.B(n_998),
.Y(n_1023)
);

NAND4xp25_ASAP7_75t_L g1024 ( 
.A(n_1022),
.B(n_1021),
.C(n_1013),
.D(n_1015),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1019),
.B(n_998),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1019),
.B(n_992),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1016),
.B(n_992),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_1014),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_1018),
.A2(n_949),
.B(n_952),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_1012),
.B(n_998),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_1020),
.A2(n_930),
.B(n_952),
.C(n_932),
.Y(n_1031)
);

OAI21xp33_ASAP7_75t_L g1032 ( 
.A1(n_1023),
.A2(n_934),
.B(n_930),
.Y(n_1032)
);

NAND2x1p5_ASAP7_75t_L g1033 ( 
.A(n_1017),
.B(n_974),
.Y(n_1033)
);

OAI21xp33_ASAP7_75t_SL g1034 ( 
.A1(n_1017),
.A2(n_957),
.B(n_994),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1020),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1022),
.B(n_984),
.Y(n_1036)
);

OAI21xp33_ASAP7_75t_SL g1037 ( 
.A1(n_1017),
.A2(n_957),
.B(n_969),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_1019),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_SL g1039 ( 
.A1(n_1020),
.A2(n_819),
.B(n_5),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1025),
.B(n_974),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1038),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1026),
.Y(n_1042)
);

INVxp67_ASAP7_75t_SL g1043 ( 
.A(n_1024),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1027),
.Y(n_1044)
);

NAND3xp33_ASAP7_75t_L g1045 ( 
.A(n_1039),
.B(n_974),
.C(n_934),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1028),
.B(n_1035),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1036),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1029),
.A2(n_974),
.B1(n_958),
.B2(n_920),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1033),
.Y(n_1049)
);

AOI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_1034),
.A2(n_940),
.B(n_12),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1033),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1030),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1032),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1031),
.B(n_969),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1037),
.A2(n_958),
.B1(n_907),
.B2(n_924),
.Y(n_1055)
);

AOI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_1024),
.A2(n_917),
.B1(n_953),
.B2(n_980),
.C(n_968),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1028),
.B(n_978),
.Y(n_1057)
);

OAI31xp33_ASAP7_75t_L g1058 ( 
.A1(n_1029),
.A2(n_978),
.A3(n_946),
.B(n_936),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1047),
.B(n_978),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1052),
.B(n_970),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_SL g1061 ( 
.A(n_1050),
.B(n_958),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1041),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_L g1063 ( 
.A(n_1046),
.B(n_15),
.Y(n_1063)
);

NAND3xp33_ASAP7_75t_L g1064 ( 
.A(n_1043),
.B(n_1056),
.C(n_1053),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1043),
.B(n_970),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_SL g1066 ( 
.A(n_1042),
.B(n_15),
.C(n_16),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1044),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1040),
.Y(n_1068)
);

OAI321xp33_ASAP7_75t_L g1069 ( 
.A1(n_1055),
.A2(n_958),
.A3(n_924),
.B1(n_941),
.B2(n_931),
.C(n_904),
.Y(n_1069)
);

OAI21xp33_ASAP7_75t_L g1070 ( 
.A1(n_1054),
.A2(n_958),
.B(n_946),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_1045),
.B(n_958),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_L g1072 ( 
.A(n_1049),
.B(n_860),
.C(n_833),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_L g1073 ( 
.A(n_1051),
.B(n_973),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1057),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1048),
.B(n_973),
.Y(n_1075)
);

OA22x2_ASAP7_75t_L g1076 ( 
.A1(n_1071),
.A2(n_1055),
.B1(n_1058),
.B2(n_936),
.Y(n_1076)
);

OAI211xp5_ASAP7_75t_SL g1077 ( 
.A1(n_1064),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_1077)
);

AOI221xp5_ASAP7_75t_L g1078 ( 
.A1(n_1064),
.A2(n_980),
.B1(n_971),
.B2(n_986),
.C(n_964),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1061),
.A2(n_926),
.B1(n_960),
.B2(n_922),
.Y(n_1079)
);

OAI221xp5_ASAP7_75t_L g1080 ( 
.A1(n_1070),
.A2(n_941),
.B1(n_931),
.B2(n_971),
.C(n_981),
.Y(n_1080)
);

OAI221xp5_ASAP7_75t_SL g1081 ( 
.A1(n_1062),
.A2(n_1074),
.B1(n_1068),
.B2(n_1060),
.C(n_1067),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1063),
.A2(n_1073),
.B(n_1065),
.Y(n_1082)
);

AOI211xp5_ASAP7_75t_L g1083 ( 
.A1(n_1072),
.A2(n_964),
.B(n_18),
.C(n_19),
.Y(n_1083)
);

AOI222xp33_ASAP7_75t_L g1084 ( 
.A1(n_1059),
.A2(n_964),
.B1(n_902),
.B2(n_961),
.C1(n_22),
.C2(n_23),
.Y(n_1084)
);

AOI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_1066),
.A2(n_981),
.B1(n_973),
.B2(n_956),
.C(n_960),
.Y(n_1085)
);

OAI221xp5_ASAP7_75t_SL g1086 ( 
.A1(n_1075),
.A2(n_931),
.B1(n_961),
.B2(n_981),
.C(n_870),
.Y(n_1086)
);

NAND4xp25_ASAP7_75t_L g1087 ( 
.A(n_1069),
.B(n_926),
.C(n_915),
.D(n_922),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1063),
.B(n_961),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1061),
.A2(n_921),
.B(n_956),
.Y(n_1089)
);

OAI322xp33_ASAP7_75t_SL g1090 ( 
.A1(n_1062),
.A2(n_944),
.A3(n_948),
.B1(n_876),
.B2(n_877),
.C1(n_25),
.C2(n_27),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1061),
.A2(n_915),
.B1(n_922),
.B2(n_955),
.Y(n_1091)
);

AND2x2_ASAP7_75t_SL g1092 ( 
.A(n_1061),
.B(n_863),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_1063),
.Y(n_1093)
);

AOI321xp33_ASAP7_75t_L g1094 ( 
.A1(n_1071),
.A2(n_955),
.A3(n_20),
.B1(n_21),
.B2(n_24),
.C(n_25),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1061),
.A2(n_915),
.B(n_944),
.Y(n_1095)
);

O2A1O1Ixp5_ASAP7_75t_L g1096 ( 
.A1(n_1071),
.A2(n_955),
.B(n_863),
.C(n_939),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1064),
.A2(n_17),
.B(n_21),
.C(n_24),
.Y(n_1097)
);

AOI221xp5_ASAP7_75t_L g1098 ( 
.A1(n_1064),
.A2(n_955),
.B1(n_28),
.B2(n_32),
.C(n_33),
.Y(n_1098)
);

OAI211xp5_ASAP7_75t_L g1099 ( 
.A1(n_1064),
.A2(n_27),
.B(n_32),
.C(n_34),
.Y(n_1099)
);

OAI211xp5_ASAP7_75t_L g1100 ( 
.A1(n_1097),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_1100)
);

OAI211xp5_ASAP7_75t_L g1101 ( 
.A1(n_1099),
.A2(n_1098),
.B(n_1077),
.C(n_1094),
.Y(n_1101)
);

AOI31xp33_ASAP7_75t_L g1102 ( 
.A1(n_1093),
.A2(n_860),
.A3(n_36),
.B(n_37),
.Y(n_1102)
);

AOI222xp33_ASAP7_75t_L g1103 ( 
.A1(n_1078),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.C1(n_41),
.C2(n_42),
.Y(n_1103)
);

NOR4xp25_ASAP7_75t_L g1104 ( 
.A(n_1081),
.B(n_41),
.C(n_42),
.D(n_43),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_SL g1105 ( 
.A(n_1082),
.B(n_815),
.Y(n_1105)
);

AOI221x1_ASAP7_75t_L g1106 ( 
.A1(n_1087),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.C(n_48),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1076),
.A2(n_870),
.B1(n_955),
.B2(n_881),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1088),
.Y(n_1108)
);

AO22x2_ASAP7_75t_L g1109 ( 
.A1(n_1090),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_1109)
);

AOI221xp5_ASAP7_75t_L g1110 ( 
.A1(n_1083),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.C(n_54),
.Y(n_1110)
);

AOI211xp5_ASAP7_75t_L g1111 ( 
.A1(n_1086),
.A2(n_51),
.B(n_54),
.C(n_829),
.Y(n_1111)
);

AOI211xp5_ASAP7_75t_L g1112 ( 
.A1(n_1085),
.A2(n_1080),
.B(n_1079),
.C(n_1095),
.Y(n_1112)
);

AOI221xp5_ASAP7_75t_L g1113 ( 
.A1(n_1096),
.A2(n_950),
.B1(n_880),
.B2(n_833),
.C(n_838),
.Y(n_1113)
);

OAI211xp5_ASAP7_75t_L g1114 ( 
.A1(n_1084),
.A2(n_833),
.B(n_838),
.C(n_888),
.Y(n_1114)
);

OAI211xp5_ASAP7_75t_SL g1115 ( 
.A1(n_1091),
.A2(n_855),
.B(n_861),
.C(n_879),
.Y(n_1115)
);

AOI211xp5_ASAP7_75t_L g1116 ( 
.A1(n_1089),
.A2(n_833),
.B(n_838),
.C(n_954),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_SL g1117 ( 
.A1(n_1092),
.A2(n_815),
.B1(n_954),
.B2(n_833),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1093),
.Y(n_1118)
);

AOI321xp33_ASAP7_75t_L g1119 ( 
.A1(n_1081),
.A2(n_954),
.A3(n_951),
.B1(n_945),
.B2(n_942),
.C(n_963),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1093),
.B(n_963),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1093),
.Y(n_1121)
);

AOI211xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1081),
.A2(n_951),
.B(n_945),
.C(n_942),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1077),
.A2(n_815),
.B1(n_951),
.B2(n_950),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1118),
.B(n_63),
.Y(n_1124)
);

OAI221xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1104),
.A2(n_1107),
.B1(n_1121),
.B2(n_1111),
.C(n_1101),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1108),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_1102),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1120),
.A2(n_1109),
.B1(n_1110),
.B2(n_1114),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1100),
.B(n_963),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1109),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1106),
.Y(n_1131)
);

BUFx4f_ASAP7_75t_SL g1132 ( 
.A(n_1105),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1123),
.B(n_966),
.Y(n_1133)
);

AND2x2_ASAP7_75t_SL g1134 ( 
.A(n_1113),
.B(n_838),
.Y(n_1134)
);

INVxp33_ASAP7_75t_L g1135 ( 
.A(n_1117),
.Y(n_1135)
);

INVxp67_ASAP7_75t_SL g1136 ( 
.A(n_1103),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1115),
.B(n_69),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_1122),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1112),
.Y(n_1139)
);

HB1xp67_ASAP7_75t_L g1140 ( 
.A(n_1116),
.Y(n_1140)
);

NOR2x1_ASAP7_75t_L g1141 ( 
.A(n_1119),
.B(n_838),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_1118),
.Y(n_1142)
);

NAND4xp75_ASAP7_75t_L g1143 ( 
.A(n_1121),
.B(n_945),
.C(n_966),
.D(n_890),
.Y(n_1143)
);

AO22x2_ASAP7_75t_L g1144 ( 
.A1(n_1121),
.A2(n_950),
.B1(n_877),
.B2(n_966),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1118),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1131),
.B(n_950),
.Y(n_1146)
);

AND2x2_ASAP7_75t_SL g1147 ( 
.A(n_1145),
.B(n_950),
.Y(n_1147)
);

AND4x2_ASAP7_75t_L g1148 ( 
.A(n_1141),
.B(n_73),
.C(n_74),
.D(n_79),
.Y(n_1148)
);

AOI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1130),
.A2(n_880),
.B1(n_898),
.B2(n_899),
.C(n_883),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1138),
.A2(n_877),
.B1(n_880),
.B2(n_886),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1142),
.B(n_883),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1139),
.A2(n_80),
.B(n_81),
.C(n_86),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1127),
.A2(n_880),
.B1(n_877),
.B2(n_871),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_1126),
.B(n_88),
.Y(n_1154)
);

AOI32xp33_ASAP7_75t_L g1155 ( 
.A1(n_1135),
.A2(n_1136),
.A3(n_1129),
.B1(n_1140),
.B2(n_1124),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1125),
.A2(n_89),
.B(n_92),
.C(n_93),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1128),
.B(n_886),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1143),
.Y(n_1158)
);

OAI211xp5_ASAP7_75t_L g1159 ( 
.A1(n_1137),
.A2(n_95),
.B(n_96),
.C(n_98),
.Y(n_1159)
);

NAND4xp75_ASAP7_75t_L g1160 ( 
.A(n_1134),
.B(n_99),
.C(n_100),
.D(n_101),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1154),
.Y(n_1161)
);

O2A1O1Ixp5_ASAP7_75t_SL g1162 ( 
.A1(n_1159),
.A2(n_1132),
.B(n_1144),
.C(n_1133),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1158),
.A2(n_1133),
.B1(n_1144),
.B2(n_880),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1146),
.B(n_102),
.Y(n_1164)
);

AOI221xp5_ASAP7_75t_L g1165 ( 
.A1(n_1156),
.A2(n_880),
.B1(n_899),
.B2(n_883),
.C(n_869),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1147),
.Y(n_1166)
);

XOR2xp5_ASAP7_75t_L g1167 ( 
.A(n_1160),
.B(n_104),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1151),
.Y(n_1168)
);

OAI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1155),
.A2(n_899),
.B1(n_880),
.B2(n_883),
.C(n_891),
.Y(n_1169)
);

XNOR2x1_ASAP7_75t_L g1170 ( 
.A(n_1157),
.B(n_105),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1150),
.B(n_1153),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1152),
.B(n_883),
.Y(n_1172)
);

AND2x2_ASAP7_75t_SL g1173 ( 
.A(n_1148),
.B(n_106),
.Y(n_1173)
);

AND2x2_ASAP7_75t_SL g1174 ( 
.A(n_1149),
.B(n_107),
.Y(n_1174)
);

XOR2xp5_ASAP7_75t_L g1175 ( 
.A(n_1146),
.B(n_113),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1173),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1161),
.Y(n_1177)
);

AOI22x1_ASAP7_75t_SL g1178 ( 
.A1(n_1166),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1175),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1174),
.A2(n_880),
.B1(n_886),
.B2(n_869),
.Y(n_1180)
);

OAI22x1_ASAP7_75t_L g1181 ( 
.A1(n_1167),
.A2(n_871),
.B1(n_869),
.B2(n_875),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1164),
.Y(n_1182)
);

OAI22xp33_ASAP7_75t_SL g1183 ( 
.A1(n_1163),
.A2(n_871),
.B1(n_891),
.B2(n_893),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1170),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1168),
.A2(n_886),
.B1(n_875),
.B2(n_873),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1176),
.A2(n_1169),
.B1(n_1172),
.B2(n_1165),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1177),
.B(n_1162),
.Y(n_1187)
);

INVxp67_ASAP7_75t_SL g1188 ( 
.A(n_1184),
.Y(n_1188)
);

NOR3xp33_ASAP7_75t_L g1189 ( 
.A(n_1179),
.B(n_1171),
.C(n_121),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1180),
.A2(n_875),
.B1(n_873),
.B2(n_893),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1178),
.Y(n_1191)
);

OAI22xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1187),
.A2(n_1182),
.B1(n_1181),
.B2(n_1183),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1191),
.A2(n_1185),
.B1(n_123),
.B2(n_124),
.Y(n_1193)
);

OAI22x1_ASAP7_75t_L g1194 ( 
.A1(n_1188),
.A2(n_1185),
.B1(n_126),
.B2(n_128),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1186),
.A2(n_875),
.B1(n_873),
.B2(n_893),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1193),
.A2(n_1189),
.B1(n_1190),
.B2(n_873),
.Y(n_1196)
);

AOI221xp5_ASAP7_75t_L g1197 ( 
.A1(n_1196),
.A2(n_1192),
.B1(n_1194),
.B2(n_1195),
.C(n_137),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_SL g1198 ( 
.A1(n_1197),
.A2(n_119),
.B(n_130),
.Y(n_1198)
);

OAI31xp33_ASAP7_75t_L g1199 ( 
.A1(n_1198),
.A2(n_135),
.A3(n_138),
.B(n_140),
.Y(n_1199)
);

OAI221xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1199),
.A2(n_142),
.B1(n_143),
.B2(n_148),
.C(n_149),
.Y(n_1200)
);

AOI211xp5_ASAP7_75t_L g1201 ( 
.A1(n_1200),
.A2(n_150),
.B(n_152),
.C(n_158),
.Y(n_1201)
);


endmodule