module fake_jpeg_14909_n_180 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_7),
.B(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_37),
.Y(n_43)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_27),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_48),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_23),
.B1(n_19),
.B2(n_22),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_46),
.B1(n_38),
.B2(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_19),
.B1(n_28),
.B2(n_15),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_24),
.C(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_21),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_57),
.B(n_61),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_66),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_73),
.Y(n_76)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_36),
.B1(n_38),
.B2(n_19),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_47),
.B1(n_30),
.B2(n_33),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_16),
.B1(n_28),
.B2(n_15),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_18),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_38),
.A3(n_26),
.B1(n_33),
.B2(n_30),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_14),
.B(n_21),
.C(n_26),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_71),
.B1(n_14),
.B2(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_52),
.B1(n_45),
.B2(n_38),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_24),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_70),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_44),
.C(n_34),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_59),
.C(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_70),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_66),
.B1(n_50),
.B2(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_85),
.B1(n_88),
.B2(n_92),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_72),
.B1(n_55),
.B2(n_43),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_51),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_56),
.B(n_51),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_35),
.B1(n_32),
.B2(n_33),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_60),
.B1(n_32),
.B2(n_63),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_97),
.C(n_110),
.Y(n_115)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_104),
.Y(n_118)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_106),
.B1(n_93),
.B2(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_109),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_60),
.B1(n_22),
.B2(n_18),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_60),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_2),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_91),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_104),
.A3(n_95),
.B1(n_111),
.B2(n_97),
.C1(n_100),
.C2(n_109),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_120),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_83),
.B1(n_98),
.B2(n_80),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_121),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_90),
.C(n_77),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_128),
.C(n_105),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_91),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_88),
.B1(n_92),
.B2(n_85),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_84),
.B1(n_112),
.B2(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_102),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_90),
.C(n_87),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_138),
.C(n_139),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_116),
.B1(n_114),
.B2(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_107),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_127),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_134),
.B(n_137),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_117),
.B1(n_125),
.B2(n_126),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_119),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_12),
.C(n_11),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_127),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_144),
.B(n_150),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_122),
.C(n_125),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_136),
.C(n_135),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_126),
.B1(n_4),
.B2(n_5),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_130),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_153),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_141),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_152),
.C(n_153),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_139),
.C(n_131),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_147),
.C(n_142),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_129),
.B1(n_12),
.B2(n_6),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_4),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_3),
.B(n_4),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_146),
.B1(n_150),
.B2(n_142),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_148),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_166),
.B(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_148),
.Y(n_168)
);

OAI21x1_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_170),
.B(n_165),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_171),
.A2(n_165),
.B(n_8),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_7),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_176),
.B(n_174),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_9),
.B(n_10),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_9),
.Y(n_180)
);


endmodule