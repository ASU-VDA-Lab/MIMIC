module real_aes_2400_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_0), .B(n_154), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_1), .A2(n_163), .B(n_168), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_2), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_3), .B(n_154), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_4), .B(n_170), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_5), .B(n_170), .Y(n_208) );
INVx1_ASAP7_75t_L g161 ( .A(n_6), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_7), .B(n_170), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_8), .Y(n_110) );
NAND2xp33_ASAP7_75t_L g197 ( .A(n_9), .B(n_172), .Y(n_197) );
AND2x2_ASAP7_75t_L g507 ( .A(n_10), .B(n_191), .Y(n_507) );
AND2x2_ASAP7_75t_L g515 ( .A(n_11), .B(n_148), .Y(n_515) );
INVx2_ASAP7_75t_L g151 ( .A(n_12), .Y(n_151) );
AOI221x1_ASAP7_75t_L g243 ( .A1(n_13), .A2(n_24), .B1(n_154), .B2(n_163), .C(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_14), .B(n_170), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_15), .B(n_109), .C(n_111), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_15), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_16), .B(n_154), .Y(n_193) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_17), .A2(n_191), .B(n_192), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_18), .B(n_174), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_19), .B(n_170), .Y(n_184) );
AO21x1_ASAP7_75t_L g203 ( .A1(n_20), .A2(n_154), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_21), .B(n_154), .Y(n_488) );
NOR2xp33_ASAP7_75t_SL g105 ( .A(n_22), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g128 ( .A(n_22), .Y(n_128) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_23), .A2(n_90), .B1(n_154), .B2(n_523), .Y(n_522) );
NAND2x1_ASAP7_75t_L g216 ( .A(n_25), .B(n_170), .Y(n_216) );
NAND2x1_ASAP7_75t_L g235 ( .A(n_26), .B(n_172), .Y(n_235) );
OAI22xp5_ASAP7_75t_SL g783 ( .A1(n_27), .A2(n_62), .B1(n_784), .B2(n_785), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_27), .Y(n_784) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_28), .A2(n_87), .B(n_151), .Y(n_150) );
OR2x2_ASAP7_75t_L g176 ( .A(n_28), .B(n_87), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_29), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_30), .B(n_170), .Y(n_196) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_31), .A2(n_148), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_32), .B(n_172), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_33), .A2(n_163), .B(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_34), .B(n_170), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_35), .A2(n_163), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g160 ( .A(n_36), .B(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g164 ( .A(n_36), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g531 ( .A(n_36), .Y(n_531) );
INVxp67_ASAP7_75t_L g111 ( .A(n_37), .Y(n_111) );
OR2x6_ASAP7_75t_L g126 ( .A(n_37), .B(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_38), .B(n_154), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_39), .B(n_154), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_40), .B(n_170), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_41), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_42), .B(n_172), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_43), .B(n_154), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_44), .A2(n_163), .B(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_45), .A2(n_163), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_46), .B(n_172), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_47), .A2(n_51), .B1(n_132), .B2(n_133), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_47), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_48), .B(n_172), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_49), .B(n_154), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_50), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_51), .Y(n_132) );
INVx1_ASAP7_75t_L g157 ( .A(n_52), .Y(n_157) );
INVx1_ASAP7_75t_L g167 ( .A(n_52), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_53), .B(n_170), .Y(n_513) );
AND2x2_ASAP7_75t_L g479 ( .A(n_54), .B(n_174), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_55), .B(n_172), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_56), .B(n_170), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_57), .B(n_172), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_58), .A2(n_163), .B(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_59), .B(n_154), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_60), .B(n_154), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_61), .A2(n_163), .B(n_472), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_62), .Y(n_785) );
AO21x1_ASAP7_75t_L g205 ( .A1(n_63), .A2(n_163), .B(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g494 ( .A(n_64), .B(n_175), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_65), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_66), .B(n_172), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_67), .B(n_154), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_68), .B(n_172), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_69), .A2(n_95), .B1(n_163), .B2(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g228 ( .A(n_70), .B(n_175), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_71), .B(n_170), .Y(n_491) );
INVx1_ASAP7_75t_L g159 ( .A(n_72), .Y(n_159) );
INVx1_ASAP7_75t_L g165 ( .A(n_72), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_73), .Y(n_790) );
AND2x2_ASAP7_75t_L g239 ( .A(n_74), .B(n_148), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_75), .B(n_172), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_76), .A2(n_163), .B(n_483), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_77), .A2(n_163), .B(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_78), .A2(n_163), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g476 ( .A(n_79), .B(n_175), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_80), .B(n_174), .Y(n_520) );
INVx1_ASAP7_75t_L g106 ( .A(n_81), .Y(n_106) );
AND2x2_ASAP7_75t_L g147 ( .A(n_82), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_83), .B(n_154), .Y(n_186) );
AND2x2_ASAP7_75t_L g555 ( .A(n_84), .B(n_191), .Y(n_555) );
AND2x2_ASAP7_75t_L g204 ( .A(n_85), .B(n_180), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_86), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_88), .B(n_172), .Y(n_185) );
AND2x2_ASAP7_75t_L g220 ( .A(n_89), .B(n_148), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_91), .B(n_170), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_92), .A2(n_163), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_93), .B(n_172), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_94), .A2(n_163), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_96), .B(n_170), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_97), .B(n_170), .Y(n_169) );
BUFx2_ASAP7_75t_L g493 ( .A(n_98), .Y(n_493) );
BUFx2_ASAP7_75t_L g116 ( .A(n_99), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_100), .A2(n_163), .B(n_195), .Y(n_194) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_112), .B(n_789), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx3_ASAP7_75t_SL g791 ( .A(n_103), .Y(n_791) );
OR2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_107), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_106), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_130), .B(n_778), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_116), .Y(n_779) );
INVxp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_118), .A2(n_781), .B(n_786), .Y(n_780) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_129), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g788 ( .A(n_123), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
OR2x6_ASAP7_75t_SL g138 ( .A(n_124), .B(n_125), .Y(n_138) );
AND2x6_ASAP7_75t_SL g768 ( .A(n_124), .B(n_126), .Y(n_768) );
OR2x2_ASAP7_75t_L g777 ( .A(n_124), .B(n_126), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
OAI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_134), .B(n_769), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_131), .A2(n_770), .B(n_774), .Y(n_769) );
INVxp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_139), .B1(n_456), .B2(n_765), .Y(n_135) );
INVx1_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g773 ( .A(n_137), .Y(n_773) );
CKINVDCx11_ASAP7_75t_R g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g772 ( .A(n_139), .Y(n_772) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_365), .Y(n_139) );
NOR4xp25_ASAP7_75t_L g140 ( .A(n_141), .B(n_283), .C(n_309), .D(n_349), .Y(n_140) );
OAI211xp5_ASAP7_75t_SL g141 ( .A1(n_142), .A2(n_198), .B(n_229), .C(n_269), .Y(n_141) );
INVxp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_177), .Y(n_143) );
AND2x2_ASAP7_75t_L g436 ( .A(n_144), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_145), .B(n_177), .Y(n_303) );
BUFx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g230 ( .A(n_146), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_146), .B(n_256), .Y(n_255) );
INVx5_ASAP7_75t_L g289 ( .A(n_146), .Y(n_289) );
NOR2x1_ASAP7_75t_SL g331 ( .A(n_146), .B(n_178), .Y(n_331) );
AND2x2_ASAP7_75t_L g387 ( .A(n_146), .B(n_190), .Y(n_387) );
OR2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_152), .Y(n_146) );
INVx3_ASAP7_75t_L g219 ( .A(n_148), .Y(n_219) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_149), .A2(n_509), .B(n_515), .Y(n_508) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_150), .Y(n_191) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_151), .B(n_176), .Y(n_175) );
AND2x4_ASAP7_75t_L g180 ( .A(n_151), .B(n_176), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_162), .B(n_174), .Y(n_152) );
AND2x4_ASAP7_75t_L g154 ( .A(n_155), .B(n_160), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_158), .Y(n_155) );
AND2x6_ASAP7_75t_L g172 ( .A(n_156), .B(n_165), .Y(n_172) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g170 ( .A(n_158), .B(n_167), .Y(n_170) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx5_ASAP7_75t_L g173 ( .A(n_160), .Y(n_173) );
AND2x2_ASAP7_75t_L g166 ( .A(n_161), .B(n_167), .Y(n_166) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_161), .Y(n_526) );
AND2x6_ASAP7_75t_L g163 ( .A(n_164), .B(n_166), .Y(n_163) );
BUFx3_ASAP7_75t_L g527 ( .A(n_164), .Y(n_527) );
INVx2_ASAP7_75t_L g533 ( .A(n_165), .Y(n_533) );
AND2x4_ASAP7_75t_L g529 ( .A(n_166), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g525 ( .A(n_167), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_171), .B(n_173), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_172), .B(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_173), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_173), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_173), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_173), .A2(n_216), .B(n_217), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_173), .A2(n_225), .B(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_173), .A2(n_235), .B(n_236), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_173), .A2(n_245), .B(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_173), .A2(n_467), .B(n_468), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_173), .A2(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_173), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_173), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_173), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_173), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_173), .A2(n_553), .B(n_554), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_174), .Y(n_238) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_174), .A2(n_243), .B(n_247), .Y(n_242) );
OA21x2_ASAP7_75t_L g282 ( .A1(n_174), .A2(n_243), .B(n_247), .Y(n_282) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_174), .A2(n_522), .B(n_528), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_174), .A2(n_550), .B(n_551), .Y(n_549) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_189), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_178), .B(n_190), .Y(n_259) );
AND2x2_ASAP7_75t_L g320 ( .A(n_178), .B(n_289), .Y(n_320) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_181), .B(n_187), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_179), .B(n_188), .Y(n_187) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_179), .A2(n_181), .B(n_187), .Y(n_273) );
INVx1_ASAP7_75t_SL g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_180), .A2(n_193), .B(n_194), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_180), .B(n_210), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_180), .A2(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_180), .A2(n_481), .B(n_482), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_186), .Y(n_181) );
AND2x2_ASAP7_75t_L g332 ( .A(n_189), .B(n_256), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_189), .B(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g376 ( .A(n_189), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g409 ( .A(n_189), .B(n_230), .Y(n_409) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g253 ( .A(n_190), .Y(n_253) );
AND2x2_ASAP7_75t_L g286 ( .A(n_190), .B(n_287), .Y(n_286) );
BUFx3_ASAP7_75t_L g321 ( .A(n_190), .Y(n_321) );
OR2x2_ASAP7_75t_L g397 ( .A(n_190), .B(n_256), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_191), .A2(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_211), .Y(n_199) );
AOI211x1_ASAP7_75t_SL g326 ( .A1(n_200), .A2(n_318), .B(n_327), .C(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_200), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_200), .B(n_369), .Y(n_416) );
BUFx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g266 ( .A(n_201), .Y(n_266) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g241 ( .A(n_202), .Y(n_241) );
OAI21x1_ASAP7_75t_SL g202 ( .A1(n_203), .A2(n_205), .B(n_209), .Y(n_202) );
INVx1_ASAP7_75t_L g210 ( .A(n_204), .Y(n_210) );
AOI322xp5_ASAP7_75t_L g229 ( .A1(n_211), .A2(n_230), .A3(n_240), .B1(n_248), .B2(n_251), .C1(n_257), .C2(n_260), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_211), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_221), .Y(n_211) );
INVx2_ASAP7_75t_L g264 ( .A(n_212), .Y(n_264) );
INVxp67_ASAP7_75t_L g306 ( .A(n_212), .Y(n_306) );
BUFx3_ASAP7_75t_L g370 ( .A(n_212), .Y(n_370) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_219), .B(n_220), .Y(n_212) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_213), .A2(n_219), .B(n_220), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_218), .Y(n_213) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_219), .A2(n_222), .B(n_228), .Y(n_221) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_219), .A2(n_222), .B(n_228), .Y(n_268) );
AO21x1_ASAP7_75t_SL g469 ( .A1(n_219), .A2(n_470), .B(n_476), .Y(n_469) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_219), .A2(n_470), .B(n_476), .Y(n_545) );
INVx2_ASAP7_75t_L g279 ( .A(n_221), .Y(n_279) );
AND2x2_ASAP7_75t_L g328 ( .A(n_221), .B(n_242), .Y(n_328) );
AND2x2_ASAP7_75t_L g372 ( .A(n_221), .B(n_281), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_223), .B(n_227), .Y(n_222) );
AND2x2_ASAP7_75t_L g257 ( .A(n_230), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_230), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_230), .B(n_286), .Y(n_451) );
INVx4_ASAP7_75t_L g256 ( .A(n_231), .Y(n_256) );
AND2x2_ASAP7_75t_L g288 ( .A(n_231), .B(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_231), .Y(n_341) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_238), .B(n_239), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_237), .Y(n_232) );
AOI21x1_ASAP7_75t_L g500 ( .A1(n_238), .A2(n_501), .B(n_507), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_240), .B(n_325), .Y(n_350) );
INVx1_ASAP7_75t_SL g389 ( .A(n_240), .Y(n_389) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
AND2x4_ASAP7_75t_L g280 ( .A(n_241), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_241), .B(n_279), .Y(n_348) );
AND2x2_ASAP7_75t_L g400 ( .A(n_241), .B(n_250), .Y(n_400) );
OR2x2_ASAP7_75t_L g424 ( .A(n_241), .B(n_242), .Y(n_424) );
AND2x2_ASAP7_75t_L g248 ( .A(n_242), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g298 ( .A(n_242), .B(n_279), .Y(n_298) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_242), .B(n_266), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_248), .B(n_361), .Y(n_378) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
BUFx2_ASAP7_75t_L g313 ( .A(n_250), .Y(n_313) );
AND2x4_ASAP7_75t_SL g353 ( .A(n_250), .B(n_267), .Y(n_353) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
OR2x2_ASAP7_75t_L g301 ( .A(n_252), .B(n_255), .Y(n_301) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g270 ( .A(n_253), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g418 ( .A(n_253), .B(n_331), .Y(n_418) );
AND2x2_ASAP7_75t_L g434 ( .A(n_253), .B(n_288), .Y(n_434) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AOI311xp33_ASAP7_75t_L g404 ( .A1(n_255), .A2(n_343), .A3(n_405), .B(n_407), .C(n_414), .Y(n_404) );
AND2x4_ASAP7_75t_L g271 ( .A(n_256), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g275 ( .A(n_256), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_256), .B(n_289), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_256), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g388 ( .A(n_256), .B(n_375), .Y(n_388) );
AND2x2_ASAP7_75t_L g274 ( .A(n_258), .B(n_275), .Y(n_274) );
INVxp67_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_259), .Y(n_292) );
OR2x2_ASAP7_75t_L g381 ( .A(n_259), .B(n_345), .Y(n_381) );
INVx1_ASAP7_75t_L g437 ( .A(n_259), .Y(n_437) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g346 ( .A(n_263), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g360 ( .A(n_263), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g435 ( .A(n_263), .B(n_308), .Y(n_435) );
BUFx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g278 ( .A(n_264), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g297 ( .A(n_264), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g359 ( .A(n_265), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_265), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_414) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AND2x2_ASAP7_75t_L g308 ( .A(n_266), .B(n_279), .Y(n_308) );
AND2x4_ASAP7_75t_L g361 ( .A(n_266), .B(n_268), .Y(n_361) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI21xp33_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_274), .B(n_276), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_270), .A2(n_356), .B1(n_360), .B2(n_362), .Y(n_355) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_271), .B(n_289), .Y(n_315) );
INVx2_ASAP7_75t_L g377 ( .A(n_271), .Y(n_377) );
AND2x2_ASAP7_75t_L g391 ( .A(n_271), .B(n_387), .Y(n_391) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g287 ( .A(n_273), .Y(n_287) );
INVx1_ASAP7_75t_L g340 ( .A(n_273), .Y(n_340) );
INVx1_ASAP7_75t_L g291 ( .A(n_275), .Y(n_291) );
AND3x2_ASAP7_75t_L g319 ( .A(n_275), .B(n_320), .C(n_321), .Y(n_319) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx1_ASAP7_75t_L g383 ( .A(n_278), .Y(n_383) );
AND2x2_ASAP7_75t_L g311 ( .A(n_280), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g382 ( .A(n_280), .B(n_383), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_280), .A2(n_394), .B1(n_398), .B2(n_401), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_280), .B(n_428), .Y(n_432) );
BUFx2_ASAP7_75t_L g323 ( .A(n_281), .Y(n_323) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g294 ( .A(n_282), .Y(n_294) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_282), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_293), .B1(n_295), .B2(n_296), .C(n_299), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_290), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g375 ( .A(n_287), .Y(n_375) );
INVx2_ASAP7_75t_SL g364 ( .A(n_288), .Y(n_364) );
AND2x2_ASAP7_75t_L g446 ( .A(n_288), .B(n_313), .Y(n_446) );
INVx4_ASAP7_75t_L g337 ( .A(n_289), .Y(n_337) );
INVx1_ASAP7_75t_L g295 ( .A(n_290), .Y(n_295) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x4_ASAP7_75t_L g406 ( .A(n_294), .B(n_361), .Y(n_406) );
INVx1_ASAP7_75t_SL g445 ( .A(n_294), .Y(n_445) );
AND2x2_ASAP7_75t_L g450 ( .A(n_294), .B(n_353), .Y(n_450) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g392 ( .A(n_298), .Y(n_392) );
OAI21xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .B(n_304), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g325 ( .A(n_306), .Y(n_325) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g322 ( .A(n_308), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g412 ( .A(n_308), .B(n_413), .Y(n_412) );
OAI211xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_314), .B(n_316), .C(n_333), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g405 ( .A(n_312), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_313), .B(n_328), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_313), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g438 ( .A(n_313), .B(n_361), .Y(n_438) );
OAI221xp5_ASAP7_75t_SL g349 ( .A1(n_314), .A2(n_338), .B1(n_350), .B2(n_351), .C(n_355), .Y(n_349) );
INVx3_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g420 ( .A(n_315), .B(n_321), .Y(n_420) );
OAI32xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_322), .A3(n_324), .B1(n_326), .B2(n_330), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVxp67_ASAP7_75t_SL g410 ( .A(n_320), .Y(n_410) );
INVx2_ASAP7_75t_L g343 ( .A(n_321), .Y(n_343) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_321), .A2(n_373), .B(n_453), .C(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g358 ( .A(n_323), .Y(n_358) );
OR2x2_ASAP7_75t_L g454 ( .A(n_323), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_327), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g415 ( .A(n_330), .Y(n_415) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g396 ( .A(n_331), .Y(n_396) );
OAI21xp33_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_342), .B(n_346), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
OR2x2_ASAP7_75t_L g373 ( .A(n_336), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_337), .B(n_340), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_339), .A2(n_371), .B1(n_440), .B2(n_443), .C(n_447), .Y(n_439) );
INVx2_ASAP7_75t_L g442 ( .A(n_339), .Y(n_442) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
OR2x2_ASAP7_75t_L g363 ( .A(n_343), .B(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g430 ( .A(n_343), .B(n_388), .Y(n_430) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g428 ( .A(n_353), .Y(n_428) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_361), .B(n_391), .Y(n_448) );
INVx2_ASAP7_75t_L g455 ( .A(n_361), .Y(n_455) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_363), .A2(n_426), .B1(n_429), .B2(n_431), .C(n_433), .Y(n_425) );
AND5x1_ASAP7_75t_L g365 ( .A(n_366), .B(n_404), .C(n_419), .D(n_439), .E(n_449), .Y(n_365) );
NOR2xp33_ASAP7_75t_SL g366 ( .A(n_367), .B(n_384), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_373), .B1(n_376), .B2(n_378), .C(n_379), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI221xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_389), .B1(n_390), .B2(n_392), .C(n_393), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_389), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
OR2x2_ASAP7_75t_L g402 ( .A(n_397), .B(n_403), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B(n_411), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_425), .Y(n_419) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_436), .B2(n_438), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_435), .A2(n_450), .B(n_451), .C(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g453 ( .A(n_446), .Y(n_453) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx4_ASAP7_75t_L g771 ( .A(n_456), .Y(n_771) );
OAI22xp5_ASAP7_75t_SL g781 ( .A1(n_456), .A2(n_771), .B1(n_782), .B2(n_783), .Y(n_781) );
AND3x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_643), .C(n_739), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_585), .C(n_612), .Y(n_457) );
OAI211xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_495), .B(n_534), .C(n_558), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_477), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_460), .A2(n_536), .B(n_540), .C(n_546), .Y(n_535) );
OR2x2_ASAP7_75t_L g658 ( .A(n_460), .B(n_595), .Y(n_658) );
INVx2_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g625 ( .A(n_461), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_461), .B(n_596), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_461), .B(n_741), .Y(n_756) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_469), .Y(n_461) );
AND2x2_ASAP7_75t_L g542 ( .A(n_462), .B(n_478), .Y(n_542) );
INVx1_ASAP7_75t_L g562 ( .A(n_462), .Y(n_562) );
OR2x2_ASAP7_75t_L g577 ( .A(n_462), .B(n_486), .Y(n_577) );
INVx2_ASAP7_75t_L g583 ( .A(n_462), .Y(n_583) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_462), .Y(n_638) );
INVx1_ASAP7_75t_L g715 ( .A(n_462), .Y(n_715) );
NOR2x1_ASAP7_75t_SL g564 ( .A(n_469), .B(n_486), .Y(n_564) );
AND2x2_ASAP7_75t_L g594 ( .A(n_469), .B(n_583), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
OR2x2_ASAP7_75t_L g588 ( .A(n_477), .B(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_477), .B(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g716 ( .A(n_477), .Y(n_716) );
NAND2x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_486), .Y(n_477) );
OR2x2_ASAP7_75t_SL g576 ( .A(n_478), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g580 ( .A(n_478), .Y(n_580) );
INVx4_ASAP7_75t_L g596 ( .A(n_478), .Y(n_596) );
OR2x2_ASAP7_75t_L g611 ( .A(n_478), .B(n_544), .Y(n_611) );
AND2x2_ASAP7_75t_L g650 ( .A(n_478), .B(n_564), .Y(n_650) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_478), .Y(n_662) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
AND2x2_ASAP7_75t_L g543 ( .A(n_486), .B(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g595 ( .A(n_486), .B(n_596), .Y(n_595) );
BUFx2_ASAP7_75t_L g610 ( .A(n_486), .Y(n_610) );
AND2x2_ASAP7_75t_L g626 ( .A(n_486), .B(n_596), .Y(n_626) );
AND2x2_ASAP7_75t_L g639 ( .A(n_486), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g671 ( .A(n_486), .B(n_583), .Y(n_671) );
INVx2_ASAP7_75t_SL g741 ( .A(n_486), .Y(n_741) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_494), .Y(n_486) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NOR2xp67_ASAP7_75t_L g496 ( .A(n_497), .B(n_516), .Y(n_496) );
OAI211xp5_ASAP7_75t_L g612 ( .A1(n_497), .A2(n_613), .B(n_617), .C(n_633), .Y(n_612) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g708 ( .A(n_498), .B(n_547), .Y(n_708) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
INVx2_ASAP7_75t_L g557 ( .A(n_499), .Y(n_557) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_499), .B(n_548), .Y(n_568) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_499), .Y(n_572) );
AND2x2_ASAP7_75t_L g630 ( .A(n_499), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g704 ( .A(n_499), .Y(n_704) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_500), .Y(n_606) );
AND2x2_ASAP7_75t_L g649 ( .A(n_500), .B(n_508), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_506), .Y(n_501) );
INVx2_ASAP7_75t_L g539 ( .A(n_508), .Y(n_539) );
AND2x2_ASAP7_75t_L g599 ( .A(n_508), .B(n_548), .Y(n_599) );
INVx2_ASAP7_75t_L g631 ( .A(n_508), .Y(n_631) );
OR2x2_ASAP7_75t_L g654 ( .A(n_508), .B(n_519), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_516), .B(n_571), .Y(n_678) );
AND2x2_ASAP7_75t_L g712 ( .A(n_516), .B(n_648), .Y(n_712) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OAI31xp33_ASAP7_75t_SL g633 ( .A1(n_517), .A2(n_614), .A3(n_634), .B(n_641), .Y(n_633) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_518), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx3_ASAP7_75t_L g567 ( .A(n_519), .Y(n_567) );
AND2x2_ASAP7_75t_L g584 ( .A(n_519), .B(n_547), .Y(n_584) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
AND2x4_ASAP7_75t_L g574 ( .A(n_520), .B(n_521), .Y(n_574) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
NOR2x1p5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g719 ( .A(n_537), .Y(n_719) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_539), .B(n_548), .Y(n_601) );
AND2x2_ASAP7_75t_L g642 ( .A(n_539), .B(n_557), .Y(n_642) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
AND2x2_ASAP7_75t_L g622 ( .A(n_543), .B(n_580), .Y(n_622) );
AND2x2_ASAP7_75t_L g581 ( .A(n_544), .B(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_544), .Y(n_590) );
INVx2_ASAP7_75t_L g640 ( .A(n_544), .Y(n_640) );
AND2x2_ASAP7_75t_L g730 ( .A(n_544), .B(n_715), .Y(n_730) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g736 ( .A(n_546), .Y(n_736) );
NAND2x1p5_ASAP7_75t_L g546 ( .A(n_547), .B(n_556), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_547), .B(n_606), .Y(n_675) );
AND2x2_ASAP7_75t_L g723 ( .A(n_547), .B(n_649), .Y(n_723) );
INVx4_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g632 ( .A(n_548), .B(n_604), .Y(n_632) );
AND2x2_ASAP7_75t_L g641 ( .A(n_548), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g653 ( .A(n_548), .Y(n_653) );
BUFx2_ASAP7_75t_L g669 ( .A(n_548), .Y(n_669) );
AND2x4_ASAP7_75t_L g703 ( .A(n_548), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g748 ( .A(n_548), .B(n_649), .Y(n_748) );
OR2x6_ASAP7_75t_L g548 ( .A(n_549), .B(n_555), .Y(n_548) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AOI222xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_565), .B1(n_569), .B2(n_575), .C1(n_578), .C2(n_584), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_560), .A2(n_624), .B1(n_627), .B2(n_632), .Y(n_623) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
AND2x2_ASAP7_75t_L g607 ( .A(n_561), .B(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_SL g621 ( .A(n_561), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_561), .B(n_626), .Y(n_759) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g720 ( .A(n_562), .B(n_626), .Y(n_720) );
OR2x2_ASAP7_75t_L g697 ( .A(n_563), .B(n_579), .Y(n_697) );
OR2x2_ASAP7_75t_L g705 ( .A(n_563), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g689 ( .A(n_564), .B(n_582), .Y(n_689) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
OR2x2_ASAP7_75t_L g597 ( .A(n_567), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g747 ( .A(n_567), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g698 ( .A(n_568), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_568), .B(n_727), .Y(n_726) );
INVx2_ASAP7_75t_SL g733 ( .A(n_568), .Y(n_733) );
INVxp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx2_ASAP7_75t_L g718 ( .A(n_571), .Y(n_718) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g620 ( .A(n_572), .B(n_599), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_573), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g619 ( .A(n_573), .Y(n_619) );
NOR2x1_ASAP7_75t_L g628 ( .A(n_573), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g722 ( .A(n_573), .B(n_594), .Y(n_722) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g656 ( .A(n_574), .B(n_642), .Y(n_656) );
AND2x2_ASAP7_75t_L g699 ( .A(n_574), .B(n_631), .Y(n_699) );
AND2x4_ASAP7_75t_L g614 ( .A(n_575), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g755 ( .A(n_577), .B(n_611), .Y(n_755) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_579), .B(n_594), .Y(n_738) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_580), .B(n_594), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g721 ( .A1(n_580), .A2(n_621), .B(n_722), .C(n_723), .Y(n_721) );
AND2x2_ASAP7_75t_L g752 ( .A(n_580), .B(n_730), .Y(n_752) );
INVx1_ASAP7_75t_L g663 ( .A(n_581), .Y(n_663) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_584), .B(n_648), .Y(n_647) );
OAI21xp33_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_597), .B(n_600), .Y(n_585) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_591), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_588), .A2(n_741), .B1(n_742), .B2(n_744), .Y(n_740) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g616 ( .A(n_590), .Y(n_616) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp67_ASAP7_75t_L g637 ( .A(n_596), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g688 ( .A(n_596), .Y(n_688) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B(n_607), .Y(n_600) );
INVx1_ASAP7_75t_L g679 ( .A(n_601), .Y(n_679) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx2_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B(n_623), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
OR2x2_ASAP7_75t_L g664 ( .A(n_619), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g701 ( .A(n_619), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_619), .B(n_649), .Y(n_737) );
INVx1_ASAP7_75t_L g757 ( .A(n_620), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_622), .A2(n_725), .B1(n_728), .B2(n_731), .C(n_734), .Y(n_724) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI321xp33_ASAP7_75t_L g745 ( .A1(n_627), .A2(n_662), .A3(n_746), .B1(n_749), .B2(n_751), .C(n_753), .Y(n_745) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g686 ( .A(n_631), .Y(n_686) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g680 ( .A(n_636), .Y(n_680) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g706 ( .A(n_637), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_639), .A2(n_667), .B1(n_671), .B2(n_672), .C(n_677), .Y(n_666) );
INVxp67_ASAP7_75t_L g695 ( .A(n_640), .Y(n_695) );
INVx1_ASAP7_75t_L g665 ( .A(n_642), .Y(n_665) );
NOR2xp67_ASAP7_75t_L g643 ( .A(n_644), .B(n_690), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_666), .C(n_681), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_650), .B1(n_651), .B2(n_657), .C(n_659), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g764 ( .A(n_649), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_652), .B(n_655), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_653), .B(n_699), .Y(n_744) );
INVx2_ASAP7_75t_SL g676 ( .A(n_654), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_655), .A2(n_660), .B1(n_661), .B2(n_664), .Y(n_659) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_663), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_664), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g670 ( .A(n_665), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g709 ( .A1(n_667), .A2(n_710), .B1(n_712), .B2(n_713), .C1(n_717), .C2(n_720), .Y(n_709) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_668), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g743 ( .A(n_668), .B(n_722), .Y(n_743) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_676), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_676), .B(n_736), .Y(n_735) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B(n_680), .Y(n_677) );
NAND2xp33_ASAP7_75t_SL g681 ( .A(n_682), .B(n_687), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_687), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
NAND4xp25_ASAP7_75t_SL g690 ( .A(n_691), .B(n_709), .C(n_721), .D(n_724), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_696), .B(n_698), .C(n_700), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_697), .A2(n_701), .B1(n_705), .B2(n_707), .Y(n_700) );
INVx1_ASAP7_75t_L g727 ( .A(n_699), .Y(n_727) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_716), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_733), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B(n_738), .Y(n_734) );
NOR4xp25_ASAP7_75t_L g739 ( .A(n_740), .B(n_745), .C(n_758), .D(n_760), .Y(n_739) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx4_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx3_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
OAI22x1_ASAP7_75t_L g770 ( .A1(n_767), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
BUFx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
endmodule