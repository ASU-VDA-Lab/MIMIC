module fake_jpeg_25078_n_173 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_21),
.B1(n_19),
.B2(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_19),
.B1(n_27),
.B2(n_16),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_21),
.B1(n_19),
.B2(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_14),
.B1(n_28),
.B2(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_15),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_14),
.B(n_1),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_28),
.B(n_27),
.C(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_48),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_37),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_38),
.B1(n_44),
.B2(n_39),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_38),
.B1(n_45),
.B2(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_70),
.B1(n_79),
.B2(n_50),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_44),
.B(n_41),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_80),
.B(n_22),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_25),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_73),
.B(n_33),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_31),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_33),
.B(n_25),
.Y(n_86)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_50),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_36),
.B1(n_18),
.B2(n_16),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_13),
.B1(n_22),
.B2(n_24),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_91),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_92),
.B(n_63),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_23),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_96),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_23),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_69),
.B(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_20),
.B1(n_25),
.B2(n_33),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_23),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_54),
.C(n_23),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_70),
.C(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_79),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_116),
.B(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_106),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_66),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_63),
.C(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_83),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_63),
.B1(n_95),
.B2(n_87),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_81),
.B1(n_99),
.B2(n_98),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_107),
.B1(n_76),
.B2(n_54),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_96),
.B1(n_86),
.B2(n_72),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_108),
.B(n_113),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_103),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_135),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_100),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_133),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_120),
.C(n_126),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_17),
.C(n_20),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_140),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_141),
.B1(n_131),
.B2(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_128),
.B(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_148),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_0),
.B(n_1),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_33),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_153),
.C(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_138),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_138),
.B1(n_136),
.B2(n_2),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_155),
.A3(n_144),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_8),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_162),
.B(n_151),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_163),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_156),
.A2(n_145),
.B(n_3),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_161),
.A2(n_9),
.B(n_10),
.Y(n_167)
);

AOI21x1_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_2),
.B(n_3),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_5),
.C(n_8),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_9),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_160),
.B(n_5),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_167),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_170),
.B(n_10),
.C(n_33),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_10),
.B(n_25),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_31),
.B1(n_169),
.B2(n_49),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_31),
.Y(n_173)
);


endmodule