module fake_netlist_1_3453_n_32 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx3_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_1), .B(n_6), .Y(n_13) );
NAND2xp5_ASAP7_75t_SL g14 ( .A(n_1), .B(n_0), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_10), .B(n_6), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_3), .B(n_2), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_7), .B(n_8), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_12), .B(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_15), .B(n_2), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_12), .B1(n_15), .B2(n_16), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_15), .B(n_17), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_12), .Y(n_22) );
HB1xp67_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_23), .B(n_21), .Y(n_25) );
OAI222xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_14), .B1(n_16), .B2(n_13), .C1(n_15), .C2(n_17), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_13), .B1(n_4), .B2(n_5), .Y(n_27) );
NAND4xp75_ASAP7_75t_L g28 ( .A(n_26), .B(n_3), .C(n_4), .D(n_7), .Y(n_28) );
NAND2xp5_ASAP7_75t_SL g29 ( .A(n_27), .B(n_11), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
AOI21xp33_ASAP7_75t_SL g32 ( .A1(n_31), .A2(n_29), .B(n_9), .Y(n_32) );
endmodule