module fake_jpeg_4118_n_108 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_13),
.B1(n_15),
.B2(n_12),
.Y(n_35)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_R g44 ( 
.A(n_35),
.B(n_30),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_17),
.B1(n_20),
.B2(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_38),
.B1(n_21),
.B2(n_12),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_17),
.B1(n_20),
.B2(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_19),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_46),
.B(n_15),
.Y(n_57)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_51),
.B1(n_19),
.B2(n_12),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_52),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_29),
.B1(n_18),
.B2(n_13),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_34),
.B1(n_36),
.B2(n_33),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_55),
.B1(n_57),
.B2(n_61),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_32),
.C(n_42),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_22),
.C(n_16),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_33),
.B1(n_45),
.B2(n_51),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_23),
.A3(n_15),
.B1(n_13),
.B2(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_73),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_68),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_24),
.B(n_16),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_41),
.B1(n_24),
.B2(n_3),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_1),
.B(n_3),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_60),
.B1(n_62),
.B2(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_84),
.Y(n_85)
);

AOI322xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_62),
.A3(n_53),
.B1(n_61),
.B2(n_59),
.C1(n_63),
.C2(n_58),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_74),
.C(n_67),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_63),
.A3(n_58),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_1),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_4),
.B(n_7),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_69),
.C(n_6),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_56),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_77),
.C(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_82),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_74),
.B1(n_75),
.B2(n_8),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_81),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_78),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_94),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_78),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_91),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_76),
.C(n_83),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_97),
.B(n_98),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_83),
.B1(n_81),
.B2(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_7),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g102 ( 
.A(n_99),
.B(n_7),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_99),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_103),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_100),
.B(n_104),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_8),
.Y(n_108)
);


endmodule