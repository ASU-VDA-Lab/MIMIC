module fake_jpeg_25881_n_25 (n_3, n_2, n_1, n_0, n_4, n_5, n_25);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_25;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

INVx8_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_13),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_9),
.B(n_1),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_6),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_8),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_15)
);

AND2x6_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_3),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_18),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_17),
.B(n_9),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_8),
.C(n_14),
.Y(n_21)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_22),
.CI(n_10),
.CON(n_23),
.SN(n_23)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_11),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_23),
.A2(n_7),
.B(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);


endmodule