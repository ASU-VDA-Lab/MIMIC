module real_aes_15913_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_1634, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_1634;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1600;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_1612;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_602;
wire n_402;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1620;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1605;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_0), .A2(n_102), .B1(n_397), .B2(n_400), .Y(n_396) );
INVxp67_ASAP7_75t_SL g453 ( .A(n_0), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_1), .A2(n_75), .B1(n_619), .B2(n_628), .Y(n_627) );
INVxp33_ASAP7_75t_SL g675 ( .A(n_1), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_2), .Y(n_1013) );
INVx1_ASAP7_75t_L g1212 ( .A(n_3), .Y(n_1212) );
AOI221xp5_ASAP7_75t_L g1260 ( .A1(n_4), .A2(n_211), .B1(n_534), .B2(n_844), .C(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1288 ( .A(n_4), .Y(n_1288) );
INVx1_ASAP7_75t_L g347 ( .A(n_5), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g1160 ( .A(n_6), .Y(n_1160) );
INVx1_ASAP7_75t_L g781 ( .A(n_7), .Y(n_781) );
OAI221xp5_ASAP7_75t_SL g816 ( .A1(n_7), .A2(n_103), .B1(n_352), .B2(n_520), .C(n_724), .Y(n_816) );
INVx1_ASAP7_75t_L g1262 ( .A(n_8), .Y(n_1262) );
AOI221xp5_ASAP7_75t_L g1291 ( .A1(n_8), .A2(n_160), .B1(n_485), .B2(n_487), .C(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g862 ( .A(n_9), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_9), .A2(n_125), .B1(n_457), .B2(n_893), .Y(n_892) );
AOI21xp33_ASAP7_75t_L g1227 ( .A1(n_10), .A2(n_529), .B(n_625), .Y(n_1227) );
INVx1_ASAP7_75t_L g1248 ( .A(n_10), .Y(n_1248) );
AOI22xp5_ASAP7_75t_SL g1339 ( .A1(n_11), .A2(n_262), .B1(n_1322), .B2(n_1330), .Y(n_1339) );
OAI221xp5_ASAP7_75t_L g852 ( .A1(n_12), .A2(n_227), .B1(n_352), .B2(n_520), .C(n_823), .Y(n_852) );
OA222x2_ASAP7_75t_L g898 ( .A1(n_12), .A2(n_58), .B1(n_232), .B2(n_430), .C1(n_660), .C2(n_663), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g1535 ( .A1(n_13), .A2(n_155), .B1(n_389), .B2(n_548), .Y(n_1535) );
INVxp67_ASAP7_75t_SL g1568 ( .A(n_13), .Y(n_1568) );
INVx1_ASAP7_75t_L g517 ( .A(n_14), .Y(n_517) );
OAI221xp5_ASAP7_75t_SL g585 ( .A1(n_14), .A2(n_269), .B1(n_586), .B2(n_590), .C(n_594), .Y(n_585) );
INVx1_ASAP7_75t_L g298 ( .A(n_15), .Y(n_298) );
AND2x2_ASAP7_75t_L g327 ( .A(n_15), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g443 ( .A(n_15), .B(n_234), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_15), .B(n_308), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g1109 ( .A(n_16), .Y(n_1109) );
OAI22xp5_ASAP7_75t_L g1586 ( .A1(n_17), .A2(n_81), .B1(n_440), .B2(n_449), .Y(n_1586) );
OAI22xp33_ASAP7_75t_L g1619 ( .A1(n_17), .A2(n_47), .B1(n_397), .B2(n_400), .Y(n_1619) );
INVx1_ASAP7_75t_L g920 ( .A(n_18), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_18), .A2(n_258), .B1(n_349), .B2(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g1076 ( .A(n_19), .Y(n_1076) );
AOI22xp5_ASAP7_75t_L g1097 ( .A1(n_19), .A2(n_42), .B1(n_603), .B2(n_1050), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_20), .A2(n_130), .B1(n_366), .B2(n_373), .Y(n_960) );
INVxp67_ASAP7_75t_SL g995 ( .A(n_20), .Y(n_995) );
INVx2_ASAP7_75t_L g1317 ( .A(n_21), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_21), .B(n_1318), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_21), .B(n_120), .Y(n_1325) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_22), .A2(n_389), .B(n_391), .Y(n_388) );
INVx1_ASAP7_75t_L g476 ( .A(n_22), .Y(n_476) );
INVx1_ASAP7_75t_L g1011 ( .A(n_23), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_24), .A2(n_161), .B1(n_382), .B2(n_412), .Y(n_411) );
AOI32xp33_ASAP7_75t_L g455 ( .A1(n_24), .A2(n_456), .A3(n_459), .B1(n_464), .B2(n_1634), .Y(n_455) );
AOI22xp5_ASAP7_75t_SL g1353 ( .A1(n_25), .A2(n_145), .B1(n_1322), .B2(n_1330), .Y(n_1353) );
XNOR2x2_ASAP7_75t_L g1255 ( .A(n_26), .B(n_1256), .Y(n_1255) );
CKINVDCx5p33_ASAP7_75t_R g1116 ( .A(n_27), .Y(n_1116) );
AOI22xp5_ASAP7_75t_SL g1348 ( .A1(n_28), .A2(n_253), .B1(n_1319), .B2(n_1324), .Y(n_1348) );
INVx1_ASAP7_75t_L g969 ( .A(n_29), .Y(n_969) );
AND2x2_ASAP7_75t_L g394 ( .A(n_30), .B(n_395), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_30), .A2(n_161), .B1(n_489), .B2(n_490), .C(n_492), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g1137 ( .A1(n_31), .A2(n_263), .B1(n_300), .B2(n_1138), .Y(n_1137) );
OAI22xp33_ASAP7_75t_L g1169 ( .A1(n_31), .A2(n_263), .B1(n_1170), .B2(n_1173), .Y(n_1169) );
INVx1_ASAP7_75t_L g1220 ( .A(n_32), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_32), .A2(n_154), .B1(n_689), .B2(n_757), .Y(n_1243) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_33), .A2(n_87), .B1(n_631), .B2(n_632), .C(n_634), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_33), .A2(n_35), .B1(n_688), .B2(n_689), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_34), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_35), .A2(n_144), .B1(n_616), .B2(n_619), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g1120 ( .A(n_36), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_37), .A2(n_177), .B1(n_395), .B2(n_618), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_37), .A2(n_151), .B1(n_1044), .B2(n_1048), .Y(n_1047) );
AOI222xp33_ASAP7_75t_L g976 ( .A1(n_38), .A2(n_186), .B1(n_224), .B2(n_375), .C1(n_529), .C2(n_871), .Y(n_976) );
INVx1_ASAP7_75t_L g1001 ( .A(n_38), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_39), .B(n_385), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_39), .A2(n_275), .B1(n_485), .B2(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g908 ( .A(n_40), .Y(n_908) );
INVx1_ASAP7_75t_L g637 ( .A(n_41), .Y(n_637) );
OA222x2_ASAP7_75t_L g659 ( .A1(n_41), .A2(n_175), .B1(n_276), .B2(n_660), .C1(n_662), .C2(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g1085 ( .A(n_42), .Y(n_1085) );
AOI22xp5_ASAP7_75t_L g1313 ( .A1(n_43), .A2(n_183), .B1(n_1314), .B2(n_1319), .Y(n_1313) );
INVx1_ASAP7_75t_L g1082 ( .A(n_44), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_44), .A2(n_184), .B1(n_485), .B2(n_603), .Y(n_1099) );
INVx1_ASAP7_75t_L g1263 ( .A(n_45), .Y(n_1263) );
AOI221xp5_ASAP7_75t_L g1282 ( .A1(n_45), .A2(n_83), .B1(n_1283), .B2(n_1285), .C(n_1287), .Y(n_1282) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_46), .A2(n_210), .B1(n_621), .B2(n_622), .C(n_625), .Y(n_620) );
INVx1_ASAP7_75t_L g683 ( .A(n_46), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g1584 ( .A1(n_47), .A2(n_657), .B(n_1585), .C(n_1602), .Y(n_1584) );
INVx1_ASAP7_75t_L g1017 ( .A(n_48), .Y(n_1017) );
INVx1_ASAP7_75t_L g1102 ( .A(n_49), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_50), .A2(n_88), .B1(n_534), .B2(n_535), .Y(n_533) );
INVxp67_ASAP7_75t_SL g598 ( .A(n_50), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g1273 ( .A1(n_51), .A2(n_72), .B1(n_349), .B2(n_354), .C(n_360), .Y(n_1273) );
INVxp67_ASAP7_75t_SL g1278 ( .A(n_51), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g1367 ( .A1(n_52), .A2(n_112), .B1(n_1322), .B2(n_1368), .Y(n_1367) );
OAI21xp33_ASAP7_75t_L g910 ( .A1(n_53), .A2(n_660), .B(n_911), .Y(n_910) );
OAI221xp5_ASAP7_75t_L g944 ( .A1(n_53), .A2(n_61), .B1(n_733), .B2(n_945), .C(n_946), .Y(n_944) );
OAI211xp5_ASAP7_75t_SL g1208 ( .A1(n_54), .A2(n_948), .B(n_1209), .C(n_1213), .Y(n_1208) );
INVx1_ASAP7_75t_L g1233 ( .A(n_54), .Y(n_1233) );
AOI22xp5_ASAP7_75t_L g1321 ( .A1(n_55), .A2(n_187), .B1(n_1322), .B2(n_1324), .Y(n_1321) );
AOI22xp5_ASAP7_75t_L g1331 ( .A1(n_56), .A2(n_99), .B1(n_1314), .B2(n_1322), .Y(n_1331) );
INVx1_ASAP7_75t_L g341 ( .A(n_57), .Y(n_341) );
INVx1_ASAP7_75t_L g359 ( .A(n_57), .Y(n_359) );
INVx1_ASAP7_75t_L g850 ( .A(n_58), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_59), .A2(n_164), .B1(n_435), .B2(n_688), .Y(n_799) );
INVx1_ASAP7_75t_L g821 ( .A(n_59), .Y(n_821) );
INVx1_ASAP7_75t_L g921 ( .A(n_60), .Y(n_921) );
INVxp67_ASAP7_75t_SL g951 ( .A(n_61), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g1333 ( .A1(n_62), .A2(n_272), .B1(n_1314), .B2(n_1319), .Y(n_1333) );
OAI221xp5_ASAP7_75t_L g1065 ( .A1(n_63), .A2(n_123), .B1(n_366), .B2(n_373), .C(n_1066), .Y(n_1065) );
INVxp67_ASAP7_75t_SL g1092 ( .A(n_63), .Y(n_1092) );
AOI221xp5_ASAP7_75t_L g962 ( .A1(n_64), .A2(n_168), .B1(n_963), .B2(n_965), .C(n_967), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_64), .A2(n_229), .B1(n_486), .B2(n_997), .C(n_999), .Y(n_996) );
OAI221xp5_ASAP7_75t_L g959 ( .A1(n_65), .A2(n_250), .B1(n_349), .B2(n_354), .C(n_360), .Y(n_959) );
OAI21xp33_ASAP7_75t_SL g987 ( .A1(n_65), .A2(n_505), .B(n_663), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g1609 ( .A1(n_66), .A2(n_245), .B1(n_366), .B2(n_373), .Y(n_1609) );
INVxp67_ASAP7_75t_SL g1621 ( .A(n_66), .Y(n_1621) );
INVx1_ASAP7_75t_L g291 ( .A(n_67), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g1272 ( .A1(n_68), .A2(n_220), .B1(n_366), .B2(n_373), .Y(n_1272) );
INVx1_ASAP7_75t_L g1281 ( .A(n_68), .Y(n_1281) );
INVx2_ASAP7_75t_L g344 ( .A(n_69), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g1117 ( .A(n_70), .Y(n_1117) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_71), .A2(n_198), .B1(n_397), .B2(n_400), .Y(n_1259) );
INVx1_ASAP7_75t_L g1279 ( .A(n_71), .Y(n_1279) );
INVx1_ASAP7_75t_L g1301 ( .A(n_72), .Y(n_1301) );
AOI22xp5_ASAP7_75t_L g1349 ( .A1(n_73), .A2(n_76), .B1(n_1314), .B2(n_1322), .Y(n_1349) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_74), .A2(n_79), .B1(n_397), .B2(n_400), .Y(n_970) );
INVxp67_ASAP7_75t_SL g982 ( .A(n_74), .Y(n_982) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_75), .Y(n_686) );
AOI22xp33_ASAP7_75t_SL g1542 ( .A1(n_77), .A2(n_80), .B1(n_389), .B2(n_1543), .Y(n_1542) );
AOI221xp5_ASAP7_75t_L g1556 ( .A1(n_77), .A2(n_155), .B1(n_486), .B2(n_1557), .C(n_1559), .Y(n_1556) );
INVx1_ASAP7_75t_L g1201 ( .A(n_78), .Y(n_1201) );
INVx1_ASAP7_75t_L g986 ( .A(n_79), .Y(n_986) );
INVxp67_ASAP7_75t_SL g1570 ( .A(n_80), .Y(n_1570) );
OAI221xp5_ASAP7_75t_L g1608 ( .A1(n_81), .A2(n_132), .B1(n_349), .B2(n_354), .C(n_360), .Y(n_1608) );
AOI22xp33_ASAP7_75t_SL g1536 ( .A1(n_82), .A2(n_196), .B1(n_1031), .B2(n_1537), .Y(n_1536) );
AOI22xp33_ASAP7_75t_L g1560 ( .A1(n_82), .A2(n_142), .B1(n_1043), .B2(n_1044), .Y(n_1560) );
AOI221xp5_ASAP7_75t_L g1264 ( .A1(n_83), .A2(n_212), .B1(n_844), .B2(n_1265), .C(n_1267), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_84), .A2(n_248), .B1(n_529), .B2(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_84), .A2(n_222), .B1(n_489), .B2(n_490), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_85), .A2(n_189), .B1(n_671), .B2(n_795), .C(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g822 ( .A(n_85), .Y(n_822) );
INVx1_ASAP7_75t_L g958 ( .A(n_86), .Y(n_958) );
OAI21xp33_ASAP7_75t_L g983 ( .A1(n_86), .A2(n_430), .B(n_984), .Y(n_983) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_87), .A2(n_210), .B1(n_669), .B2(n_671), .C(n_672), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_88), .A2(n_109), .B1(n_569), .B2(n_574), .C(n_576), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g856 ( .A(n_89), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_90), .A2(n_255), .B1(n_1142), .B2(n_1145), .Y(n_1141) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_90), .A2(n_255), .B1(n_1191), .B2(n_1193), .Y(n_1190) );
INVx1_ASAP7_75t_L g866 ( .A(n_91), .Y(n_866) );
AOI221x1_ASAP7_75t_SL g883 ( .A1(n_91), .A2(n_110), .B1(n_435), .B2(n_795), .C(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g650 ( .A(n_92), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_92), .B(n_657), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g1544 ( .A1(n_93), .A2(n_268), .B1(n_1545), .B2(n_1548), .Y(n_1544) );
INVx1_ASAP7_75t_L g1563 ( .A(n_93), .Y(n_1563) );
INVx1_ASAP7_75t_L g1083 ( .A(n_94), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_94), .A2(n_236), .B1(n_435), .B2(n_688), .Y(n_1098) );
AOI22xp5_ASAP7_75t_L g1329 ( .A1(n_95), .A2(n_195), .B1(n_1319), .B2(n_1330), .Y(n_1329) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_96), .A2(n_106), .B1(n_1021), .B2(n_1023), .Y(n_1020) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_96), .A2(n_136), .B1(n_456), .B2(n_486), .C(n_576), .Y(n_1041) );
INVx1_ASAP7_75t_L g1230 ( .A(n_97), .Y(n_1230) );
XOR2x1_ASAP7_75t_L g318 ( .A(n_98), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g1598 ( .A(n_100), .Y(n_1598) );
AOI221xp5_ASAP7_75t_L g1221 ( .A1(n_101), .A2(n_149), .B1(n_634), .B2(n_1222), .C(n_1223), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_101), .A2(n_201), .B1(n_566), .B2(n_757), .Y(n_1249) );
INVx1_ASAP7_75t_L g320 ( .A(n_102), .Y(n_320) );
INVx1_ASAP7_75t_L g790 ( .A(n_103), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_104), .Y(n_1072) );
INVx1_ASAP7_75t_L g847 ( .A(n_105), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_105), .A2(n_227), .B1(n_895), .B2(n_897), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g1049 ( .A1(n_106), .A2(n_213), .B1(n_574), .B2(n_1050), .C(n_1051), .Y(n_1049) );
INVx1_ASAP7_75t_L g651 ( .A(n_107), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_107), .A2(n_192), .B1(n_440), .B2(n_449), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g777 ( .A1(n_108), .A2(n_279), .B1(n_674), .B2(n_778), .C(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g806 ( .A(n_108), .Y(n_806) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_109), .A2(n_171), .B1(n_524), .B2(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g878 ( .A(n_110), .Y(n_878) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_111), .Y(n_293) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_111), .B(n_291), .Y(n_1315) );
CKINVDCx5p33_ASAP7_75t_R g732 ( .A(n_113), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_114), .A2(n_169), .B1(n_538), .B2(n_632), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_114), .A2(n_115), .B1(n_689), .B2(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g735 ( .A(n_115), .Y(n_735) );
OAI21xp5_ASAP7_75t_SL g1055 ( .A1(n_116), .A2(n_557), .B(n_1056), .Y(n_1055) );
AOI22xp5_ASAP7_75t_L g1370 ( .A1(n_117), .A2(n_170), .B1(n_1314), .B2(n_1319), .Y(n_1370) );
AOI22xp33_ASAP7_75t_SL g917 ( .A1(n_118), .A2(n_191), .B1(n_485), .B2(n_797), .Y(n_917) );
AOI221xp5_ASAP7_75t_L g937 ( .A1(n_118), .A2(n_179), .B1(n_625), .B2(n_631), .C(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g527 ( .A(n_119), .Y(n_527) );
INVx1_ASAP7_75t_L g1318 ( .A(n_120), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_120), .B(n_1317), .Y(n_1323) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_121), .A2(n_275), .B1(n_404), .B2(n_409), .C(n_410), .Y(n_403) );
INVx1_ASAP7_75t_L g478 ( .A(n_121), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_122), .A2(n_696), .B1(n_697), .B2(n_765), .Y(n_695) );
INVx1_ASAP7_75t_L g765 ( .A(n_122), .Y(n_765) );
INVx1_ASAP7_75t_L g1101 ( .A(n_123), .Y(n_1101) );
AOI22xp5_ASAP7_75t_L g1340 ( .A1(n_124), .A2(n_193), .B1(n_1314), .B2(n_1319), .Y(n_1340) );
INVx1_ASAP7_75t_L g872 ( .A(n_125), .Y(n_872) );
XNOR2xp5_ASAP7_75t_L g1007 ( .A(n_126), .B(n_1008), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_127), .A2(n_265), .B1(n_366), .B2(n_373), .Y(n_365) );
INVxp33_ASAP7_75t_L g503 ( .A(n_127), .Y(n_503) );
INVx1_ASAP7_75t_L g785 ( .A(n_128), .Y(n_785) );
OAI21xp33_ASAP7_75t_L g814 ( .A1(n_128), .A2(n_552), .B(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g346 ( .A(n_129), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_129), .B(n_344), .Y(n_369) );
INVx1_ASAP7_75t_L g415 ( .A(n_129), .Y(n_415) );
INVxp67_ASAP7_75t_SL g979 ( .A(n_130), .Y(n_979) );
INVxp67_ASAP7_75t_SL g1226 ( .A(n_131), .Y(n_1226) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_131), .A2(n_149), .B1(n_1239), .B2(n_1241), .Y(n_1238) );
INVxp67_ASAP7_75t_SL g1604 ( .A(n_132), .Y(n_1604) );
OAI221xp5_ASAP7_75t_L g348 ( .A1(n_133), .A2(n_166), .B1(n_349), .B2(n_354), .C(n_360), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_133), .B(n_461), .Y(n_460) );
XOR2xp5_ASAP7_75t_L g837 ( .A(n_134), .B(n_838), .Y(n_837) );
AOI221xp5_ASAP7_75t_L g1599 ( .A1(n_135), .A2(n_156), .B1(n_466), .B2(n_1594), .C(n_1600), .Y(n_1599) );
AOI221xp5_ASAP7_75t_L g1616 ( .A1(n_135), .A2(n_167), .B1(n_389), .B2(n_619), .C(n_1617), .Y(n_1616) );
AOI221xp5_ASAP7_75t_L g1028 ( .A1(n_136), .A2(n_151), .B1(n_534), .B2(n_1023), .C(n_1029), .Y(n_1028) );
OA22x2_ASAP7_75t_L g1580 ( .A1(n_137), .A2(n_1581), .B1(n_1622), .B2(n_1623), .Y(n_1580) );
CKINVDCx5p33_ASAP7_75t_R g1622 ( .A(n_137), .Y(n_1622) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_138), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_138), .Y(n_772) );
AOI22xp33_ASAP7_75t_SL g918 ( .A1(n_139), .A2(n_259), .B1(n_689), .B2(n_803), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_139), .A2(n_219), .B1(n_389), .B2(n_631), .C(n_634), .Y(n_939) );
CKINVDCx5p33_ASAP7_75t_R g868 ( .A(n_140), .Y(n_868) );
INVx1_ASAP7_75t_L g1086 ( .A(n_141), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_141), .A2(n_197), .B1(n_489), .B2(n_490), .Y(n_1100) );
AOI22xp33_ASAP7_75t_SL g1539 ( .A1(n_142), .A2(n_243), .B1(n_1031), .B2(n_1537), .Y(n_1539) );
INVx1_ASAP7_75t_L g1597 ( .A(n_143), .Y(n_1597) );
AOI221xp5_ASAP7_75t_L g1611 ( .A1(n_143), .A2(n_281), .B1(n_381), .B2(n_619), .C(n_1612), .Y(n_1611) );
INVxp67_ASAP7_75t_SL g673 ( .A(n_144), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g848 ( .A1(n_146), .A2(n_152), .B1(n_407), .B2(n_623), .Y(n_848) );
INVx1_ASAP7_75t_L g901 ( .A(n_146), .Y(n_901) );
INVx1_ASAP7_75t_L g1271 ( .A(n_147), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_148), .A2(n_199), .B1(n_749), .B2(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g832 ( .A(n_148), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_150), .A2(n_1206), .B1(n_1253), .B2(n_1254), .Y(n_1205) );
INVx1_ASAP7_75t_L g1254 ( .A(n_150), .Y(n_1254) );
INVx1_ASAP7_75t_L g900 ( .A(n_152), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g1552 ( .A1(n_153), .A2(n_178), .B1(n_557), .B2(n_701), .Y(n_1552) );
OAI211xp5_ASAP7_75t_SL g1554 ( .A1(n_153), .A2(n_564), .B(n_1555), .C(n_1561), .Y(n_1554) );
AOI22xp33_ASAP7_75t_SL g1228 ( .A1(n_154), .A2(n_201), .B1(n_412), .B2(n_632), .Y(n_1228) );
INVx1_ASAP7_75t_L g1615 ( .A(n_156), .Y(n_1615) );
INVx1_ASAP7_75t_L g1214 ( .A(n_157), .Y(n_1214) );
OAI221xp5_ASAP7_75t_L g1235 ( .A1(n_157), .A2(n_200), .B1(n_897), .B2(n_1236), .C(n_1237), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_158), .A2(n_218), .B1(n_803), .B2(n_924), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_158), .A2(n_259), .B1(n_389), .B2(n_412), .Y(n_936) );
AOI221xp5_ASAP7_75t_SL g794 ( .A1(n_159), .A2(n_180), .B1(n_671), .B2(n_795), .C(n_798), .Y(n_794) );
INVx1_ASAP7_75t_L g825 ( .A(n_159), .Y(n_825) );
INVx1_ASAP7_75t_L g1268 ( .A(n_160), .Y(n_1268) );
AOI22xp5_ASAP7_75t_L g1371 ( .A1(n_162), .A2(n_190), .B1(n_1322), .B2(n_1368), .Y(n_1371) );
BUFx3_ASAP7_75t_L g338 ( .A(n_163), .Y(n_338) );
INVx1_ASAP7_75t_L g834 ( .A(n_164), .Y(n_834) );
INVx1_ASAP7_75t_L g1215 ( .A(n_165), .Y(n_1215) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_166), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g1592 ( .A1(n_167), .A2(n_215), .B1(n_492), .B2(n_1593), .C(n_1594), .Y(n_1592) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_168), .B(n_602), .Y(n_989) );
AOI22xp33_ASAP7_75t_SL g747 ( .A1(n_169), .A2(n_240), .B1(n_748), .B2(n_749), .Y(n_747) );
INVxp67_ASAP7_75t_SL g600 ( .A(n_171), .Y(n_600) );
INVx1_ASAP7_75t_L g968 ( .A(n_172), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g1334 ( .A1(n_173), .A2(n_223), .B1(n_1322), .B2(n_1330), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_174), .Y(n_305) );
INVx1_ASAP7_75t_L g653 ( .A(n_175), .Y(n_653) );
INVx1_ASAP7_75t_L g912 ( .A(n_176), .Y(n_912) );
AOI22xp33_ASAP7_75t_SL g1042 ( .A1(n_177), .A2(n_267), .B1(n_1043), .B2(n_1044), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_179), .A2(n_219), .B1(n_927), .B2(n_928), .Y(n_926) );
INVx1_ASAP7_75t_L g831 ( .A(n_180), .Y(n_831) );
OAI222xp33_ASAP7_75t_L g550 ( .A1(n_181), .A2(n_221), .B1(n_241), .B2(n_551), .C1(n_557), .C2(n_559), .Y(n_550) );
OAI211xp5_ASAP7_75t_L g563 ( .A1(n_181), .A2(n_564), .B(n_567), .C(n_579), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_182), .Y(n_792) );
INVx1_ASAP7_75t_L g1075 ( .A(n_184), .Y(n_1075) );
INVx1_ASAP7_75t_L g1164 ( .A(n_185), .Y(n_1164) );
OAI211xp5_ASAP7_75t_L g1176 ( .A1(n_185), .A2(n_1177), .B(n_1179), .C(n_1181), .Y(n_1176) );
INVx1_ASAP7_75t_L g992 ( .A(n_186), .Y(n_992) );
INVx1_ASAP7_75t_L g712 ( .A(n_188), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g750 ( .A1(n_188), .A2(n_663), .B1(n_751), .B2(n_759), .C(n_760), .Y(n_750) );
INVx1_ASAP7_75t_L g835 ( .A(n_189), .Y(n_835) );
XOR2xp5_ASAP7_75t_L g1527 ( .A(n_190), .B(n_1528), .Y(n_1527) );
AOI22xp5_ASAP7_75t_L g1578 ( .A1(n_190), .A2(n_1579), .B1(n_1625), .B2(n_1628), .Y(n_1578) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_191), .A2(n_218), .B1(n_412), .B2(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g636 ( .A(n_192), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g1110 ( .A(n_194), .Y(n_1110) );
AOI221xp5_ASAP7_75t_L g1571 ( .A1(n_196), .A2(n_243), .B1(n_602), .B2(n_604), .C(n_928), .Y(n_1571) );
INVx1_ASAP7_75t_L g1079 ( .A(n_197), .Y(n_1079) );
INVxp67_ASAP7_75t_SL g1299 ( .A(n_198), .Y(n_1299) );
INVx1_ASAP7_75t_L g828 ( .A(n_199), .Y(n_828) );
INVx1_ASAP7_75t_L g1231 ( .A(n_200), .Y(n_1231) );
CKINVDCx5p33_ASAP7_75t_R g703 ( .A(n_202), .Y(n_703) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_203), .Y(n_304) );
INVx1_ASAP7_75t_L g1068 ( .A(n_204), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_204), .A2(n_206), .B1(n_440), .B2(n_449), .Y(n_1095) );
OAI211xp5_ASAP7_75t_L g1151 ( .A1(n_205), .A2(n_1152), .B(n_1155), .C(n_1158), .Y(n_1151) );
INVx1_ASAP7_75t_L g1189 ( .A(n_205), .Y(n_1189) );
INVx1_ASAP7_75t_L g1071 ( .A(n_206), .Y(n_1071) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_207), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g1121 ( .A(n_208), .Y(n_1121) );
CKINVDCx5p33_ASAP7_75t_R g1551 ( .A(n_209), .Y(n_1551) );
INVx1_ASAP7_75t_L g1293 ( .A(n_211), .Y(n_1293) );
INVx1_ASAP7_75t_L g1296 ( .A(n_212), .Y(n_1296) );
AOI22xp33_ASAP7_75t_SL g1030 ( .A1(n_213), .A2(n_267), .B1(n_1021), .B2(n_1031), .Y(n_1030) );
CKINVDCx5p33_ASAP7_75t_R g1114 ( .A(n_214), .Y(n_1114) );
INVx1_ASAP7_75t_L g1613 ( .A(n_215), .Y(n_1613) );
INVx1_ASAP7_75t_L g379 ( .A(n_216), .Y(n_379) );
INVx1_ASAP7_75t_L g1603 ( .A(n_217), .Y(n_1603) );
INVxp67_ASAP7_75t_SL g1275 ( .A(n_220), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_222), .A2(n_246), .B1(n_541), .B2(n_543), .Y(n_540) );
AOI21xp33_ASAP7_75t_L g993 ( .A1(n_224), .A2(n_456), .B(n_994), .Y(n_993) );
OAI211xp5_ASAP7_75t_L g1069 ( .A1(n_225), .A2(n_335), .B(n_360), .C(n_1070), .Y(n_1069) );
INVxp33_ASAP7_75t_SL g1094 ( .A(n_225), .Y(n_1094) );
INVx1_ASAP7_75t_L g1532 ( .A(n_226), .Y(n_1532) );
OAI221xp5_ASAP7_75t_SL g1564 ( .A1(n_226), .A2(n_278), .B1(n_1565), .B2(n_1566), .C(n_1567), .Y(n_1564) );
INVx1_ASAP7_75t_L g1035 ( .A(n_228), .Y(n_1035) );
AOI21xp33_ASAP7_75t_L g971 ( .A1(n_229), .A2(n_972), .B(n_975), .Y(n_971) );
INVx1_ASAP7_75t_L g699 ( .A(n_230), .Y(n_699) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_231), .Y(n_704) );
OAI221xp5_ASAP7_75t_L g720 ( .A1(n_231), .A2(n_360), .B1(n_366), .B2(n_721), .C(n_730), .Y(n_720) );
INVx1_ASAP7_75t_L g845 ( .A(n_232), .Y(n_845) );
INVx1_ASAP7_75t_L g1016 ( .A(n_233), .Y(n_1016) );
BUFx3_ASAP7_75t_L g308 ( .A(n_234), .Y(n_308) );
INVx1_ASAP7_75t_L g328 ( .A(n_234), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g1112 ( .A(n_235), .Y(n_1112) );
INVx1_ASAP7_75t_L g1078 ( .A(n_236), .Y(n_1078) );
INVx1_ASAP7_75t_L g693 ( .A(n_237), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_238), .A2(n_541), .B(n_625), .Y(n_718) );
INVx1_ASAP7_75t_L g745 ( .A(n_238), .Y(n_745) );
INVx1_ASAP7_75t_L g1210 ( .A(n_239), .Y(n_1210) );
INVx1_ASAP7_75t_L g729 ( .A(n_240), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g709 ( .A(n_242), .Y(n_709) );
INVx1_ASAP7_75t_L g325 ( .A(n_244), .Y(n_325) );
INVx2_ASAP7_75t_L g419 ( .A(n_244), .Y(n_419) );
INVx1_ASAP7_75t_L g434 ( .A(n_244), .Y(n_434) );
INVxp67_ASAP7_75t_SL g1605 ( .A(n_245), .Y(n_1605) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_246), .A2(n_248), .B1(n_456), .B2(n_602), .C(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g1269 ( .A(n_247), .Y(n_1269) );
INVx1_ASAP7_75t_L g1038 ( .A(n_249), .Y(n_1038) );
INVx1_ASAP7_75t_L g985 ( .A(n_250), .Y(n_985) );
INVx1_ASAP7_75t_L g522 ( .A(n_251), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g1352 ( .A1(n_252), .A2(n_271), .B1(n_1314), .B2(n_1319), .Y(n_1352) );
XOR2x2_ASAP7_75t_L g954 ( .A(n_254), .B(n_955), .Y(n_954) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_256), .Y(n_714) );
INVx1_ASAP7_75t_L g1365 ( .A(n_257), .Y(n_1365) );
INVx1_ASAP7_75t_L g913 ( .A(n_258), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_260), .B(n_762), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_261), .Y(n_874) );
OAI21xp33_ASAP7_75t_SL g1063 ( .A1(n_264), .A2(n_657), .B(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1067 ( .A(n_264), .Y(n_1067) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_265), .Y(n_421) );
INVx1_ASAP7_75t_L g1218 ( .A(n_266), .Y(n_1218) );
INVx1_ASAP7_75t_L g1562 ( .A(n_268), .Y(n_1562) );
INVx1_ASAP7_75t_L g514 ( .A(n_269), .Y(n_514) );
XNOR2xp5_ASAP7_75t_L g509 ( .A(n_270), .B(n_510), .Y(n_509) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_272), .Y(n_904) );
NAND2xp33_ASAP7_75t_SL g1591 ( .A(n_273), .B(n_680), .Y(n_1591) );
INVx1_ASAP7_75t_L g1618 ( .A(n_273), .Y(n_1618) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_274), .Y(n_780) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_276), .A2(n_280), .B1(n_644), .B2(n_645), .C(n_649), .Y(n_643) );
INVx1_ASAP7_75t_L g711 ( .A(n_277), .Y(n_711) );
INVx1_ASAP7_75t_L g1533 ( .A(n_278), .Y(n_1533) );
INVx1_ASAP7_75t_L g808 ( .A(n_279), .Y(n_808) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_280), .Y(n_665) );
INVx1_ASAP7_75t_L g1589 ( .A(n_281), .Y(n_1589) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_309), .B(n_1304), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx4f_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_294), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g1577 ( .A(n_288), .B(n_297), .Y(n_1577) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g1627 ( .A(n_290), .B(n_293), .Y(n_1627) );
INVx1_ASAP7_75t_L g1630 ( .A(n_290), .Y(n_1630) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g1632 ( .A(n_293), .B(n_1630), .Y(n_1632) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g1166 ( .A(n_297), .B(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x4_ASAP7_75t_L g496 ( .A(n_298), .B(n_308), .Y(n_496) );
AND2x4_ASAP7_75t_L g605 ( .A(n_298), .B(n_307), .Y(n_605) );
AND2x4_ASAP7_75t_SL g1576 ( .A(n_299), .B(n_1577), .Y(n_1576) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x6_ASAP7_75t_L g300 ( .A(n_301), .B(n_306), .Y(n_300) );
BUFx4f_ASAP7_75t_L g477 ( .A(n_301), .Y(n_477) );
OR2x6_ASAP7_75t_L g1144 ( .A(n_301), .B(n_1140), .Y(n_1144) );
INVx1_ASAP7_75t_L g1295 ( .A(n_301), .Y(n_1295) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx4f_ASAP7_75t_L g597 ( .A(n_302), .Y(n_597) );
INVx3_ASAP7_75t_L g886 ( .A(n_302), .Y(n_886) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx2_ASAP7_75t_L g330 ( .A(n_304), .Y(n_330) );
AND2x2_ASAP7_75t_L g425 ( .A(n_304), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g438 ( .A(n_304), .Y(n_438) );
INVx1_ASAP7_75t_L g452 ( .A(n_304), .Y(n_452) );
AND2x2_ASAP7_75t_L g458 ( .A(n_304), .B(n_305), .Y(n_458) );
NAND2x1_ASAP7_75t_L g463 ( .A(n_304), .B(n_305), .Y(n_463) );
INVx1_ASAP7_75t_L g331 ( .A(n_305), .Y(n_331) );
INVx2_ASAP7_75t_L g426 ( .A(n_305), .Y(n_426) );
AND2x2_ASAP7_75t_L g437 ( .A(n_305), .B(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g446 ( .A(n_305), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_305), .B(n_438), .Y(n_483) );
OR2x2_ASAP7_75t_L g682 ( .A(n_305), .B(n_330), .Y(n_682) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g1157 ( .A(n_307), .Y(n_1157) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx2_ASAP7_75t_L g1150 ( .A(n_308), .Y(n_1150) );
AND2x4_ASAP7_75t_L g1163 ( .A(n_308), .B(n_451), .Y(n_1163) );
OAI22xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_1057), .B2(n_1058), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B1(n_1004), .B2(n_1005), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
XNOR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_767), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_609), .B2(n_766), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OA22x2_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_508), .B2(n_509), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AO211x2_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_321), .B(n_332), .C(n_427), .Y(n_319) );
INVx3_ASAP7_75t_L g657 ( .A(n_321), .Y(n_657) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_321), .A2(n_422), .B1(n_699), .B2(n_700), .C1(n_703), .C2(n_704), .Y(n_698) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_321), .A2(n_422), .B1(n_900), .B2(n_901), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_321), .B(n_908), .Y(n_907) );
AOI211xp5_ASAP7_75t_L g981 ( .A1(n_321), .A2(n_982), .B(n_983), .C(n_987), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g1250 ( .A1(n_321), .A2(n_1210), .B1(n_1230), .B2(n_1251), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_321), .B(n_1299), .Y(n_1298) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
AND2x4_ASAP7_75t_L g422 ( .A(n_322), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g449 ( .A(n_323), .B(n_450), .Y(n_449) );
INVxp67_ASAP7_75t_L g560 ( .A(n_323), .Y(n_560) );
OR2x2_ASAP7_75t_L g897 ( .A(n_323), .B(n_450), .Y(n_897) );
INVx1_ASAP7_75t_L g1167 ( .A(n_323), .Y(n_1167) );
BUFx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g495 ( .A(n_324), .Y(n_495) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g581 ( .A(n_326), .Y(n_581) );
BUFx6f_ASAP7_75t_L g1037 ( .A(n_326), .Y(n_1037) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_L g423 ( .A(n_327), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_327), .B(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g565 ( .A(n_327), .B(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g584 ( .A(n_327), .B(n_424), .Y(n_584) );
AND2x4_ASAP7_75t_SL g589 ( .A(n_327), .B(n_457), .Y(n_589) );
BUFx2_ASAP7_75t_L g782 ( .A(n_327), .Y(n_782) );
HB1xp67_ASAP7_75t_L g1140 ( .A(n_328), .Y(n_1140) );
INVx3_ASAP7_75t_L g491 ( .A(n_329), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_329), .B(n_443), .Y(n_502) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_329), .Y(n_688) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_376), .B(n_416), .C(n_420), .Y(n_332) );
AOI211xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_347), .B(n_348), .C(n_365), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_334), .A2(n_640), .B1(n_643), .B2(n_653), .Y(n_639) );
INVx2_ASAP7_75t_L g948 ( .A(n_334), .Y(n_948) );
AOI211xp5_ASAP7_75t_SL g957 ( .A1(n_334), .A2(n_958), .B(n_959), .C(n_960), .Y(n_957) );
AOI211xp5_ASAP7_75t_SL g1270 ( .A1(n_334), .A2(n_1271), .B(n_1272), .C(n_1273), .Y(n_1270) );
AOI211xp5_ASAP7_75t_SL g1607 ( .A1(n_334), .A2(n_1603), .B(n_1608), .C(n_1609), .Y(n_1607) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x6_ASAP7_75t_L g559 ( .A(n_335), .B(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g701 ( .A(n_335), .B(n_560), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_336), .B(n_342), .Y(n_335) );
INVx8_ASAP7_75t_L g390 ( .A(n_336), .Y(n_390) );
AND2x2_ASAP7_75t_L g398 ( .A(n_336), .B(n_399), .Y(n_398) );
BUFx3_ASAP7_75t_L g618 ( .A(n_336), .Y(n_618) );
BUFx3_ASAP7_75t_L g633 ( .A(n_336), .Y(n_633) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
AND2x4_ASAP7_75t_L g371 ( .A(n_337), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_338), .Y(n_353) );
AND2x4_ASAP7_75t_L g402 ( .A(n_338), .B(n_358), .Y(n_402) );
OR2x2_ASAP7_75t_L g408 ( .A(n_338), .B(n_340), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_338), .B(n_359), .Y(n_555) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g372 ( .A(n_341), .Y(n_372) );
AND2x6_ASAP7_75t_L g350 ( .A(n_342), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g355 ( .A(n_342), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
AND2x4_ASAP7_75t_L g516 ( .A(n_342), .B(n_500), .Y(n_516) );
AND2x4_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_343), .B(n_415), .Y(n_414) );
NAND3x1_ASAP7_75t_L g545 ( .A(n_343), .B(n_415), .C(n_546), .Y(n_545) );
OR2x4_ASAP7_75t_L g1172 ( .A(n_343), .B(n_408), .Y(n_1172) );
INVx1_ASAP7_75t_L g1175 ( .A(n_343), .Y(n_1175) );
AND2x4_ASAP7_75t_L g1180 ( .A(n_343), .B(n_402), .Y(n_1180) );
OR2x6_ASAP7_75t_L g1195 ( .A(n_343), .B(n_648), .Y(n_1195) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g393 ( .A(n_344), .Y(n_393) );
NAND2xp33_ASAP7_75t_SL g626 ( .A(n_344), .B(n_346), .Y(n_626) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g392 ( .A(n_346), .B(n_393), .Y(n_392) );
AND3x4_ASAP7_75t_L g532 ( .A(n_346), .B(n_393), .C(n_418), .Y(n_532) );
HB1xp67_ASAP7_75t_L g1198 ( .A(n_346), .Y(n_1198) );
AOI222xp33_ASAP7_75t_L g428 ( .A1(n_347), .A2(n_429), .B1(n_439), .B2(n_447), .C1(n_448), .C2(n_453), .Y(n_428) );
INVx4_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_350), .A2(n_355), .B1(n_636), .B2(n_637), .C(n_638), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_350), .A2(n_355), .B1(n_711), .B2(n_712), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_350), .A2(n_355), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
AOI221xp5_ASAP7_75t_L g1213 ( .A1(n_350), .A2(n_355), .B1(n_638), .B2(n_1214), .C(n_1215), .Y(n_1213) );
AND2x2_ASAP7_75t_L g515 ( .A(n_351), .B(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_353), .B(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g375 ( .A(n_353), .B(n_357), .Y(n_375) );
BUFx2_ASAP7_75t_L g1185 ( .A(n_353), .Y(n_1185) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g934 ( .A(n_355), .Y(n_934) );
INVx1_ASAP7_75t_L g520 ( .A(n_356), .Y(n_520) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g363 ( .A(n_359), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_360), .Y(n_638) );
OR2x6_ASAP7_75t_L g360 ( .A(n_361), .B(n_364), .Y(n_360) );
INVx1_ASAP7_75t_L g409 ( .A(n_361), .Y(n_409) );
INVx1_ASAP7_75t_L g974 ( .A(n_361), .Y(n_974) );
INVx1_ASAP7_75t_L g1178 ( .A(n_361), .Y(n_1178) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_362), .Y(n_387) );
BUFx3_ASAP7_75t_L g724 ( .A(n_362), .Y(n_724) );
BUFx2_ASAP7_75t_L g1188 ( .A(n_363), .Y(n_1188) );
INVx1_ASAP7_75t_L g853 ( .A(n_364), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_366), .Y(n_1211) );
OR2x6_ASAP7_75t_SL g366 ( .A(n_367), .B(n_370), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g374 ( .A(n_368), .B(n_375), .Y(n_374) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_368), .Y(n_642) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g399 ( .A(n_369), .Y(n_399) );
OR2x2_ASAP7_75t_L g526 ( .A(n_369), .B(n_495), .Y(n_526) );
INVx3_ASAP7_75t_L g810 ( .A(n_370), .Y(n_810) );
BUFx2_ASAP7_75t_L g1022 ( .A(n_370), .Y(n_1022) );
BUFx2_ASAP7_75t_L g1538 ( .A(n_370), .Y(n_1538) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_371), .Y(n_382) );
BUFx8_ASAP7_75t_L g529 ( .A(n_371), .Y(n_529) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_371), .Y(n_624) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_374), .B(n_655), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_374), .A2(n_1210), .B1(n_1211), .B2(n_1212), .Y(n_1209) );
BUFx3_ASAP7_75t_L g395 ( .A(n_375), .Y(n_395) );
BUFx12f_ASAP7_75t_L g412 ( .A(n_375), .Y(n_412) );
INVx5_ASAP7_75t_L g539 ( .A(n_375), .Y(n_539) );
BUFx2_ASAP7_75t_L g619 ( .A(n_375), .Y(n_619) );
BUFx3_ASAP7_75t_L g844 ( .A(n_375), .Y(n_844) );
NOR3xp33_ASAP7_75t_L g376 ( .A(n_377), .B(n_396), .C(n_403), .Y(n_376) );
NOR3xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_383), .C(n_394), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_379), .B(n_460), .Y(n_471) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g1113 ( .A(n_381), .Y(n_1113) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g877 ( .A(n_382), .Y(n_877) );
INVx2_ASAP7_75t_L g945 ( .A(n_382), .Y(n_945) );
INVx1_ASAP7_75t_L g964 ( .A(n_382), .Y(n_964) );
AND2x4_ASAP7_75t_L g1174 ( .A(n_382), .B(n_1175), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g1119 ( .A1(n_386), .A2(n_865), .B1(n_1120), .B2(n_1121), .Y(n_1119) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g558 ( .A(n_387), .B(n_526), .Y(n_558) );
INVx3_ASAP7_75t_L g717 ( .A(n_387), .Y(n_717) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_387), .Y(n_823) );
INVx4_ASAP7_75t_L g864 ( .A(n_387), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_389), .A2(n_621), .B1(n_703), .B2(n_709), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g815 ( .A1(n_389), .A2(n_516), .B(n_780), .C(n_816), .Y(n_815) );
INVx8_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g524 ( .A(n_390), .Y(n_524) );
INVx2_ASAP7_75t_L g534 ( .A(n_390), .Y(n_534) );
INVx3_ASAP7_75t_L g851 ( .A(n_390), .Y(n_851) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g873 ( .A1(n_392), .A2(n_874), .B1(n_875), .B2(n_876), .C(n_878), .Y(n_873) );
OAI221xp5_ASAP7_75t_L g967 ( .A1(n_392), .A2(n_539), .B1(n_617), .B2(n_968), .C(n_969), .Y(n_967) );
OAI221xp5_ASAP7_75t_L g1074 ( .A1(n_392), .A2(n_823), .B1(n_942), .B2(n_1075), .C(n_1076), .Y(n_1074) );
OAI221xp5_ASAP7_75t_L g1261 ( .A1(n_392), .A2(n_623), .B1(n_724), .B2(n_1262), .C(n_1263), .Y(n_1261) );
OAI221xp5_ASAP7_75t_L g1617 ( .A1(n_392), .A2(n_1266), .B1(n_1598), .B2(n_1614), .C(n_1618), .Y(n_1617) );
INVx3_ASAP7_75t_L g1184 ( .A(n_393), .Y(n_1184) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g1066 ( .A1(n_398), .A2(n_401), .B1(n_1067), .B2(n_1068), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_398), .A2(n_401), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
AND2x2_ASAP7_75t_L g401 ( .A(n_399), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g536 ( .A(n_402), .Y(n_536) );
BUFx2_ASAP7_75t_L g549 ( .A(n_402), .Y(n_549) );
BUFx2_ASAP7_75t_L g621 ( .A(n_402), .Y(n_621) );
BUFx3_ASAP7_75t_L g631 ( .A(n_402), .Y(n_631) );
BUFx2_ASAP7_75t_L g652 ( .A(n_402), .Y(n_652) );
BUFx2_ASAP7_75t_L g1222 ( .A(n_402), .Y(n_1222) );
BUFx2_ASAP7_75t_L g1543 ( .A(n_402), .Y(n_1543) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g1081 ( .A1(n_407), .A2(n_413), .B1(n_875), .B2(n_1082), .C(n_1083), .Y(n_1081) );
BUFx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx4f_ASAP7_75t_L g728 ( .A(n_408), .Y(n_728) );
BUFx3_ASAP7_75t_L g865 ( .A(n_408), .Y(n_865) );
INVx2_ASAP7_75t_L g871 ( .A(n_408), .Y(n_871) );
OR2x4_ASAP7_75t_L g1192 ( .A(n_408), .B(n_1175), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_412), .Y(n_1031) );
INVx3_ASAP7_75t_L g634 ( .A(n_413), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_413), .A2(n_722), .B1(n_725), .B2(n_726), .C(n_729), .Y(n_721) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_413), .A2(n_862), .B1(n_863), .B2(n_865), .C(n_866), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_413), .B(n_976), .Y(n_975) );
OAI221xp5_ASAP7_75t_L g1267 ( .A1(n_413), .A2(n_724), .B1(n_728), .B2(n_1268), .C(n_1269), .Y(n_1267) );
OAI221xp5_ASAP7_75t_L g1612 ( .A1(n_413), .A2(n_726), .B1(n_1613), .B2(n_1614), .C(n_1615), .Y(n_1612) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g836 ( .A(n_414), .B(n_468), .Y(n_836) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g608 ( .A(n_417), .Y(n_608) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g929 ( .A1(n_418), .A2(n_930), .B1(n_949), .B2(n_951), .Y(n_929) );
INVx2_ASAP7_75t_SL g977 ( .A(n_418), .Y(n_977) );
OAI31xp33_ASAP7_75t_SL g1064 ( .A1(n_418), .A2(n_1065), .A3(n_1069), .B(n_1073), .Y(n_1064) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_419), .B(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g468 ( .A(n_419), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_422), .Y(n_666) );
INVx1_ASAP7_75t_L g950 ( .A(n_422), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_422), .B(n_979), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_422), .B(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1252 ( .A(n_422), .Y(n_1252) );
INVx2_ASAP7_75t_L g474 ( .A(n_424), .Y(n_474) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_424), .Y(n_603) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx3_ASAP7_75t_L g487 ( .A(n_425), .Y(n_487) );
INVx2_ASAP7_75t_L g670 ( .A(n_425), .Y(n_670) );
AND2x4_ASAP7_75t_L g1139 ( .A(n_425), .B(n_1140), .Y(n_1139) );
NAND3xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_454), .C(n_497), .Y(n_427) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g662 ( .A(n_431), .Y(n_662) );
INVx1_ASAP7_75t_L g702 ( .A(n_431), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_431), .A2(n_912), .B1(n_913), .B2(n_914), .Y(n_911) );
AOI21xp33_ASAP7_75t_L g1093 ( .A1(n_431), .A2(n_1094), .B(n_1095), .Y(n_1093) );
AOI222xp33_ASAP7_75t_L g1232 ( .A1(n_431), .A2(n_498), .B1(n_914), .B2(n_1212), .C1(n_1215), .C2(n_1233), .Y(n_1232) );
AOI222xp33_ASAP7_75t_L g1277 ( .A1(n_431), .A2(n_439), .B1(n_448), .B2(n_1271), .C1(n_1278), .C2(n_1279), .Y(n_1277) );
AOI222xp33_ASAP7_75t_L g1602 ( .A1(n_431), .A2(n_498), .B1(n_914), .B2(n_1603), .C1(n_1604), .C2(n_1605), .Y(n_1602) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g461 ( .A(n_433), .B(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g663 ( .A(n_433), .B(n_462), .Y(n_663) );
INVx1_ASAP7_75t_L g500 ( .A(n_434), .Y(n_500) );
INVx1_ASAP7_75t_L g546 ( .A(n_434), .Y(n_546) );
INVx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g489 ( .A(n_437), .Y(n_489) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_437), .Y(n_566) );
BUFx3_ASAP7_75t_L g689 ( .A(n_437), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_439), .A2(n_448), .B1(n_709), .B2(n_711), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g919 ( .A1(n_439), .A2(n_448), .B1(n_920), .B2(n_921), .Y(n_919) );
AOI22xp5_ASAP7_75t_L g984 ( .A1(n_439), .A2(n_448), .B1(n_985), .B2(n_986), .Y(n_984) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g896 ( .A(n_440), .Y(n_896) );
HB1xp67_ASAP7_75t_L g1236 ( .A(n_440), .Y(n_1236) );
NAND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_444), .Y(n_440) );
INVx1_ASAP7_75t_L g507 ( .A(n_441), .Y(n_507) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_443), .B(n_451), .Y(n_450) );
AND2x6_ASAP7_75t_L g578 ( .A(n_443), .B(n_457), .Y(n_578) );
INVx1_ASAP7_75t_L g593 ( .A(n_443), .Y(n_593) );
AND2x2_ASAP7_75t_L g788 ( .A(n_443), .B(n_789), .Y(n_788) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g592 ( .A(n_446), .Y(n_592) );
BUFx2_ASAP7_75t_L g789 ( .A(n_446), .Y(n_789) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_446), .B(n_1150), .Y(n_1159) );
INVx2_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g557 ( .A(n_449), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g791 ( .A(n_450), .Y(n_791) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_470), .B1(n_484), .B2(n_488), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_456), .A2(n_489), .B1(n_780), .B2(n_781), .Y(n_779) );
A2O1A1Ixp33_ASAP7_75t_L g784 ( .A1(n_456), .A2(n_757), .B(n_785), .C(n_786), .Y(n_784) );
BUFx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g485 ( .A(n_457), .Y(n_485) );
BUFx3_ASAP7_75t_L g671 ( .A(n_457), .Y(n_671) );
BUFx6f_ASAP7_75t_L g998 ( .A(n_457), .Y(n_998) );
BUFx3_ASAP7_75t_L g1050 ( .A(n_457), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_457), .B(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1284 ( .A(n_457), .Y(n_1284) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g573 ( .A(n_458), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_459), .A2(n_471), .B1(n_472), .B2(n_475), .Y(n_470) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g914 ( .A(n_461), .Y(n_914) );
BUFx3_ASAP7_75t_L g887 ( .A(n_462), .Y(n_887) );
INVx2_ASAP7_75t_SL g1131 ( .A(n_462), .Y(n_1131) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_463), .Y(n_506) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g741 ( .A(n_466), .Y(n_741) );
INVx4_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g691 ( .A(n_467), .Y(n_691) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_467), .Y(n_882) );
AOI31xp33_ASAP7_75t_L g916 ( .A1(n_467), .A2(n_504), .A3(n_917), .B(n_918), .Y(n_916) );
INVx2_ASAP7_75t_L g994 ( .A(n_467), .Y(n_994) );
INVx1_ASAP7_75t_L g1123 ( .A(n_467), .Y(n_1123) );
AOI222xp33_ASAP7_75t_L g1280 ( .A1(n_467), .A2(n_498), .B1(n_676), .B2(n_1281), .C1(n_1282), .C2(n_1291), .Y(n_1280) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g655 ( .A(n_468), .Y(n_655) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g575 ( .A(n_473), .Y(n_575) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_478), .B2(n_479), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_477), .A2(n_479), .B1(n_969), .B2(n_992), .Y(n_991) );
INVx5_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx6_ASAP7_75t_L g599 ( .A(n_480), .Y(n_599) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g1002 ( .A(n_481), .Y(n_1002) );
INVx1_ASAP7_75t_L g1135 ( .A(n_481), .Y(n_1135) );
INVx4_ASAP7_75t_L g1290 ( .A(n_481), .Y(n_1290) );
INVx2_ASAP7_75t_SL g1297 ( .A(n_481), .Y(n_1297) );
INVx1_ASAP7_75t_L g1569 ( .A(n_481), .Y(n_1569) );
INVx2_ASAP7_75t_L g1601 ( .A(n_481), .Y(n_1601) );
INVx8_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_482), .B(n_1150), .Y(n_1149) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g1240 ( .A(n_487), .Y(n_1240) );
INVx1_ASAP7_75t_L g1286 ( .A(n_487), .Y(n_1286) );
BUFx3_ASAP7_75t_L g1044 ( .A(n_489), .Y(n_1044) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g748 ( .A(n_491), .Y(n_748) );
INVx2_ASAP7_75t_L g893 ( .A(n_491), .Y(n_893) );
INVx2_ASAP7_75t_L g1043 ( .A(n_491), .Y(n_1043) );
INVx1_ASAP7_75t_L g1048 ( .A(n_491), .Y(n_1048) );
INVx1_ASAP7_75t_L g1242 ( .A(n_492), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .Y(n_492) );
AND2x4_ASAP7_75t_L g676 ( .A(n_493), .B(n_496), .Y(n_676) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g819 ( .A(n_495), .B(n_626), .Y(n_819) );
HB1xp67_ASAP7_75t_L g1200 ( .A(n_495), .Y(n_1200) );
INVx4_ASAP7_75t_L g576 ( .A(n_496), .Y(n_576) );
INVx4_ASAP7_75t_L g801 ( .A(n_496), .Y(n_801) );
INVx1_ASAP7_75t_SL g1559 ( .A(n_496), .Y(n_1559) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_503), .B(n_504), .Y(n_497) );
AOI322xp5_ASAP7_75t_L g988 ( .A1(n_498), .A2(n_676), .A3(n_989), .B1(n_990), .B2(n_993), .C1(n_995), .C2(n_996), .Y(n_988) );
AOI332xp33_ASAP7_75t_L g1096 ( .A1(n_498), .A2(n_676), .A3(n_741), .B1(n_1097), .B2(n_1098), .B3(n_1099), .C1(n_1100), .C2(n_1101), .Y(n_1096) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g556 ( .A(n_500), .B(n_502), .Y(n_556) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g1090 ( .A1(n_504), .A2(n_914), .B(n_1072), .Y(n_1090) );
AOI21xp5_ASAP7_75t_L g1300 ( .A1(n_504), .A2(n_914), .B(n_1301), .Y(n_1300) );
NOR3xp33_ASAP7_75t_L g1585 ( .A(n_504), .B(n_1586), .C(n_1587), .Y(n_1585) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g677 ( .A1(n_505), .A2(n_678), .B(n_690), .Y(n_677) );
OAI21xp5_ASAP7_75t_SL g738 ( .A1(n_505), .A2(n_739), .B(n_742), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g888 ( .A1(n_505), .A2(n_759), .B(n_889), .Y(n_888) );
OAI21xp5_ASAP7_75t_L g1244 ( .A1(n_505), .A2(n_1245), .B(n_1247), .Y(n_1244) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx4_ASAP7_75t_L g685 ( .A(n_506), .Y(n_685) );
BUFx4f_ASAP7_75t_L g746 ( .A(n_506), .Y(n_746) );
BUFx4f_ASAP7_75t_L g755 ( .A(n_506), .Y(n_755) );
BUFx4f_ASAP7_75t_L g1154 ( .A(n_506), .Y(n_1154) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_562), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_550), .C(n_561), .Y(n_511) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_521), .C(n_530), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_517), .B2(n_518), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_515), .A2(n_518), .B1(n_1016), .B2(n_1017), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1531 ( .A1(n_515), .A2(n_518), .B1(n_1532), .B2(n_1533), .Y(n_1531) );
AND2x4_ASAP7_75t_L g518 ( .A(n_516), .B(n_519), .Y(n_518) );
AND2x4_ASAP7_75t_L g561 ( .A(n_516), .B(n_549), .Y(n_561) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_527), .B2(n_528), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_522), .A2(n_527), .B1(n_580), .B2(n_582), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_523), .B(n_806), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_523), .A2(n_528), .B1(n_1035), .B2(n_1038), .Y(n_1056) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
AND2x4_ASAP7_75t_L g528 ( .A(n_525), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g552 ( .A(n_526), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g811 ( .A(n_526), .Y(n_811) );
INVx2_ASAP7_75t_L g1548 ( .A(n_528), .Y(n_1548) );
INVx3_ASAP7_75t_L g542 ( .A(n_529), .Y(n_542) );
INVx2_ASAP7_75t_SL g731 ( .A(n_529), .Y(n_731) );
INVx3_ASAP7_75t_L g942 ( .A(n_529), .Y(n_942) );
INVx2_ASAP7_75t_SL g1266 ( .A(n_529), .Y(n_1266) );
AOI33xp33_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_533), .A3(n_537), .B1(n_540), .B2(n_544), .B3(n_547), .Y(n_530) );
INVx1_ASAP7_75t_L g1029 ( .A(n_531), .Y(n_1029) );
AOI33xp33_ASAP7_75t_L g1534 ( .A1(n_531), .A2(n_1535), .A3(n_1536), .B1(n_1539), .B2(n_1540), .B3(n_1542), .Y(n_1534) );
BUFx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_534), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g846 ( .A(n_536), .Y(n_846) );
INVx2_ASAP7_75t_L g1023 ( .A(n_536), .Y(n_1023) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g543 ( .A(n_539), .Y(n_543) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g1118 ( .A(n_544), .Y(n_1118) );
CKINVDCx5p33_ASAP7_75t_R g1541 ( .A(n_544), .Y(n_1541) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx3_ASAP7_75t_L g1026 ( .A(n_545), .Y(n_1026) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_549), .A2(n_851), .B1(n_908), .B2(n_921), .Y(n_946) );
INVx8_ASAP7_75t_L g1012 ( .A(n_551), .Y(n_1012) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_556), .Y(n_551) );
INVx1_ASAP7_75t_L g1088 ( .A(n_553), .Y(n_1088) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_554), .Y(n_734) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g648 ( .A(n_555), .Y(n_648) );
INVx1_ASAP7_75t_L g661 ( .A(n_556), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_556), .B(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g812 ( .A(n_558), .Y(n_812) );
INVx3_ASAP7_75t_L g1010 ( .A(n_559), .Y(n_1010) );
INVx3_ASAP7_75t_L g1018 ( .A(n_561), .Y(n_1018) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_585), .B(n_606), .Y(n_562) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g1040 ( .A1(n_565), .A2(n_578), .B1(n_1011), .B2(n_1041), .C(n_1042), .Y(n_1040) );
BUFx2_ASAP7_75t_L g749 ( .A(n_566), .Y(n_749) );
INVx1_ASAP7_75t_L g925 ( .A(n_566), .Y(n_925) );
AOI21xp5_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_577), .B(n_578), .Y(n_567) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g928 ( .A(n_572), .Y(n_928) );
INVx1_ASAP7_75t_L g1241 ( .A(n_572), .Y(n_1241) );
BUFx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g1555 ( .A1(n_578), .A2(n_1556), .B(n_1560), .Y(n_1555) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g1561 ( .A1(n_582), .A2(n_1036), .B1(n_1562), .B2(n_1563), .Y(n_1561) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx6f_ASAP7_75t_L g1039 ( .A(n_584), .Y(n_1039) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g1565 ( .A(n_587), .Y(n_1565) );
INVx4_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx3_ASAP7_75t_L g1046 ( .A(n_589), .Y(n_1046) );
BUFx2_ASAP7_75t_L g1566 ( .A(n_590), .Y(n_1566) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2x1_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g786 ( .A(n_593), .Y(n_786) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_598), .B1(n_599), .B2(n_600), .C(n_601), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g1567 ( .A1(n_595), .A2(n_1568), .B1(n_1569), .B2(n_1570), .C(n_1571), .Y(n_1567) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g1125 ( .A(n_596), .Y(n_1125) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx3_ASAP7_75t_L g674 ( .A(n_597), .Y(n_674) );
INVx4_ASAP7_75t_L g1289 ( .A(n_597), .Y(n_1289) );
OAI22xp33_ASAP7_75t_L g672 ( .A1(n_599), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g889 ( .A1(n_599), .A2(n_859), .B1(n_874), .B2(n_890), .C(n_892), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_599), .A2(n_1109), .B1(n_1120), .B2(n_1125), .Y(n_1124) );
BUFx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx3_ASAP7_75t_L g798 ( .A(n_605), .Y(n_798) );
INVx1_ASAP7_75t_L g1051 ( .A(n_605), .Y(n_1051) );
OAI21xp5_ASAP7_75t_L g1553 ( .A1(n_606), .A2(n_1554), .B(n_1564), .Y(n_1553) );
A2O1A1Ixp33_ASAP7_75t_SL g1606 ( .A1(n_606), .A2(n_1607), .B(n_1610), .C(n_1620), .Y(n_1606) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g736 ( .A(n_608), .Y(n_736) );
INVx2_ASAP7_75t_SL g766 ( .A(n_609), .Y(n_766) );
XNOR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_695), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_693), .B(n_694), .Y(n_610) );
AND3x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_658), .C(n_667), .Y(n_611) );
AOI31xp33_ASAP7_75t_L g694 ( .A1(n_612), .A2(n_658), .A3(n_667), .B(n_693), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_654), .B(n_656), .Y(n_612) );
NAND3xp33_ASAP7_75t_SL g613 ( .A(n_614), .B(n_635), .C(n_639), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_620), .B1(n_627), .B2(n_630), .Y(n_614) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_SL g629 ( .A(n_624), .Y(n_629) );
INVx3_ASAP7_75t_L g644 ( .A(n_624), .Y(n_644) );
INVx5_ASAP7_75t_L g826 ( .A(n_624), .Y(n_826) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_624), .Y(n_858) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g1224 ( .A(n_633), .Y(n_1224) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_638), .B(n_932), .Y(n_931) );
INVxp67_ASAP7_75t_L g707 ( .A(n_640), .Y(n_707) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx2_ASAP7_75t_L g842 ( .A(n_642), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_645), .A2(n_868), .B1(n_869), .B2(n_872), .Y(n_867) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g827 ( .A(n_647), .Y(n_827) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx3_ASAP7_75t_L g860 ( .A(n_648), .Y(n_860) );
INVx2_ASAP7_75t_L g1054 ( .A(n_654), .Y(n_1054) );
OAI21xp5_ASAP7_75t_L g1207 ( .A1(n_654), .A2(n_1208), .B(n_1216), .Y(n_1207) );
BUFx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI21xp5_ASAP7_75t_SL g775 ( .A1(n_655), .A2(n_776), .B(n_793), .Y(n_775) );
INVx1_ASAP7_75t_L g880 ( .A(n_655), .Y(n_880) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_664), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g1620 ( .A(n_666), .B(n_1621), .Y(n_1620) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_676), .B(n_677), .C(n_692), .Y(n_667) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g797 ( .A(n_670), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_676), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g922 ( .A(n_676), .B(n_923), .C(n_926), .Y(n_922) );
INVx2_ASAP7_75t_L g1132 ( .A(n_676), .Y(n_1132) );
OAI221xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_683), .B1(n_684), .B2(n_686), .C(n_687), .Y(n_678) );
OAI221xp5_ASAP7_75t_L g1596 ( .A1(n_679), .A2(n_746), .B1(n_1597), .B2(n_1598), .C(n_1599), .Y(n_1596) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
BUFx3_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g744 ( .A(n_682), .Y(n_744) );
BUFx2_ASAP7_75t_L g754 ( .A(n_682), .Y(n_754) );
INVx1_ASAP7_75t_L g891 ( .A(n_682), .Y(n_891) );
OAI221xp5_ASAP7_75t_L g1247 ( .A1(n_684), .A2(n_752), .B1(n_1218), .B2(n_1248), .C(n_1249), .Y(n_1247) );
INVx1_ASAP7_75t_L g1593 ( .A(n_684), .Y(n_1593) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx3_ASAP7_75t_L g758 ( .A(n_688), .Y(n_758) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_688), .Y(n_803) );
INVx1_ASAP7_75t_L g1246 ( .A(n_690), .Y(n_1246) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_705), .C(n_737), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_720), .B(n_736), .Y(n_705) );
OAI211xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B(n_710), .C(n_713), .Y(n_706) );
OAI211xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B(n_718), .C(n_719), .Y(n_713) );
OAI221xp5_ASAP7_75t_L g751 ( .A1(n_714), .A2(n_725), .B1(n_752), .B2(n_755), .C(n_756), .Y(n_751) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI211xp5_ASAP7_75t_L g1225 ( .A1(n_716), .A2(n_1226), .B(n_1227), .C(n_1228), .Y(n_1225) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g1108 ( .A1(n_722), .A2(n_865), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI22xp33_ASAP7_75t_L g833 ( .A1(n_724), .A2(n_728), .B1(n_834), .B2(n_835), .Y(n_833) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI22xp33_ASAP7_75t_L g820 ( .A1(n_728), .A2(n_821), .B1(n_822), .B2(n_823), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_733), .B2(n_735), .Y(n_730) );
OAI221xp5_ASAP7_75t_L g742 ( .A1(n_732), .A2(n_743), .B1(n_745), .B2(n_746), .C(n_747), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_733), .A2(n_1112), .B1(n_1113), .B2(n_1114), .Y(n_1111) );
CKINVDCx8_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
INVx3_ASAP7_75t_L g1080 ( .A(n_734), .Y(n_1080) );
INVx3_ASAP7_75t_L g1219 ( .A(n_734), .Y(n_1219) );
NOR3xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_750), .C(n_761), .Y(n_737) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_743), .A2(n_746), .B1(n_1112), .B2(n_1116), .Y(n_1126) );
INVx1_ASAP7_75t_L g1129 ( .A(n_743), .Y(n_1129) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g778 ( .A(n_753), .Y(n_778) );
INVx4_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
XNOR2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_902), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
XNOR2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_837), .Y(n_770) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_804), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_782), .B(n_783), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_787), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_788), .A2(n_790), .B1(n_791), .B2(n_792), .Y(n_787) );
INVx1_ASAP7_75t_L g1053 ( .A(n_788), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_792), .A2(n_808), .B1(n_809), .B2(n_812), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_799), .B1(n_800), .B2(n_802), .Y(n_793) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g927 ( .A(n_796), .Y(n_927) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NAND3xp33_ASAP7_75t_SL g804 ( .A(n_805), .B(n_807), .C(n_813), .Y(n_804) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx2_ASAP7_75t_L g830 ( .A(n_810), .Y(n_830) );
INVxp67_ASAP7_75t_L g1547 ( .A(n_811), .Y(n_1547) );
NOR2xp33_ASAP7_75t_SL g813 ( .A(n_814), .B(n_817), .Y(n_813) );
OAI33xp33_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_820), .A3(n_824), .B1(n_829), .B2(n_833), .B3(n_836), .Y(n_817) );
BUFx4f_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
BUFx8_ASAP7_75t_L g1107 ( .A(n_819), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_826), .B1(n_827), .B2(n_828), .Y(n_824) );
INVx8_ASAP7_75t_L g938 ( .A(n_826), .Y(n_938) );
OAI221xp5_ASAP7_75t_L g1217 ( .A1(n_826), .A2(n_1218), .B1(n_1219), .B2(n_1220), .C(n_1221), .Y(n_1217) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_827), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_830), .A2(n_860), .B1(n_1116), .B2(n_1117), .Y(n_1115) );
NAND4xp75_ASAP7_75t_L g838 ( .A(n_839), .B(n_881), .C(n_898), .D(n_899), .Y(n_838) );
OAI21x1_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_854), .B(n_879), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_843), .B(n_849), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_842), .A2(n_912), .B1(n_944), .B2(n_947), .Y(n_943) );
AOI221xp5_ASAP7_75t_SL g843 ( .A1(n_844), .A2(n_845), .B1(n_846), .B2(n_847), .C(n_848), .Y(n_843) );
A2O1A1Ixp33_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_851), .B(n_852), .C(n_853), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_861), .B1(n_867), .B2(n_873), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_857), .B1(n_859), .B2(n_860), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_856), .A2(n_868), .B1(n_885), .B2(n_887), .Y(n_884) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g875 ( .A(n_864), .Y(n_875) );
INVx2_ASAP7_75t_L g966 ( .A(n_864), .Y(n_966) );
INVx2_ASAP7_75t_L g1614 ( .A(n_864), .Y(n_1614) );
BUFx4f_ASAP7_75t_SL g869 ( .A(n_870), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_870), .A2(n_1078), .B1(n_1079), .B2(n_1080), .Y(n_1077) );
INVx3_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx2_ASAP7_75t_SL g1546 ( .A(n_871), .Y(n_1546) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
AOI211x1_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_883), .B(n_888), .C(n_894), .Y(n_881) );
BUFx3_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
BUFx3_ASAP7_75t_L g1000 ( .A(n_886), .Y(n_1000) );
BUFx6f_ASAP7_75t_L g1595 ( .A(n_886), .Y(n_1595) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_953), .B1(n_954), .B2(n_1003), .Y(n_902) );
INVx1_ASAP7_75t_L g1003 ( .A(n_903), .Y(n_1003) );
OAI21x1_ASAP7_75t_SL g903 ( .A1(n_904), .A2(n_905), .B(n_952), .Y(n_903) );
NAND4xp25_ASAP7_75t_L g952 ( .A(n_904), .B(n_907), .C(n_909), .D(n_929), .Y(n_952) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
NAND3xp33_ASAP7_75t_L g906 ( .A(n_907), .B(n_909), .C(n_929), .Y(n_906) );
NOR2xp33_ASAP7_75t_L g909 ( .A(n_910), .B(n_915), .Y(n_909) );
NAND3xp33_ASAP7_75t_SL g915 ( .A(n_916), .B(n_919), .C(n_922), .Y(n_915) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
NAND3xp33_ASAP7_75t_L g930 ( .A(n_931), .B(n_935), .C(n_943), .Y(n_930) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B1(n_939), .B2(n_940), .Y(n_935) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_942), .A2(n_1085), .B1(n_1086), .B2(n_1087), .Y(n_1084) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_949), .B(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx2_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
NOR2x1_ASAP7_75t_L g955 ( .A(n_956), .B(n_980), .Y(n_955) );
A2O1A1Ixp33_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_961), .B(n_977), .C(n_978), .Y(n_956) );
NOR3xp33_ASAP7_75t_SL g961 ( .A(n_962), .B(n_970), .C(n_971), .Y(n_961) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_968), .A2(n_1000), .B1(n_1001), .B2(n_1002), .Y(n_999) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_988), .Y(n_980) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
BUFx2_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1558 ( .A(n_998), .Y(n_1558) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
NAND2xp67_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1032), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g1009 ( .A1(n_1010), .A2(n_1011), .B1(n_1012), .B2(n_1013), .C(n_1014), .Y(n_1009) );
AOI21xp5_ASAP7_75t_L g1550 ( .A1(n_1012), .A2(n_1551), .B(n_1552), .Y(n_1550) );
NAND3xp33_ASAP7_75t_SL g1014 ( .A(n_1015), .B(n_1018), .C(n_1019), .Y(n_1014) );
AOI222xp33_ASAP7_75t_L g1045 ( .A1(n_1016), .A2(n_1017), .B1(n_1046), .B2(n_1047), .C1(n_1049), .C2(n_1052), .Y(n_1045) );
INVx2_ASAP7_75t_SL g1549 ( .A(n_1018), .Y(n_1549) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1024), .B1(n_1028), .B2(n_1030), .Y(n_1019) );
INVx2_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1027), .Y(n_1024) );
BUFx2_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
AOI21xp5_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1054), .B(n_1055), .Y(n_1032) );
NAND3xp33_ASAP7_75t_SL g1033 ( .A(n_1034), .B(n_1040), .C(n_1045), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1036), .B1(n_1038), .B2(n_1039), .Y(n_1034) );
HB1xp67_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
A2O1A1Ixp33_ASAP7_75t_L g1257 ( .A1(n_1054), .A2(n_1258), .B(n_1270), .C(n_1274), .Y(n_1257) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g1058 ( .A1(n_1059), .A2(n_1203), .B1(n_1302), .B2(n_1303), .Y(n_1058) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1059), .Y(n_1302) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_1060), .A2(n_1061), .B1(n_1103), .B2(n_1202), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
XOR2x2_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1102), .Y(n_1061) );
NOR2xp33_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1089), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_1074), .A2(n_1077), .B1(n_1081), .B2(n_1084), .Y(n_1073) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
NAND4xp25_ASAP7_75t_SL g1089 ( .A(n_1090), .B(n_1091), .C(n_1093), .D(n_1096), .Y(n_1089) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1103), .Y(n_1202) );
XOR2x2_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1201), .Y(n_1103) );
AND3x1_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1136), .C(n_1168), .Y(n_1104) );
NOR2xp33_ASAP7_75t_SL g1105 ( .A(n_1106), .B(n_1122), .Y(n_1105) );
OAI33xp33_ASAP7_75t_L g1106 ( .A1(n_1107), .A2(n_1108), .A3(n_1111), .B1(n_1115), .B2(n_1118), .B3(n_1119), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1127 ( .A1(n_1110), .A2(n_1121), .B1(n_1128), .B2(n_1130), .Y(n_1127) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_1114), .A2(n_1117), .B1(n_1125), .B2(n_1134), .Y(n_1133) );
OAI33xp33_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1124), .A3(n_1126), .B1(n_1127), .B2(n_1132), .B3(n_1133), .Y(n_1122) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
INVx5_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
BUFx3_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
OAI31xp33_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1141), .A3(n_1151), .B(n_1165), .Y(n_1136) );
INVx4_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx2_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx3_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_1159), .A2(n_1160), .B1(n_1161), .B2(n_1164), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_1160), .A2(n_1182), .B1(n_1186), .B2(n_1189), .Y(n_1181) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
BUFx3_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
OAI31xp33_ASAP7_75t_L g1168 ( .A1(n_1169), .A2(n_1176), .A3(n_1190), .B(n_1196), .Y(n_1168) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx2_ASAP7_75t_SL g1171 ( .A(n_1172), .Y(n_1171) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVxp67_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
CKINVDCx8_ASAP7_75t_R g1179 ( .A(n_1180), .Y(n_1179) );
BUFx3_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1185), .Y(n_1183) );
AND2x4_ASAP7_75t_L g1187 ( .A(n_1184), .B(n_1188), .Y(n_1187) );
BUFx6f_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
BUFx2_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
AND2x2_ASAP7_75t_SL g1196 ( .A(n_1197), .B(n_1199), .Y(n_1196) );
INVx1_ASAP7_75t_SL g1197 ( .A(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1203), .Y(n_1303) );
XOR2x2_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1255), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1206), .Y(n_1253) );
NAND4xp25_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1232), .C(n_1234), .D(n_1250), .Y(n_1206) );
NAND3xp33_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1225), .C(n_1229), .Y(n_1216) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1244), .Y(n_1234) );
NAND3xp33_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1242), .C(n_1243), .Y(n_1237) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
OAI221xp5_ASAP7_75t_L g1363 ( .A1(n_1254), .A2(n_1364), .B1(n_1365), .B2(n_1366), .C(n_1367), .Y(n_1363) );
OR2x2_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1276), .Y(n_1256) );
NOR3xp33_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1260), .C(n_1264), .Y(n_1258) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
OAI22xp5_ASAP7_75t_L g1287 ( .A1(n_1269), .A2(n_1288), .B1(n_1289), .B2(n_1290), .Y(n_1287) );
NAND4xp25_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1280), .C(n_1298), .D(n_1300), .Y(n_1276) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
HB1xp67_ASAP7_75t_L g1590 ( .A(n_1290), .Y(n_1590) );
OAI22xp5_ASAP7_75t_L g1292 ( .A1(n_1293), .A2(n_1294), .B1(n_1296), .B2(n_1297), .Y(n_1292) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
OAI221xp5_ASAP7_75t_L g1304 ( .A1(n_1305), .A2(n_1522), .B1(n_1525), .B2(n_1572), .C(n_1578), .Y(n_1304) );
AND3x1_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1451), .C(n_1487), .Y(n_1305) );
NOR3xp33_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1382), .C(n_1440), .Y(n_1306) );
OAI221xp5_ASAP7_75t_L g1307 ( .A1(n_1308), .A2(n_1310), .B1(n_1360), .B2(n_1372), .C(n_1375), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g1308 ( .A1(n_1309), .A2(n_1335), .B1(n_1341), .B2(n_1350), .C(n_1354), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1326), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1311), .B(n_1400), .Y(n_1399) );
CKINVDCx5p33_ASAP7_75t_R g1435 ( .A(n_1311), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1311), .B(n_1454), .Y(n_1453) );
OAI211xp5_ASAP7_75t_SL g1488 ( .A1(n_1311), .A2(n_1489), .B(n_1492), .C(n_1504), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1501 ( .A(n_1311), .B(n_1386), .Y(n_1501) );
NOR2xp33_ASAP7_75t_L g1519 ( .A(n_1311), .B(n_1520), .Y(n_1519) );
INVx4_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx4_ASAP7_75t_L g1343 ( .A(n_1312), .Y(n_1343) );
NAND2xp5_ASAP7_75t_SL g1358 ( .A(n_1312), .B(n_1359), .Y(n_1358) );
OR2x2_ASAP7_75t_L g1390 ( .A(n_1312), .B(n_1359), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1312), .B(n_1443), .Y(n_1442) );
NOR2xp33_ASAP7_75t_L g1450 ( .A(n_1312), .B(n_1374), .Y(n_1450) );
NAND2xp5_ASAP7_75t_L g1497 ( .A(n_1312), .B(n_1410), .Y(n_1497) );
AND2x4_ASAP7_75t_SL g1312 ( .A(n_1313), .B(n_1321), .Y(n_1312) );
AND2x4_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1316), .Y(n_1314) );
AND2x6_ASAP7_75t_L g1319 ( .A(n_1315), .B(n_1320), .Y(n_1319) );
AND2x6_ASAP7_75t_L g1322 ( .A(n_1315), .B(n_1323), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1315), .B(n_1325), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1315), .B(n_1325), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_1315), .B(n_1316), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1315), .B(n_1325), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1318), .Y(n_1316) );
INVx2_ASAP7_75t_L g1366 ( .A(n_1319), .Y(n_1366) );
INVx2_ASAP7_75t_L g1524 ( .A(n_1322), .Y(n_1524) );
OAI21xp5_ASAP7_75t_L g1629 ( .A1(n_1323), .A2(n_1630), .B(n_1631), .Y(n_1629) );
INVxp67_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
NOR2xp33_ASAP7_75t_L g1485 ( .A(n_1327), .B(n_1343), .Y(n_1485) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1332), .Y(n_1327) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1328), .Y(n_1357) );
OR2x2_ASAP7_75t_L g1391 ( .A(n_1328), .B(n_1351), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1328), .B(n_1359), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1328), .B(n_1350), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1328), .B(n_1351), .Y(n_1414) );
NOR2xp33_ASAP7_75t_L g1496 ( .A(n_1328), .B(n_1497), .Y(n_1496) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1328), .Y(n_1507) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1331), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1381 ( .A(n_1332), .B(n_1356), .Y(n_1381) );
OR2x2_ASAP7_75t_L g1412 ( .A(n_1332), .B(n_1413), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_1332), .B(n_1408), .Y(n_1432) );
AOI222xp33_ASAP7_75t_L g1518 ( .A1(n_1332), .A2(n_1454), .B1(n_1460), .B2(n_1468), .C1(n_1519), .C2(n_1521), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1334), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1333), .B(n_1334), .Y(n_1359) );
OAI321xp33_ASAP7_75t_L g1440 ( .A1(n_1335), .A2(n_1441), .A3(n_1444), .B1(n_1445), .B2(n_1446), .C(n_1447), .Y(n_1440) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1336), .B(n_1369), .Y(n_1404) );
NOR2xp33_ASAP7_75t_L g1474 ( .A(n_1336), .B(n_1343), .Y(n_1474) );
NOR2xp33_ASAP7_75t_L g1477 ( .A(n_1336), .B(n_1478), .Y(n_1477) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1337), .B(n_1346), .Y(n_1345) );
OR2x2_ASAP7_75t_L g1374 ( .A(n_1337), .B(n_1347), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1337), .B(n_1377), .Y(n_1392) );
OR2x2_ASAP7_75t_L g1394 ( .A(n_1337), .B(n_1387), .Y(n_1394) );
INVx2_ASAP7_75t_L g1423 ( .A(n_1337), .Y(n_1423) );
OR2x2_ASAP7_75t_L g1431 ( .A(n_1337), .B(n_1369), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1337), .B(n_1369), .Y(n_1499) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
OR2x2_ASAP7_75t_L g1439 ( .A(n_1338), .B(n_1387), .Y(n_1439) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1340), .Y(n_1338) );
NOR2xp33_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1344), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1342), .B(n_1373), .Y(n_1396) );
NAND3xp33_ASAP7_75t_L g1403 ( .A(n_1342), .B(n_1401), .C(n_1404), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1342), .B(n_1346), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1521 ( .A(n_1342), .B(n_1345), .Y(n_1521) );
CKINVDCx5p33_ASAP7_75t_R g1342 ( .A(n_1343), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1343), .B(n_1346), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1343), .B(n_1363), .Y(n_1434) );
NAND2x1_ASAP7_75t_L g1511 ( .A(n_1343), .B(n_1512), .Y(n_1511) );
NOR2xp33_ASAP7_75t_L g1354 ( .A(n_1344), .B(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1345), .B(n_1443), .Y(n_1446) );
INVx2_ASAP7_75t_L g1410 ( .A(n_1346), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_1346), .B(n_1377), .Y(n_1456) );
OAI31xp33_ASAP7_75t_L g1502 ( .A1(n_1346), .A2(n_1351), .A3(n_1395), .B(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1347), .Y(n_1387) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1349), .Y(n_1347) );
NOR2xp33_ASAP7_75t_L g1400 ( .A(n_1350), .B(n_1401), .Y(n_1400) );
OR2x2_ASAP7_75t_L g1449 ( .A(n_1350), .B(n_1359), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1350), .B(n_1359), .Y(n_1483) );
INVx2_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1351), .B(n_1357), .Y(n_1356) );
NAND2x1p5_ASAP7_75t_L g1351 ( .A(n_1352), .B(n_1353), .Y(n_1351) );
OR2x2_ASAP7_75t_L g1355 ( .A(n_1356), .B(n_1358), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1356), .B(n_1407), .Y(n_1406) );
OR2x2_ASAP7_75t_L g1455 ( .A(n_1356), .B(n_1401), .Y(n_1455) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1356), .Y(n_1490) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1358), .Y(n_1419) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1359), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1359), .B(n_1507), .Y(n_1506) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1359), .B(n_1414), .Y(n_1512) );
OR2x2_ASAP7_75t_L g1520 ( .A(n_1359), .B(n_1507), .Y(n_1520) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
NOR2xp33_ASAP7_75t_SL g1361 ( .A(n_1362), .B(n_1369), .Y(n_1361) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1362), .Y(n_1422) );
A2O1A1Ixp33_ASAP7_75t_L g1428 ( .A1(n_1362), .A2(n_1410), .B(n_1429), .C(n_1431), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1362), .B(n_1376), .Y(n_1509) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1369), .Y(n_1373) );
INVx3_ASAP7_75t_L g1377 ( .A(n_1369), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1371), .Y(n_1369) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1372), .Y(n_1491) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1373), .B(n_1374), .Y(n_1372) );
NAND3xp33_ASAP7_75t_L g1503 ( .A(n_1373), .B(n_1380), .C(n_1408), .Y(n_1503) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1378), .Y(n_1375) );
NAND3xp33_ASAP7_75t_L g1500 ( .A(n_1376), .B(n_1408), .C(n_1501), .Y(n_1500) );
CKINVDCx14_ASAP7_75t_R g1376 ( .A(n_1377), .Y(n_1376) );
OR2x2_ASAP7_75t_L g1430 ( .A(n_1377), .B(n_1386), .Y(n_1430) );
OR2x2_ASAP7_75t_L g1438 ( .A(n_1377), .B(n_1439), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1377), .B(n_1460), .Y(n_1459) );
NOR2xp33_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1381), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
NAND3xp33_ASAP7_75t_L g1382 ( .A(n_1383), .B(n_1409), .C(n_1424), .Y(n_1382) );
AOI21xp5_ASAP7_75t_L g1383 ( .A1(n_1384), .A2(n_1392), .B(n_1393), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1385), .B(n_1388), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1416 ( .A(n_1385), .B(n_1417), .Y(n_1416) );
O2A1O1Ixp33_ASAP7_75t_L g1481 ( .A1(n_1385), .A2(n_1482), .B(n_1484), .C(n_1486), .Y(n_1481) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1386), .B(n_1392), .Y(n_1402) );
OAI22xp5_ASAP7_75t_SL g1433 ( .A1(n_1386), .A2(n_1421), .B1(n_1434), .B2(n_1435), .Y(n_1433) );
OAI221xp5_ASAP7_75t_L g1510 ( .A1(n_1386), .A2(n_1511), .B1(n_1513), .B2(n_1514), .C(n_1518), .Y(n_1510) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
AOI222xp33_ASAP7_75t_L g1504 ( .A1(n_1388), .A2(n_1404), .B1(n_1432), .B2(n_1459), .C1(n_1505), .C2(n_1506), .Y(n_1504) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
OR2x2_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1391), .Y(n_1389) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1390), .Y(n_1427) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1391), .Y(n_1418) );
OAI211xp5_ASAP7_75t_SL g1457 ( .A1(n_1391), .A2(n_1458), .B(n_1461), .C(n_1463), .Y(n_1457) );
OR2x2_ASAP7_75t_L g1465 ( .A(n_1391), .B(n_1401), .Y(n_1465) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1392), .Y(n_1486) );
OAI322xp33_ASAP7_75t_L g1393 ( .A1(n_1394), .A2(n_1395), .A3(n_1397), .B1(n_1398), .B2(n_1402), .C1(n_1403), .C2(n_1405), .Y(n_1393) );
CKINVDCx5p33_ASAP7_75t_R g1460 ( .A(n_1394), .Y(n_1460) );
CKINVDCx14_ASAP7_75t_R g1395 ( .A(n_1396), .Y(n_1395) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1397), .Y(n_1479) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1401), .B(n_1418), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1401), .B(n_1408), .Y(n_1443) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1408), .B(n_1427), .Y(n_1467) );
A2O1A1Ixp33_ASAP7_75t_R g1409 ( .A1(n_1410), .A2(n_1411), .B(n_1415), .C(n_1420), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1410), .B(n_1462), .Y(n_1461) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_1410), .B(n_1431), .Y(n_1475) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1410), .Y(n_1513) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
AOI21xp33_ASAP7_75t_SL g1452 ( .A1(n_1412), .A2(n_1453), .B(n_1456), .Y(n_1452) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1414), .B(n_1427), .Y(n_1426) );
AOI211xp5_ASAP7_75t_L g1492 ( .A1(n_1414), .A2(n_1493), .B(n_1494), .C(n_1502), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1414), .B(n_1419), .Y(n_1517) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1419), .Y(n_1417) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1422), .B(n_1423), .Y(n_1421) );
INVx2_ASAP7_75t_L g1445 ( .A(n_1422), .Y(n_1445) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1423), .Y(n_1505) );
AOI222xp33_ASAP7_75t_L g1424 ( .A1(n_1425), .A2(n_1428), .B1(n_1432), .B2(n_1433), .C1(n_1436), .C2(n_1437), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
OAI21xp5_ASAP7_75t_L g1447 ( .A1(n_1432), .A2(n_1448), .B(n_1450), .Y(n_1447) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1432), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1435), .B(n_1436), .Y(n_1462) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1436), .Y(n_1471) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
CKINVDCx5p33_ASAP7_75t_R g1468 ( .A(n_1439), .Y(n_1468) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
AOI22xp5_ASAP7_75t_L g1487 ( .A1(n_1444), .A2(n_1488), .B1(n_1508), .B2(n_1510), .Y(n_1487) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
OAI31xp33_ASAP7_75t_L g1451 ( .A1(n_1445), .A2(n_1452), .A3(n_1457), .B(n_1469), .Y(n_1451) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
OAI221xp5_ASAP7_75t_L g1469 ( .A1(n_1455), .A2(n_1470), .B1(n_1473), .B2(n_1475), .C(n_1476), .Y(n_1469) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
OAI21xp33_ASAP7_75t_L g1463 ( .A1(n_1464), .A2(n_1466), .B(n_1468), .Y(n_1463) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1515 ( .A(n_1465), .B(n_1516), .Y(n_1515) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1472), .Y(n_1470) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1475), .Y(n_1493) );
NOR2xp33_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1481), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1480), .Y(n_1478) );
CKINVDCx14_ASAP7_75t_R g1482 ( .A(n_1483), .Y(n_1482) );
INVxp67_ASAP7_75t_SL g1484 ( .A(n_1485), .Y(n_1484) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1490), .B(n_1491), .Y(n_1489) );
OAI21xp33_ASAP7_75t_L g1494 ( .A1(n_1495), .A2(n_1498), .B(n_1500), .Y(n_1494) );
INVxp33_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
INVxp67_ASAP7_75t_SL g1514 ( .A(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
CKINVDCx20_ASAP7_75t_R g1522 ( .A(n_1523), .Y(n_1522) );
CKINVDCx20_ASAP7_75t_R g1523 ( .A(n_1524), .Y(n_1523) );
INVx2_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
INVx2_ASAP7_75t_SL g1526 ( .A(n_1527), .Y(n_1526) );
NAND3xp33_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1550), .C(n_1553), .Y(n_1528) );
NOR3xp33_ASAP7_75t_L g1529 ( .A(n_1530), .B(n_1544), .C(n_1549), .Y(n_1529) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1534), .Y(n_1530) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
OR2x6_ASAP7_75t_L g1545 ( .A(n_1546), .B(n_1547), .Y(n_1545) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
CKINVDCx20_ASAP7_75t_R g1572 ( .A(n_1573), .Y(n_1572) );
CKINVDCx20_ASAP7_75t_R g1573 ( .A(n_1574), .Y(n_1573) );
INVx3_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
BUFx3_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
CKINVDCx5p33_ASAP7_75t_R g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1582), .Y(n_1624) );
BUFx4_ASAP7_75t_R g1582 ( .A(n_1583), .Y(n_1582) );
NOR2x1_ASAP7_75t_SL g1583 ( .A(n_1584), .B(n_1606), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1587 ( .A(n_1588), .B(n_1596), .Y(n_1587) );
OAI211xp5_ASAP7_75t_L g1588 ( .A1(n_1589), .A2(n_1590), .B(n_1591), .C(n_1592), .Y(n_1588) );
INVx2_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVxp33_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
NOR3xp33_ASAP7_75t_L g1610 ( .A(n_1611), .B(n_1616), .C(n_1619), .Y(n_1610) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
BUFx3_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
BUFx3_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
HB1xp67_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
endmodule