module fake_jpeg_8602_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_49),
.B(n_33),
.Y(n_90)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_20),
.B1(n_23),
.B2(n_21),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_59),
.B1(n_33),
.B2(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_16),
.B1(n_21),
.B2(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_26),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_28),
.B(n_26),
.Y(n_73)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_18),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_70),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_73),
.B(n_86),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_44),
.B(n_25),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_0),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_51),
.B1(n_60),
.B2(n_32),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_18),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_25),
.B(n_29),
.Y(n_115)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_79),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_88),
.B1(n_60),
.B2(n_47),
.Y(n_100)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_55),
.B1(n_48),
.B2(n_54),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_114),
.B1(n_81),
.B2(n_87),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_89),
.B1(n_91),
.B2(n_56),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_71),
.B(n_30),
.C(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_99),
.B(n_101),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_100),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_51),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_104),
.A2(n_112),
.B(n_115),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_24),
.B(n_29),
.C(n_60),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_70),
.B1(n_79),
.B2(n_83),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_32),
.B1(n_30),
.B2(n_17),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_43),
.C(n_24),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_1),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_88),
.B1(n_65),
.B2(n_67),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_122),
.A2(n_125),
.B1(n_127),
.B2(n_135),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_141),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_116),
.B1(n_97),
.B2(n_113),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_126),
.B1(n_131),
.B2(n_150),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_81),
.B1(n_66),
.B2(n_68),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_68),
.B1(n_66),
.B2(n_84),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_128),
.A2(n_140),
.B1(n_144),
.B2(n_4),
.Y(n_183)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_97),
.A3(n_104),
.B1(n_115),
.B2(n_99),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_2),
.C(n_3),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_85),
.B1(n_77),
.B2(n_78),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_136),
.B(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_151),
.Y(n_153)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_143),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_82),
.B1(n_80),
.B2(n_15),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_146),
.B1(n_4),
.B2(n_5),
.Y(n_185)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_15),
.B1(n_14),
.B2(n_3),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_147),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_102),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_117),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_154),
.B(n_155),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_138),
.A2(n_110),
.B1(n_119),
.B2(n_111),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_180),
.B1(n_152),
.B2(n_158),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_102),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_172),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_169),
.C(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_108),
.C(n_95),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_145),
.B(n_108),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_6),
.B(n_7),
.Y(n_199)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_134),
.B(n_136),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_176),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_104),
.Y(n_174)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_104),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_127),
.B(n_98),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_182),
.B(n_5),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_95),
.C(n_111),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_8),
.C(n_9),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_110),
.B1(n_106),
.B2(n_107),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_110),
.Y(n_181)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_3),
.B(n_4),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_172),
.A2(n_135),
.B1(n_129),
.B2(n_131),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_205),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_155),
.A2(n_135),
.B1(n_124),
.B2(n_144),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_184),
.A2(n_151),
.B1(n_150),
.B2(n_7),
.Y(n_194)
);

AO22x1_ASAP7_75t_SL g196 ( 
.A1(n_166),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_202),
.B1(n_207),
.B2(n_174),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_214),
.B(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_181),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_154),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_212),
.C(n_171),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_166),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_161),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_208),
.B1(n_211),
.B2(n_213),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_176),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_12),
.B1(n_13),
.B2(n_167),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_13),
.C(n_179),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_164),
.B1(n_162),
.B2(n_159),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_177),
.B(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_222),
.B(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_157),
.Y(n_220)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_153),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_221),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_169),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_175),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_237),
.C(n_212),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_191),
.A2(n_177),
.B1(n_171),
.B2(n_182),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_153),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_188),
.C(n_233),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_239),
.B(n_199),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_243),
.C(n_246),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_242),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_197),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_209),
.C(n_203),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_227),
.B(n_192),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_194),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_250),
.C(n_256),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_196),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_219),
.B(n_196),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_229),
.C(n_209),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_239),
.C(n_203),
.Y(n_272)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_217),
.B1(n_225),
.B2(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_253),
.A2(n_225),
.B1(n_230),
.B2(n_226),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_246),
.B1(n_256),
.B2(n_244),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_221),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_268),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_257),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_186),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_275),
.B(n_254),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_220),
.C(n_188),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_171),
.C(n_160),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_208),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_261),
.A2(n_196),
.B1(n_245),
.B2(n_251),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_163),
.Y(n_298)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_267),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_270),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_274),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_250),
.B1(n_255),
.B2(n_249),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_284),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_263),
.B1(n_271),
.B2(n_205),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_241),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_288),
.C(n_262),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_242),
.C(n_211),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_210),
.B(n_207),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_266),
.B(n_210),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_291),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_272),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_297),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_295),
.B1(n_278),
.B2(n_282),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_206),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_288),
.C(n_289),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_163),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_298),
.B(n_281),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_306),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_283),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_307),
.A2(n_308),
.B(n_299),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_283),
.B(n_285),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_309),
.B(n_312),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_303),
.A2(n_292),
.B(n_291),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_305),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_305),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_313),
.B(n_314),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_310),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_318),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_302),
.B(n_296),
.Y(n_321)
);


endmodule