module fake_jpeg_19498_n_298 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_265;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_123;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_39),
.Y(n_88)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_48),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_51),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_19),
.B(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_57),
.B(n_60),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_25),
.B1(n_34),
.B2(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_58),
.A2(n_63),
.B1(n_66),
.B2(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_70),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_25),
.B1(n_34),
.B2(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_65),
.B(n_67),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_25),
.B1(n_20),
.B2(n_38),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_36),
.Y(n_67)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_21),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_72),
.B(n_75),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_36),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_29),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_43),
.A2(n_52),
.B1(n_40),
.B2(n_20),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_82),
.B1(n_97),
.B2(n_4),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_23),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_80),
.B(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_23),
.B1(n_32),
.B2(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_45),
.B(n_37),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_37),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_41),
.B(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_42),
.B(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_13),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_91),
.Y(n_129)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_39),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_94),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_32),
.B1(n_30),
.B2(n_22),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_51),
.B(n_13),
.Y(n_98)
);

CKINVDCx12_ASAP7_75t_R g99 ( 
.A(n_49),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_50),
.A2(n_32),
.B1(n_30),
.B2(n_22),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_51),
.B(n_12),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_10),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_31),
.B(n_28),
.C(n_17),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_102),
.A2(n_116),
.B(n_106),
.Y(n_163)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_53),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_58),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_71),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_4),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_0),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_88),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_64),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_77),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_131),
.Y(n_143)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_91),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_67),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_134),
.B(n_151),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_136),
.B(n_137),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_118),
.B(n_116),
.C(n_131),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_139),
.A2(n_121),
.B(n_125),
.C(n_7),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_100),
.B1(n_66),
.B2(n_97),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_147),
.B1(n_148),
.B2(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_149),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_96),
.B1(n_73),
.B2(n_56),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_62),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_156),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_76),
.C(n_94),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_162),
.C(n_74),
.Y(n_174)
);

OAI22x1_ASAP7_75t_SL g154 ( 
.A1(n_110),
.A2(n_56),
.B1(n_73),
.B2(n_81),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_62),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_155),
.B(n_159),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_105),
.B(n_89),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_69),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_163),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_102),
.A2(n_84),
.B1(n_61),
.B2(n_54),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_161),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_95),
.C(n_93),
.Y(n_162)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_105),
.B(n_61),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_156),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_108),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_171),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_108),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_181),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_149),
.B(n_153),
.Y(n_180)
);

NOR4xp25_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_140),
.C(n_121),
.D(n_151),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_115),
.C(n_126),
.Y(n_181)
);

NOR4xp25_ASAP7_75t_SL g185 ( 
.A(n_154),
.B(n_114),
.C(n_6),
.D(n_7),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_6),
.C(n_7),
.Y(n_220)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_144),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_187),
.B(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_4),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_150),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_145),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_195),
.B(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_202),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_152),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_163),
.B(n_143),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_189),
.B(n_166),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_135),
.B1(n_147),
.B2(n_141),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_206),
.A2(n_207),
.B1(n_175),
.B2(n_181),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_148),
.B1(n_135),
.B2(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_209),
.B(n_215),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_162),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_210),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_166),
.A2(n_148),
.B(n_137),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_219),
.B(n_220),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_171),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_183),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_176),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_172),
.C(n_183),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_217),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_222),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_179),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_226),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_216),
.B(n_197),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_229),
.B(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_219),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_194),
.B(n_187),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_239),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_170),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_214),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_178),
.B(n_191),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_241),
.A2(n_254),
.B1(n_235),
.B2(n_228),
.Y(n_259)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_167),
.B(n_168),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_249),
.B1(n_253),
.B2(n_238),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_204),
.B1(n_169),
.B2(n_212),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_203),
.B1(n_177),
.B2(n_196),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_223),
.B(n_236),
.C(n_224),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_6),
.B(n_10),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_209),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_206),
.C(n_208),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_227),
.C(n_231),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g252 ( 
.A1(n_236),
.A2(n_218),
.A3(n_198),
.B1(n_200),
.B2(n_186),
.C1(n_177),
.C2(n_178),
.Y(n_252)
);

OAI322xp33_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_235),
.A3(n_228),
.B1(n_198),
.B2(n_238),
.C1(n_237),
.C2(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_200),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_264),
.B1(n_241),
.B2(n_254),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_230),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_261),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_232),
.B1(n_225),
.B2(n_226),
.Y(n_257)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

OAI21x1_ASAP7_75t_SL g258 ( 
.A1(n_251),
.A2(n_227),
.B(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_266),
.B(n_240),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_263),
.Y(n_269)
);

XOR2x2_ASAP7_75t_SL g262 ( 
.A(n_251),
.B(n_230),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_247),
.B(n_246),
.Y(n_272)
);

NAND4xp25_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_237),
.C(n_203),
.D(n_167),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_267),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_264),
.A2(n_243),
.B1(n_253),
.B2(n_240),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_275),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_168),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_267),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_263),
.C(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_281),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_259),
.C(n_261),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_244),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_10),
.B(n_11),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_283),
.A2(n_284),
.B1(n_270),
.B2(n_276),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_257),
.A3(n_262),
.B1(n_258),
.B2(n_256),
.C1(n_265),
.C2(n_188),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_268),
.B1(n_274),
.B2(n_279),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_288),
.B1(n_289),
.B2(n_117),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_11),
.B(n_12),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_SL g288 ( 
.A1(n_284),
.A2(n_270),
.B(n_271),
.C(n_167),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_188),
.C(n_161),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_126),
.C(n_123),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_293),
.A2(n_117),
.B(n_103),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_295),
.B(n_12),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_123),
.C(n_115),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_297),
.Y(n_298)
);


endmodule