module fake_jpeg_30667_n_41 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

INVx4_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_1),
.Y(n_18)
);

OAI21xp33_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_21),
.B(n_22),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_4),
.Y(n_23)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_25),
.B1(n_26),
.B2(n_7),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_11),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_16),
.B1(n_8),
.B2(n_7),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22x1_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_14),
.B1(n_16),
.B2(n_11),
.Y(n_28)
);

NAND5xp2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.C(n_12),
.D(n_17),
.E(n_31),
.Y(n_36)
);

AOI321xp33_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_27),
.A3(n_29),
.B1(n_18),
.B2(n_19),
.C(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_22),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_36),
.C(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_36),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_40),
.B(n_12),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_32),
.B(n_17),
.Y(n_40)
);


endmodule