module real_aes_10044_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_265;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g1073 ( .A(n_0), .Y(n_1073) );
AO22x2_ASAP7_75t_L g1008 ( .A1(n_1), .A2(n_1009), .B1(n_1055), .B2(n_1056), .Y(n_1008) );
INVxp67_ASAP7_75t_L g1055 ( .A(n_1), .Y(n_1055) );
AOI22xp5_ASAP7_75t_L g1190 ( .A1(n_1), .A2(n_2), .B1(n_1162), .B2(n_1191), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1449 ( .A1(n_3), .A2(n_217), .B1(n_886), .B2(n_1002), .Y(n_1449) );
INVx1_ASAP7_75t_L g1455 ( .A(n_3), .Y(n_1455) );
CKINVDCx5p33_ASAP7_75t_R g1091 ( .A(n_4), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_5), .B(n_189), .Y(n_363) );
AND2x2_ASAP7_75t_L g375 ( .A(n_5), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g403 ( .A(n_5), .Y(n_403) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_5), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_6), .A2(n_148), .B1(n_325), .B2(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g434 ( .A(n_6), .Y(n_434) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_7), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_7), .A2(n_236), .B1(n_733), .B2(n_735), .C(n_736), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g1195 ( .A1(n_8), .A2(n_216), .B1(n_1174), .B2(n_1180), .Y(n_1195) );
INVx1_ASAP7_75t_L g785 ( .A(n_9), .Y(n_785) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_9), .A2(n_131), .B1(n_826), .B2(n_829), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_10), .Y(n_1090) );
INVx1_ASAP7_75t_L g1434 ( .A(n_11), .Y(n_1434) );
OAI22xp5_ASAP7_75t_L g1453 ( .A1(n_11), .A2(n_62), .B1(n_861), .B2(n_912), .Y(n_1453) );
CKINVDCx14_ASAP7_75t_R g1199 ( .A(n_12), .Y(n_1199) );
INVxp33_ASAP7_75t_SL g683 ( .A(n_13), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_13), .A2(n_66), .B1(n_658), .B2(n_720), .C(n_722), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_14), .A2(n_97), .B1(n_541), .B2(n_658), .Y(n_1387) );
INVxp67_ASAP7_75t_SL g1411 ( .A(n_14), .Y(n_1411) );
INVx1_ASAP7_75t_L g1390 ( .A(n_15), .Y(n_1390) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_16), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_17), .Y(n_671) );
INVxp67_ASAP7_75t_SL g761 ( .A(n_18), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_18), .A2(n_225), .B1(n_659), .B2(n_812), .Y(n_820) );
OAI221xp5_ASAP7_75t_L g582 ( .A1(n_19), .A2(n_81), .B1(n_583), .B2(n_590), .C(n_593), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_19), .A2(n_81), .B1(n_643), .B2(n_646), .Y(n_642) );
INVx1_ASAP7_75t_L g915 ( .A(n_20), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_20), .A2(n_187), .B1(n_541), .B2(n_886), .Y(n_941) );
OR2x2_ASAP7_75t_L g269 ( .A(n_21), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g308 ( .A(n_21), .Y(n_308) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_22), .A2(n_67), .B1(n_797), .B2(n_802), .Y(n_801) );
INVxp33_ASAP7_75t_L g834 ( .A(n_22), .Y(n_834) );
INVx1_ASAP7_75t_L g477 ( .A(n_23), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_23), .A2(n_165), .B1(n_544), .B2(n_547), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_24), .Y(n_297) );
INVx1_ASAP7_75t_L g741 ( .A(n_25), .Y(n_741) );
INVx1_ASAP7_75t_L g271 ( .A(n_26), .Y(n_271) );
BUFx2_ASAP7_75t_L g323 ( .A(n_26), .Y(n_323) );
BUFx2_ASAP7_75t_L g345 ( .A(n_26), .Y(n_345) );
OR2x2_ASAP7_75t_L g589 ( .A(n_26), .B(n_363), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g871 ( .A1(n_27), .A2(n_184), .B1(n_872), .B2(n_873), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_27), .A2(n_184), .B1(n_553), .B2(n_880), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g1376 ( .A1(n_28), .A2(n_138), .B1(n_639), .B2(n_1002), .Y(n_1376) );
INVxp33_ASAP7_75t_SL g1401 ( .A(n_28), .Y(n_1401) );
INVx1_ASAP7_75t_L g461 ( .A(n_29), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_29), .A2(n_137), .B1(n_342), .B2(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g1388 ( .A(n_30), .Y(n_1388) );
INVx1_ASAP7_75t_L g777 ( .A(n_31), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_31), .A2(n_55), .B1(n_331), .B2(n_818), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_32), .A2(n_212), .B1(n_829), .B2(n_1018), .C(n_1019), .Y(n_1017) );
INVx1_ASAP7_75t_L g1026 ( .A(n_32), .Y(n_1026) );
OAI221xp5_ASAP7_75t_L g687 ( .A1(n_33), .A2(n_50), .B1(n_583), .B2(n_593), .C(n_688), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_33), .A2(n_50), .B1(n_643), .B2(n_730), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_34), .A2(n_89), .B1(n_815), .B2(n_903), .Y(n_1066) );
AOI221xp5_ASAP7_75t_L g1085 ( .A1(n_34), .A2(n_89), .B1(n_471), .B2(n_472), .C(n_574), .Y(n_1085) );
OAI22xp33_ASAP7_75t_L g862 ( .A1(n_35), .A2(n_53), .B1(n_771), .B2(n_775), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_35), .A2(n_163), .B1(n_738), .B2(n_884), .Y(n_883) );
CKINVDCx5p33_ASAP7_75t_R g981 ( .A(n_36), .Y(n_981) );
CKINVDCx5p33_ASAP7_75t_R g1074 ( .A(n_37), .Y(n_1074) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_38), .Y(n_951) );
AOI22xp33_ASAP7_75t_SL g1070 ( .A1(n_39), .A2(n_43), .B1(n_292), .B2(n_813), .Y(n_1070) );
INVx1_ASAP7_75t_L g1081 ( .A(n_39), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_40), .A2(n_246), .B1(n_872), .B2(n_926), .Y(n_925) );
AOI22xp33_ASAP7_75t_SL g935 ( .A1(n_40), .A2(n_246), .B1(n_650), .B2(n_936), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_41), .A2(n_68), .B1(n_797), .B2(n_799), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_41), .A2(n_68), .B1(n_812), .B2(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g1438 ( .A(n_42), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g1443 ( .A1(n_42), .A2(n_227), .B1(n_928), .B2(n_930), .Y(n_1443) );
INVx1_ASAP7_75t_L g1080 ( .A(n_43), .Y(n_1080) );
INVx1_ASAP7_75t_L g897 ( .A(n_44), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_44), .A2(n_141), .B1(n_928), .B2(n_930), .Y(n_927) );
INVx1_ASAP7_75t_L g1391 ( .A(n_45), .Y(n_1391) );
AOI221xp5_ASAP7_75t_L g1126 ( .A1(n_46), .A2(n_61), .B1(n_471), .B2(n_472), .C(n_780), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_46), .A2(n_61), .B1(n_331), .B2(n_1133), .Y(n_1132) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_47), .Y(n_619) );
INVx1_ASAP7_75t_L g706 ( .A(n_48), .Y(n_706) );
INVx1_ASAP7_75t_L g281 ( .A(n_49), .Y(n_281) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_49), .A2(n_51), .B1(n_394), .B2(n_396), .C(n_399), .Y(n_393) );
INVx1_ASAP7_75t_L g272 ( .A(n_51), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_52), .A2(n_78), .B1(n_794), .B2(n_805), .Y(n_804) );
INVxp67_ASAP7_75t_SL g823 ( .A(n_52), .Y(n_823) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_53), .A2(n_208), .B1(n_854), .B2(n_856), .Y(n_853) );
INVx1_ASAP7_75t_L g902 ( .A(n_54), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_54), .A2(n_104), .B1(n_778), .B2(n_932), .Y(n_931) );
INVxp33_ASAP7_75t_L g769 ( .A(n_55), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g1196 ( .A1(n_56), .A2(n_80), .B1(n_1162), .B2(n_1191), .Y(n_1196) );
AO221x1_ASAP7_75t_L g1088 ( .A1(n_57), .A2(n_75), .B1(n_494), .B2(n_495), .C(n_806), .Y(n_1088) );
INVx1_ASAP7_75t_L g1100 ( .A(n_57), .Y(n_1100) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_58), .A2(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g504 ( .A(n_58), .Y(n_504) );
INVx1_ASAP7_75t_L g944 ( .A(n_59), .Y(n_944) );
AOI22xp5_ASAP7_75t_SL g1183 ( .A1(n_59), .A2(n_73), .B1(n_1162), .B2(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1024 ( .A(n_60), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_60), .A2(n_194), .B1(n_292), .B2(n_1002), .Y(n_1054) );
INVx1_ASAP7_75t_L g1435 ( .A(n_62), .Y(n_1435) );
CKINVDCx16_ASAP7_75t_R g1222 ( .A(n_63), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_64), .A2(n_205), .B1(n_797), .B2(n_1037), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_64), .A2(n_205), .B1(n_812), .B2(n_1002), .Y(n_1044) );
INVx1_ASAP7_75t_L g964 ( .A(n_65), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_65), .A2(n_82), .B1(n_658), .B2(n_1002), .Y(n_1001) );
INVxp33_ASAP7_75t_L g685 ( .A(n_66), .Y(n_685) );
INVxp67_ASAP7_75t_SL g835 ( .A(n_67), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_69), .A2(n_107), .B1(n_851), .B2(n_852), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_69), .A2(n_107), .B1(n_486), .B2(n_873), .Y(n_874) );
XNOR2x2_ASAP7_75t_L g892 ( .A(n_70), .B(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g848 ( .A(n_71), .Y(n_848) );
OAI222xp33_ASAP7_75t_L g859 ( .A1(n_71), .A2(n_163), .B1(n_177), .B2(n_492), .C1(n_860), .C2(n_861), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_72), .A2(n_155), .B1(n_341), .B2(n_343), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_72), .A2(n_155), .B1(n_442), .B2(n_447), .Y(n_441) );
INVxp33_ASAP7_75t_L g691 ( .A(n_74), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_74), .A2(n_112), .B1(n_541), .B2(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g1102 ( .A(n_75), .Y(n_1102) );
AOI221xp5_ASAP7_75t_L g1114 ( .A1(n_76), .A2(n_86), .B1(n_399), .B2(n_1115), .C(n_1116), .Y(n_1114) );
INVx1_ASAP7_75t_L g1138 ( .A(n_76), .Y(n_1138) );
INVx1_ASAP7_75t_L g270 ( .A(n_77), .Y(n_270) );
INVx1_ASAP7_75t_L g321 ( .A(n_77), .Y(n_321) );
INVxp33_ASAP7_75t_L g831 ( .A(n_78), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g1093 ( .A(n_79), .Y(n_1093) );
AOI222xp33_ASAP7_75t_L g1367 ( .A1(n_80), .A2(n_1368), .B1(n_1417), .B2(n_1421), .C1(n_1461), .C2(n_1465), .Y(n_1367) );
INVx1_ASAP7_75t_L g1416 ( .A(n_80), .Y(n_1416) );
INVx1_ASAP7_75t_L g971 ( .A(n_82), .Y(n_971) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_83), .A2(n_221), .B1(n_486), .B2(n_487), .C(n_490), .Y(n_485) );
INVx1_ASAP7_75t_L g509 ( .A(n_83), .Y(n_509) );
AOI22x1_ASAP7_75t_L g1059 ( .A1(n_84), .A2(n_1060), .B1(n_1061), .B2(n_1103), .Y(n_1059) );
INVxp67_ASAP7_75t_SL g1103 ( .A(n_84), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1441 ( .A1(n_85), .A2(n_130), .B1(n_876), .B2(n_924), .Y(n_1441) );
AOI22xp33_ASAP7_75t_L g1446 ( .A1(n_85), .A2(n_130), .B1(n_939), .B2(n_1384), .Y(n_1446) );
INVx1_ASAP7_75t_L g1140 ( .A(n_86), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_87), .A2(n_220), .B1(n_1174), .B2(n_1235), .Y(n_1234) );
CKINVDCx20_ASAP7_75t_R g1244 ( .A(n_88), .Y(n_1244) );
INVx1_ASAP7_75t_L g967 ( .A(n_90), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g998 ( .A1(n_90), .A2(n_211), .B1(n_630), .B2(n_720), .C(n_999), .Y(n_998) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_91), .Y(n_614) );
INVx1_ASAP7_75t_L g1122 ( .A(n_92), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_92), .A2(n_218), .B1(n_630), .B2(n_993), .Y(n_1135) );
INVx1_ASAP7_75t_L g572 ( .A(n_93), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_93), .A2(n_207), .B1(n_633), .B2(n_634), .C(n_636), .Y(n_632) );
INVx1_ASAP7_75t_L g712 ( .A(n_94), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_95), .A2(n_203), .B1(n_1112), .B2(n_1128), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_95), .A2(n_203), .B1(n_630), .B2(n_641), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_96), .A2(n_242), .B1(n_794), .B2(n_795), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_96), .A2(n_242), .B1(n_635), .B2(n_815), .Y(n_814) );
INVxp33_ASAP7_75t_L g1406 ( .A(n_97), .Y(n_1406) );
INVx1_ASAP7_75t_L g1377 ( .A(n_98), .Y(n_1377) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_99), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_100), .A2(n_174), .B1(n_1046), .B2(n_1068), .Y(n_1067) );
OAI221xp5_ASAP7_75t_L g1087 ( .A1(n_100), .A2(n_371), .B1(n_1088), .B2(n_1089), .C(n_1092), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_101), .A2(n_197), .B1(n_343), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_SL g1083 ( .A1(n_101), .A2(n_197), .B1(n_489), .B2(n_1084), .Y(n_1083) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_102), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g1442 ( .A1(n_103), .A2(n_224), .B1(n_872), .B2(n_926), .Y(n_1442) );
AOI22xp33_ASAP7_75t_L g1447 ( .A1(n_103), .A2(n_224), .B1(n_639), .B2(n_1002), .Y(n_1447) );
INVx1_ASAP7_75t_L g896 ( .A(n_104), .Y(n_896) );
INVx1_ASAP7_75t_L g1152 ( .A(n_105), .Y(n_1152) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_106), .Y(n_484) );
AOI21xp33_ASAP7_75t_L g470 ( .A1(n_108), .A2(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g539 ( .A(n_108), .Y(n_539) );
XOR2xp5_ASAP7_75t_L g563 ( .A(n_109), .B(n_564), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g1429 ( .A(n_110), .Y(n_1429) );
INVx1_ASAP7_75t_L g1020 ( .A(n_111), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_111), .A2(n_136), .B1(n_794), .B2(n_869), .Y(n_1042) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_112), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g980 ( .A(n_113), .Y(n_980) );
XNOR2xp5_ASAP7_75t_L g255 ( .A(n_114), .B(n_256), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_115), .A2(n_206), .B1(n_1112), .B2(n_1113), .Y(n_1111) );
INVx1_ASAP7_75t_L g1141 ( .A(n_115), .Y(n_1141) );
INVx1_ASAP7_75t_L g1125 ( .A(n_116), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_116), .A2(n_237), .B1(n_283), .B2(n_350), .Y(n_1134) );
INVx1_ASAP7_75t_L g601 ( .A(n_117), .Y(n_601) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_117), .A2(n_162), .B1(n_650), .B2(n_652), .C(n_654), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g1173 ( .A1(n_118), .A2(n_204), .B1(n_1174), .B2(n_1180), .Y(n_1173) );
INVx1_ASAP7_75t_L g610 ( .A(n_119), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_119), .A2(n_152), .B1(n_658), .B2(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g910 ( .A(n_120), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_120), .A2(n_190), .B1(n_658), .B2(n_845), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g1448 ( .A1(n_121), .A2(n_228), .B1(n_658), .B2(n_1384), .Y(n_1448) );
INVx1_ASAP7_75t_L g1458 ( .A(n_121), .Y(n_1458) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_122), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g975 ( .A(n_123), .Y(n_975) );
INVx1_ASAP7_75t_L g579 ( .A(n_124), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_124), .A2(n_245), .B1(n_639), .B2(n_640), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_125), .A2(n_126), .B1(n_1184), .B2(n_1237), .Y(n_1236) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_127), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g1378 ( .A1(n_128), .A2(n_180), .B1(n_1379), .B2(n_1380), .Y(n_1378) );
OAI221xp5_ASAP7_75t_L g1402 ( .A1(n_128), .A2(n_180), .B1(n_583), .B2(n_590), .C(n_1403), .Y(n_1402) );
XNOR2xp5_ASAP7_75t_L g1422 ( .A(n_129), .B(n_1423), .Y(n_1422) );
INVxp67_ASAP7_75t_SL g781 ( .A(n_131), .Y(n_781) );
CKINVDCx14_ASAP7_75t_R g1201 ( .A(n_132), .Y(n_1201) );
INVx1_ASAP7_75t_L g1033 ( .A(n_133), .Y(n_1033) );
AOI22xp33_ASAP7_75t_SL g1052 ( .A1(n_133), .A2(n_139), .B1(n_1046), .B2(n_1053), .Y(n_1052) );
AOI22xp5_ASAP7_75t_L g1189 ( .A1(n_134), .A2(n_156), .B1(n_1174), .B2(n_1180), .Y(n_1189) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_135), .A2(n_200), .B1(n_409), .B2(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1144 ( .A(n_135), .Y(n_1144) );
INVx1_ASAP7_75t_L g1012 ( .A(n_136), .Y(n_1012) );
INVx1_ASAP7_75t_L g462 ( .A(n_137), .Y(n_462) );
INVxp33_ASAP7_75t_L g1396 ( .A(n_138), .Y(n_1396) );
INVx1_ASAP7_75t_L g1028 ( .A(n_139), .Y(n_1028) );
INVx1_ASAP7_75t_L g949 ( .A(n_140), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_140), .A2(n_232), .B1(n_651), .B2(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g900 ( .A(n_141), .Y(n_900) );
INVx1_ASAP7_75t_L g1145 ( .A(n_142), .Y(n_1145) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_143), .Y(n_899) );
INVx1_ASAP7_75t_L g864 ( .A(n_144), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_144), .A2(n_147), .B1(n_541), .B2(n_886), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_145), .A2(n_175), .B1(n_396), .B2(n_869), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_145), .A2(n_175), .B1(n_815), .B2(n_1046), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_146), .A2(n_172), .B1(n_876), .B2(n_924), .Y(n_923) );
AOI22xp33_ASAP7_75t_SL g938 ( .A1(n_146), .A2(n_172), .B1(n_845), .B2(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g865 ( .A(n_147), .Y(n_865) );
INVx1_ASAP7_75t_L g436 ( .A(n_148), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_149), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_150), .A2(n_196), .B1(n_331), .B2(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g420 ( .A(n_150), .Y(n_420) );
INVx1_ASAP7_75t_L g1392 ( .A(n_151), .Y(n_1392) );
INVx1_ASAP7_75t_L g598 ( .A(n_152), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g977 ( .A(n_153), .Y(n_977) );
AOI22x1_ASAP7_75t_SL g839 ( .A1(n_154), .A2(n_840), .B1(n_887), .B2(n_888), .Y(n_839) );
INVx1_ASAP7_75t_L g887 ( .A(n_154), .Y(n_887) );
AO221x2_ASAP7_75t_L g1197 ( .A1(n_154), .A2(n_231), .B1(n_1162), .B2(n_1191), .C(n_1198), .Y(n_1197) );
CKINVDCx16_ASAP7_75t_R g1223 ( .A(n_157), .Y(n_1223) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_158), .Y(n_290) );
INVx1_ASAP7_75t_L g710 ( .A(n_159), .Y(n_710) );
INVx1_ASAP7_75t_L g844 ( .A(n_160), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_160), .A2(n_208), .B1(n_869), .B2(n_876), .Y(n_875) );
HB1xp67_ASAP7_75t_L g1154 ( .A(n_161), .Y(n_1154) );
AND3x2_ASAP7_75t_L g1165 ( .A(n_161), .B(n_1152), .C(n_1166), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_161), .B(n_1152), .Y(n_1179) );
INVx1_ASAP7_75t_L g604 ( .A(n_162), .Y(n_604) );
AOI22xp5_ASAP7_75t_SL g1240 ( .A1(n_164), .A2(n_176), .B1(n_1162), .B2(n_1184), .Y(n_1240) );
INVx1_ASAP7_75t_L g466 ( .A(n_165), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_166), .Y(n_491) );
AOI221xp5_ASAP7_75t_L g1375 ( .A1(n_167), .A2(n_214), .B1(n_337), .B2(n_903), .C(n_996), .Y(n_1375) );
INVxp33_ASAP7_75t_L g1398 ( .A(n_167), .Y(n_1398) );
INVx2_ASAP7_75t_L g367 ( .A(n_168), .Y(n_367) );
AOI22xp5_ASAP7_75t_SL g1239 ( .A1(n_169), .A2(n_226), .B1(n_1174), .B2(n_1180), .Y(n_1239) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_170), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_171), .Y(n_481) );
XOR2xp5_ASAP7_75t_L g676 ( .A(n_173), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g1086 ( .A(n_174), .Y(n_1086) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_177), .Y(n_847) );
INVx1_ASAP7_75t_L g904 ( .A(n_178), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_178), .A2(n_199), .B1(n_912), .B2(n_913), .Y(n_911) );
INVx1_ASAP7_75t_L g1166 ( .A(n_179), .Y(n_1166) );
INVx1_ASAP7_75t_L g353 ( .A(n_181), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g751 ( .A(n_182), .Y(n_751) );
AOI221xp5_ASAP7_75t_L g1383 ( .A1(n_183), .A2(n_241), .B1(n_630), .B2(n_1384), .C(n_1386), .Y(n_1383) );
INVxp67_ASAP7_75t_SL g1409 ( .A(n_183), .Y(n_1409) );
AO221x2_ASAP7_75t_L g1241 ( .A1(n_185), .A2(n_248), .B1(n_1237), .B2(n_1242), .C(n_1243), .Y(n_1241) );
AOI22xp33_ASAP7_75t_SL g868 ( .A1(n_186), .A2(n_223), .B1(n_471), .B2(n_869), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_186), .A2(n_223), .B1(n_658), .B2(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g916 ( .A(n_187), .Y(n_916) );
OAI221xp5_ASAP7_75t_L g956 ( .A1(n_188), .A2(n_192), .B1(n_583), .B2(n_590), .C(n_957), .Y(n_956) );
OAI221xp5_ASAP7_75t_L g986 ( .A1(n_188), .A2(n_192), .B1(n_646), .B2(n_987), .C(n_989), .Y(n_986) );
INVx2_ASAP7_75t_L g376 ( .A(n_189), .Y(n_376) );
INVx1_ASAP7_75t_L g432 ( .A(n_189), .Y(n_432) );
INVx1_ASAP7_75t_L g918 ( .A(n_190), .Y(n_918) );
CKINVDCx14_ASAP7_75t_R g1246 ( .A(n_191), .Y(n_1246) );
AO22x2_ASAP7_75t_L g452 ( .A1(n_193), .A2(n_453), .B1(n_557), .B2(n_558), .Y(n_452) );
INVxp67_ASAP7_75t_SL g557 ( .A(n_193), .Y(n_557) );
INVx1_ASAP7_75t_L g1023 ( .A(n_194), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_195), .B(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g426 ( .A(n_196), .Y(n_426) );
INVx1_ASAP7_75t_L g715 ( .A(n_198), .Y(n_715) );
INVx1_ASAP7_75t_L g907 ( .A(n_199), .Y(n_907) );
INVx1_ASAP7_75t_L g1143 ( .A(n_200), .Y(n_1143) );
CKINVDCx16_ASAP7_75t_R g1219 ( .A(n_201), .Y(n_1219) );
INVx1_ASAP7_75t_L g1437 ( .A(n_202), .Y(n_1437) );
AOI22xp33_ASAP7_75t_L g1444 ( .A1(n_202), .A2(n_209), .B1(n_876), .B2(n_924), .Y(n_1444) );
INVx1_ASAP7_75t_L g1137 ( .A(n_206), .Y(n_1137) );
INVx1_ASAP7_75t_L g576 ( .A(n_207), .Y(n_576) );
INVx1_ASAP7_75t_L g1432 ( .A(n_209), .Y(n_1432) );
INVx1_ASAP7_75t_L g773 ( .A(n_210), .Y(n_773) );
INVx1_ASAP7_75t_L g965 ( .A(n_211), .Y(n_965) );
INVx1_ASAP7_75t_L g1027 ( .A(n_212), .Y(n_1027) );
INVxp33_ASAP7_75t_SL g686 ( .A(n_213), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_213), .A2(n_219), .B1(n_726), .B2(n_728), .Y(n_725) );
INVxp33_ASAP7_75t_L g1400 ( .A(n_214), .Y(n_1400) );
INVx1_ASAP7_75t_L g1164 ( .A(n_215), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_215), .B(n_1177), .Y(n_1182) );
INVx1_ASAP7_75t_L g1456 ( .A(n_217), .Y(n_1456) );
INVx1_ASAP7_75t_L g1123 ( .A(n_218), .Y(n_1123) );
INVxp33_ASAP7_75t_SL g681 ( .A(n_219), .Y(n_681) );
INVx1_ASAP7_75t_L g517 ( .A(n_221), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_222), .Y(n_261) );
INVx1_ASAP7_75t_L g758 ( .A(n_225), .Y(n_758) );
INVx1_ASAP7_75t_L g1430 ( .A(n_227), .Y(n_1430) );
INVx1_ASAP7_75t_L g1452 ( .A(n_228), .Y(n_1452) );
INVx1_ASAP7_75t_L g953 ( .A(n_229), .Y(n_953) );
AOI21xp33_ASAP7_75t_L g994 ( .A1(n_229), .A2(n_995), .B(n_996), .Y(n_994) );
INVx2_ASAP7_75t_L g368 ( .A(n_230), .Y(n_368) );
INVx1_ASAP7_75t_L g954 ( .A(n_232), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_233), .A2(n_234), .B1(n_332), .B2(n_337), .Y(n_336) );
OAI211xp5_ASAP7_75t_SL g370 ( .A1(n_233), .A2(n_371), .B(n_381), .C(n_404), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_234), .A2(n_412), .B1(n_414), .B2(n_433), .C(n_439), .Y(n_411) );
INVx1_ASAP7_75t_L g1016 ( .A(n_235), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_235), .A2(n_239), .B1(n_797), .B2(n_1041), .Y(n_1040) );
INVxp33_ASAP7_75t_SL g695 ( .A(n_236), .Y(n_695) );
INVx1_ASAP7_75t_L g1117 ( .A(n_237), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g983 ( .A(n_238), .Y(n_983) );
INVx1_ASAP7_75t_L g1013 ( .A(n_239), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g1216 ( .A(n_240), .Y(n_1216) );
INVxp33_ASAP7_75t_SL g1407 ( .A(n_241), .Y(n_1407) );
INVx1_ASAP7_75t_L g267 ( .A(n_243), .Y(n_267) );
BUFx3_ASAP7_75t_L g287 ( .A(n_243), .Y(n_287) );
BUFx3_ASAP7_75t_L g266 ( .A(n_244), .Y(n_266) );
INVx1_ASAP7_75t_L g279 ( .A(n_244), .Y(n_279) );
INVx1_ASAP7_75t_L g568 ( .A(n_245), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_247), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_1148), .B(n_1158), .Y(n_249) );
XNOR2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_745), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AOI22x1_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_561), .B1(n_743), .B2(n_744), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g743 ( .A(n_254), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_452), .B1(n_559), .B2(n_560), .Y(n_254) );
INVx1_ASAP7_75t_L g559 ( .A(n_255), .Y(n_559) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND3xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_352), .C(n_369), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_295), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_280), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B1(n_272), .B2(n_273), .Y(n_260) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_261), .A2(n_290), .B1(n_382), .B2(n_387), .C(n_393), .Y(n_381) );
AOI222xp33_ASAP7_75t_L g1099 ( .A1(n_262), .A2(n_282), .B1(n_355), .B2(n_1090), .C1(n_1093), .C2(n_1100), .Y(n_1099) );
AOI22xp5_ASAP7_75t_L g1136 ( .A1(n_262), .A2(n_273), .B1(n_1137), .B2(n_1138), .Y(n_1136) );
CKINVDCx6p67_ASAP7_75t_R g262 ( .A(n_263), .Y(n_262) );
OR2x6_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
INVx2_ASAP7_75t_L g641 ( .A(n_264), .Y(n_641) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g329 ( .A(n_265), .Y(n_329) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_265), .Y(n_519) );
INVx1_ASAP7_75t_L g542 ( .A(n_265), .Y(n_542) );
BUFx6f_ASAP7_75t_L g993 ( .A(n_265), .Y(n_993) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g288 ( .A(n_266), .Y(n_288) );
AND2x2_ASAP7_75t_L g335 ( .A(n_266), .B(n_287), .Y(n_335) );
INVx1_ASAP7_75t_L g277 ( .A(n_267), .Y(n_277) );
OR2x6_ASAP7_75t_L g274 ( .A(n_268), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g289 ( .A(n_268), .Y(n_289) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx2_ASAP7_75t_L g631 ( .A(n_269), .Y(n_631) );
OR2x2_ASAP7_75t_L g668 ( .A(n_269), .B(n_538), .Y(n_668) );
OR2x2_ASAP7_75t_L g670 ( .A(n_269), .B(n_329), .Y(n_670) );
INVx1_ASAP7_75t_L g306 ( .A(n_270), .Y(n_306) );
INVx1_ASAP7_75t_L g309 ( .A(n_271), .Y(n_309) );
AND2x4_ASAP7_75t_L g571 ( .A(n_271), .B(n_375), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g1101 ( .A1(n_273), .A2(n_291), .B1(n_1091), .B2(n_1102), .Y(n_1101) );
CKINVDCx6p67_ASAP7_75t_R g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g551 ( .A(n_276), .Y(n_551) );
BUFx4f_ASAP7_75t_L g991 ( .A(n_276), .Y(n_991) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OR2x2_ASAP7_75t_L g538 ( .A(n_277), .B(n_278), .Y(n_538) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g294 ( .A(n_279), .B(n_287), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_290), .B2(n_291), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g1139 ( .A1(n_282), .A2(n_291), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_289), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g658 ( .A(n_284), .Y(n_658) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
INVx6_ASAP7_75t_L g339 ( .A(n_285), .Y(n_339) );
AND2x2_ASAP7_75t_L g356 ( .A(n_285), .B(n_305), .Y(n_356) );
AND2x4_ASAP7_75t_L g514 ( .A(n_285), .B(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g315 ( .A(n_286), .Y(n_315) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g302 ( .A(n_288), .Y(n_302) );
AND2x2_ASAP7_75t_L g291 ( .A(n_289), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g1065 ( .A(n_293), .Y(n_1065) );
INVx2_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_L g325 ( .A(n_294), .Y(n_325) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_294), .Y(n_342) );
AND2x6_ASAP7_75t_L g510 ( .A(n_294), .B(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_294), .Y(n_546) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_294), .Y(n_630) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_294), .Y(n_651) );
BUFx2_ASAP7_75t_L g812 ( .A(n_294), .Y(n_812) );
NAND3xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_316), .C(n_347), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B1(n_310), .B2(n_311), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_297), .A2(n_310), .B1(n_405), .B2(n_408), .Y(n_404) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g1072 ( .A(n_299), .Y(n_1072) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g645 ( .A(n_301), .Y(n_645) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g526 ( .A(n_302), .Y(n_526) );
INVx2_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
OR2x6_ASAP7_75t_L g312 ( .A(n_304), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g351 ( .A(n_304), .Y(n_351) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_305), .B(n_309), .Y(n_304) );
AND2x4_ASAP7_75t_L g644 ( .A(n_305), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g647 ( .A(n_305), .B(n_314), .Y(n_647) );
INVx1_ASAP7_75t_L g664 ( .A(n_305), .Y(n_664) );
AND2x4_ASAP7_75t_L g988 ( .A(n_305), .B(n_645), .Y(n_988) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_305), .B(n_314), .Y(n_1381) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x4_ASAP7_75t_L g346 ( .A(n_307), .B(n_321), .Y(n_346) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g320 ( .A(n_308), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g507 ( .A(n_308), .Y(n_507) );
INVx1_ASAP7_75t_L g512 ( .A(n_308), .Y(n_512) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_308), .Y(n_516) );
OR2x6_ASAP7_75t_L g623 ( .A(n_309), .B(n_401), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g1071 ( .A1(n_311), .A2(n_1072), .B1(n_1073), .B2(n_1074), .C(n_1075), .Y(n_1071) );
AOI221xp5_ASAP7_75t_L g1142 ( .A1(n_311), .A2(n_1072), .B1(n_1075), .B2(n_1143), .C(n_1144), .Y(n_1142) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g730 ( .A(n_313), .B(n_664), .Y(n_730) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x6_ASAP7_75t_L g527 ( .A(n_315), .B(n_512), .Y(n_527) );
AOI33xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_324), .A3(n_330), .B1(n_336), .B2(n_340), .B3(n_344), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_318), .A2(n_534), .B1(n_548), .B2(n_554), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g878 ( .A(n_318), .Y(n_878) );
OR2x6_ASAP7_75t_L g318 ( .A(n_319), .B(n_322), .Y(n_318) );
OR2x2_ASAP7_75t_L g810 ( .A(n_319), .B(n_322), .Y(n_810) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_SL g656 ( .A(n_320), .Y(n_656) );
INVx1_ASAP7_75t_L g736 ( .A(n_320), .Y(n_736) );
BUFx3_ASAP7_75t_L g1000 ( .A(n_320), .Y(n_1000) );
INVx1_ASAP7_75t_L g1050 ( .A(n_320), .Y(n_1050) );
INVx1_ASAP7_75t_L g500 ( .A(n_321), .Y(n_500) );
INVx2_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
BUFx2_ASAP7_75t_L g451 ( .A(n_322), .Y(n_451) );
AND2x4_ASAP7_75t_L g792 ( .A(n_322), .B(n_429), .Y(n_792) );
AND2x4_ASAP7_75t_L g922 ( .A(n_322), .B(n_429), .Y(n_922) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_322), .B(n_1050), .Y(n_1049) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx2_ASAP7_75t_L g501 ( .A(n_323), .Y(n_501) );
OR2x6_ASAP7_75t_L g596 ( .A(n_323), .B(n_472), .Y(n_596) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g343 ( .A(n_327), .Y(n_343) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g728 ( .A(n_328), .Y(n_728) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g845 ( .A(n_333), .Y(n_845) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_334), .Y(n_350) );
INVx1_ASAP7_75t_L g522 ( .A(n_334), .Y(n_522) );
AND2x4_ASAP7_75t_L g661 ( .A(n_334), .B(n_631), .Y(n_661) );
INVx1_ASAP7_75t_L g819 ( .A(n_334), .Y(n_819) );
BUFx3_ASAP7_75t_L g882 ( .A(n_334), .Y(n_882) );
BUFx4f_ASAP7_75t_L g903 ( .A(n_334), .Y(n_903) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_335), .Y(n_532) );
INVx4_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g633 ( .A(n_338), .Y(n_633) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g508 ( .A(n_339), .Y(n_508) );
INVx2_ASAP7_75t_L g739 ( .A(n_339), .Y(n_739) );
INVx2_ASAP7_75t_L g816 ( .A(n_339), .Y(n_816) );
INVx2_ASAP7_75t_SL g995 ( .A(n_339), .Y(n_995) );
INVx1_ASAP7_75t_L g1053 ( .A(n_339), .Y(n_1053) );
BUFx4f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g886 ( .A(n_342), .Y(n_886) );
AOI33xp33_ASAP7_75t_L g808 ( .A1(n_344), .A2(n_809), .A3(n_811), .B1(n_814), .B2(n_817), .B3(n_820), .Y(n_808) );
NAND3xp33_ASAP7_75t_L g1051 ( .A(n_344), .B(n_1052), .C(n_1054), .Y(n_1051) );
AOI33xp33_ASAP7_75t_L g1063 ( .A1(n_344), .A2(n_809), .A3(n_1064), .B1(n_1066), .B2(n_1067), .B3(n_1070), .Y(n_1063) );
AOI33xp33_ASAP7_75t_L g1130 ( .A1(n_344), .A2(n_1048), .A3(n_1131), .B1(n_1132), .B2(n_1134), .B3(n_1135), .Y(n_1130) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
AND2x4_ASAP7_75t_L g355 ( .A(n_345), .B(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g556 ( .A(n_345), .B(n_346), .Y(n_556) );
OR2x6_ASAP7_75t_L g754 ( .A(n_345), .B(n_755), .Y(n_754) );
OR2x2_ASAP7_75t_L g1460 ( .A(n_345), .B(n_755), .Y(n_1460) );
INVx2_ASAP7_75t_L g637 ( .A(n_346), .Y(n_637) );
INVx2_ASAP7_75t_SL g724 ( .A(n_346), .Y(n_724) );
CKINVDCx5p33_ASAP7_75t_R g996 ( .A(n_346), .Y(n_996) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_350), .Y(n_547) );
BUFx2_ASAP7_75t_SL g735 ( .A(n_350), .Y(n_735) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_351), .B(n_1076), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g1108 ( .A(n_354), .Y(n_1108) );
OR2x6_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx2_ASAP7_75t_L g675 ( .A(n_355), .Y(n_675) );
NOR2xp67_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx2_ASAP7_75t_L g626 ( .A(n_358), .Y(n_626) );
INVx1_ASAP7_75t_L g457 ( .A(n_359), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
AND2x2_ASAP7_75t_L g405 ( .A(n_360), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x6_ASAP7_75t_L g409 ( .A(n_361), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g439 ( .A(n_361), .B(n_440), .Y(n_439) );
OR2x6_ASAP7_75t_L g497 ( .A(n_361), .B(n_440), .Y(n_497) );
INVx1_ASAP7_75t_L g1096 ( .A(n_361), .Y(n_1096) );
INVx1_ASAP7_75t_L g1120 ( .A(n_361), .Y(n_1120) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g794 ( .A(n_364), .Y(n_794) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g494 ( .A(n_365), .Y(n_494) );
INVx2_ASAP7_75t_SL g578 ( .A(n_365), .Y(n_578) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_366), .Y(n_398) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx2_ASAP7_75t_L g380 ( .A(n_367), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_367), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g407 ( .A(n_367), .Y(n_407) );
INVx1_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_367), .B(n_368), .Y(n_425) );
INVx1_ASAP7_75t_L g446 ( .A(n_367), .Y(n_446) );
INVx1_ASAP7_75t_L g379 ( .A(n_368), .Y(n_379) );
INVx2_ASAP7_75t_L g386 ( .A(n_368), .Y(n_386) );
AND2x4_ASAP7_75t_L g392 ( .A(n_368), .B(n_380), .Y(n_392) );
INVx1_ASAP7_75t_L g419 ( .A(n_368), .Y(n_419) );
OAI31xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_411), .A3(n_441), .B(n_449), .Y(n_369) );
INVx8_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_372), .A2(n_413), .B1(n_456), .B2(n_457), .C1(n_458), .C2(n_459), .Y(n_455) );
AOI221xp5_ASAP7_75t_SL g1110 ( .A1(n_372), .A2(n_1111), .B1(n_1114), .B2(n_1117), .C(n_1118), .Y(n_1110) );
AND2x4_ASAP7_75t_L g372 ( .A(n_373), .B(n_377), .Y(n_372) );
AND2x4_ASAP7_75t_L g448 ( .A(n_373), .B(n_390), .Y(n_448) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g413 ( .A(n_375), .B(n_398), .Y(n_413) );
AND2x2_ASAP7_75t_L g443 ( .A(n_375), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g402 ( .A(n_376), .Y(n_402) );
INVx1_ASAP7_75t_L g473 ( .A(n_376), .Y(n_473) );
INVx1_ASAP7_75t_L g395 ( .A(n_377), .Y(n_395) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx3_ASAP7_75t_L g574 ( .A(n_378), .Y(n_574) );
AND2x4_ASAP7_75t_L g765 ( .A(n_378), .B(n_766), .Y(n_765) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_378), .Y(n_780) );
BUFx6f_ASAP7_75t_L g806 ( .A(n_378), .Y(n_806) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_378), .Y(n_1031) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
BUFx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g435 ( .A(n_384), .Y(n_435) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g476 ( .A(n_385), .Y(n_476) );
INVx1_ASAP7_75t_L g609 ( .A(n_385), .Y(n_609) );
INVx1_ASAP7_75t_L g410 ( .A(n_386), .Y(n_410) );
AND2x4_ASAP7_75t_L g444 ( .A(n_386), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g1128 ( .A(n_391), .Y(n_1128) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g438 ( .A(n_392), .Y(n_438) );
INVx3_ASAP7_75t_L g480 ( .A(n_392), .Y(n_480) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_392), .Y(n_489) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g1116 ( .A(n_395), .Y(n_1116) );
A2O1A1Ixp33_ASAP7_75t_L g1092 ( .A1(n_396), .A2(n_1093), .B(n_1094), .C(n_1096), .Y(n_1092) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_398), .Y(n_471) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_398), .Y(n_1115) );
INVx2_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g495 ( .A(n_401), .Y(n_495) );
NAND2x1p5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g767 ( .A(n_402), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_405), .A2(n_408), .B1(n_483), .B2(n_484), .Y(n_482) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g587 ( .A(n_407), .Y(n_587) );
AND2x4_ASAP7_75t_L g784 ( .A(n_407), .B(n_772), .Y(n_784) );
CKINVDCx11_ASAP7_75t_R g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g592 ( .A(n_410), .Y(n_592) );
CKINVDCx6p67_ASAP7_75t_R g412 ( .A(n_413), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g1082 ( .A1(n_413), .A2(n_1083), .B1(n_1085), .B2(n_1086), .Y(n_1082) );
AOI221xp5_ASAP7_75t_L g1124 ( .A1(n_413), .A2(n_496), .B1(n_1125), .B2(n_1126), .C(n_1127), .Y(n_1124) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_420), .B1(n_421), .B2(n_426), .C(n_427), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g961 ( .A1(n_415), .A2(n_962), .B1(n_964), .B2(n_965), .Y(n_961) );
OAI22xp33_ASAP7_75t_L g978 ( .A1(n_415), .A2(n_979), .B1(n_980), .B2(n_981), .Y(n_978) );
OAI22xp33_ASAP7_75t_L g1415 ( .A1(n_415), .A2(n_979), .B1(n_1388), .B2(n_1390), .Y(n_1415) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g440 ( .A(n_417), .Y(n_440) );
INVx2_ASAP7_75t_L g492 ( .A(n_417), .Y(n_492) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_418), .B(n_419), .Y(n_469) );
INVx1_ASAP7_75t_L g788 ( .A(n_419), .Y(n_788) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g979 ( .A(n_423), .Y(n_979) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g600 ( .A(n_424), .Y(n_600) );
OR2x2_ASAP7_75t_L g674 ( .A(n_424), .B(n_589), .Y(n_674) );
INVx2_ASAP7_75t_SL g694 ( .A(n_424), .Y(n_694) );
OR2x6_ASAP7_75t_L g771 ( .A(n_424), .B(n_772), .Y(n_771) );
OR2x6_ASAP7_75t_L g775 ( .A(n_424), .B(n_760), .Y(n_775) );
INVx2_ASAP7_75t_SL g963 ( .A(n_424), .Y(n_963) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_430), .Y(n_755) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g472 ( .A(n_431), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_SL g772 ( .A(n_432), .Y(n_772) );
OR2x2_ASAP7_75t_L g861 ( .A(n_432), .B(n_788), .Y(n_861) );
OR2x2_ASAP7_75t_L g913 ( .A(n_432), .B(n_788), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_436), .B2(n_437), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_435), .A2(n_800), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
INVx1_ASAP7_75t_L g612 ( .A(n_437), .Y(n_612) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g763 ( .A(n_438), .Y(n_763) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_440), .Y(n_696) );
INVx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_443), .A2(n_448), .B1(n_461), .B2(n_462), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_443), .A2(n_448), .B1(n_1080), .B2(n_1081), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_443), .A2(n_448), .B1(n_1122), .B2(n_1123), .Y(n_1121) );
BUFx2_ASAP7_75t_L g486 ( .A(n_444), .Y(n_486) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_444), .Y(n_581) );
AND2x4_ASAP7_75t_L g759 ( .A(n_444), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g798 ( .A(n_444), .Y(n_798) );
BUFx2_ASAP7_75t_L g872 ( .A(n_444), .Y(n_872) );
BUFx6f_ASAP7_75t_L g1084 ( .A(n_444), .Y(n_1084) );
BUFx6f_ASAP7_75t_L g1112 ( .A(n_444), .Y(n_1112) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI31xp33_ASAP7_75t_L g984 ( .A1(n_449), .A2(n_985), .A3(n_997), .B(n_1003), .Y(n_984) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
CKINVDCx8_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
AOI221x1_ASAP7_75t_SL g453 ( .A1(n_451), .A2(n_454), .B1(n_498), .B2(n_502), .C(n_533), .Y(n_453) );
INVx2_ASAP7_75t_SL g560 ( .A(n_452), .Y(n_560) );
INVx1_ASAP7_75t_L g558 ( .A(n_453), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_460), .C(n_463), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_456), .A2(n_514), .B1(n_517), .B2(n_518), .Y(n_513) );
OAI221xp5_ASAP7_75t_L g548 ( .A1(n_458), .A2(n_459), .B1(n_536), .B2(n_549), .C(n_552), .Y(n_548) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_485), .C(n_496), .Y(n_463) );
OAI21xp5_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_474), .B(n_482), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_470), .Y(n_465) );
BUFx3_ASAP7_75t_L g602 ( .A(n_467), .Y(n_602) );
BUFx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g714 ( .A(n_468), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_468), .B(n_1095), .Y(n_1094) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g933 ( .A(n_471), .Y(n_933) );
INVx1_ASAP7_75t_L g760 ( .A(n_473), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_477), .B1(n_478), .B2(n_481), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_475), .A2(n_706), .B1(n_707), .B2(n_710), .Y(n_705) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g570 ( .A(n_479), .B(n_571), .Y(n_570) );
BUFx3_ASAP7_75t_L g1414 ( .A(n_479), .Y(n_1414) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g704 ( .A(n_480), .Y(n_704) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_480), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g534 ( .A1(n_481), .A2(n_535), .B1(n_539), .B2(n_540), .C(n_543), .Y(n_534) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_483), .A2(n_484), .B1(n_491), .B2(n_521), .C1(n_523), .C2(n_527), .Y(n_520) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_SL g926 ( .A(n_488), .Y(n_926) );
INVx4_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g615 ( .A(n_489), .Y(n_615) );
BUFx3_ASAP7_75t_L g930 ( .A(n_489), .Y(n_930) );
OAI21xp5_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_492), .B(n_493), .Y(n_490) );
OAI22xp33_ASAP7_75t_L g617 ( .A1(n_492), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g1405 ( .A1(n_492), .A2(n_979), .B1(n_1406), .B2(n_1407), .Y(n_1405) );
BUFx3_ASAP7_75t_L g876 ( .A(n_494), .Y(n_876) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI211x1_ASAP7_75t_L g893 ( .A1(n_498), .A2(n_894), .B(n_908), .C(n_919), .Y(n_893) );
AOI221x1_ASAP7_75t_L g1009 ( .A1(n_498), .A2(n_753), .B1(n_1010), .B2(n_1021), .C(n_1034), .Y(n_1009) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AOI211x1_ASAP7_75t_SL g1426 ( .A1(n_499), .A2(n_1427), .B(n_1439), .C(n_1450), .Y(n_1426) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
AND2x4_ASAP7_75t_L g837 ( .A(n_500), .B(n_501), .Y(n_837) );
INVx2_ASAP7_75t_L g1098 ( .A(n_501), .Y(n_1098) );
NAND4xp25_ASAP7_75t_SL g502 ( .A(n_503), .B(n_513), .C(n_520), .D(n_528), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B1(n_509), .B2(n_510), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_505), .A2(n_510), .B1(n_896), .B2(n_897), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_505), .A2(n_518), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_505), .A2(n_510), .B1(n_1437), .B2(n_1438), .Y(n_1436) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
AND2x6_ASAP7_75t_L g518 ( .A(n_506), .B(n_519), .Y(n_518) );
AND2x4_ASAP7_75t_L g832 ( .A(n_506), .B(n_508), .Y(n_832) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g827 ( .A(n_507), .B(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_510), .A2(n_518), .B1(n_834), .B2(n_835), .Y(n_833) );
CKINVDCx6p67_ASAP7_75t_R g851 ( .A(n_510), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g1014 ( .A1(n_510), .A2(n_514), .B1(n_1015), .B2(n_1016), .C(n_1017), .Y(n_1014) );
INVx1_ASAP7_75t_L g531 ( .A(n_511), .Y(n_531) );
AND2x2_ASAP7_75t_L g824 ( .A(n_511), .B(n_635), .Y(n_824) );
INVx1_ASAP7_75t_L g855 ( .A(n_511), .Y(n_855) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_514), .A2(n_773), .B1(n_831), .B2(n_832), .Y(n_830) );
INVx4_ASAP7_75t_L g856 ( .A(n_514), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_514), .A2(n_518), .B1(n_899), .B2(n_900), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_514), .A2(n_518), .B1(n_1429), .B2(n_1430), .Y(n_1428) );
AND2x4_ASAP7_75t_L g524 ( .A(n_515), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx4_ASAP7_75t_L g852 ( .A(n_518), .Y(n_852) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_519), .Y(n_659) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_519), .Y(n_813) );
INVx2_ASAP7_75t_L g937 ( .A(n_519), .Y(n_937) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AOI222xp33_ASAP7_75t_L g1431 ( .A1(n_523), .A2(n_527), .B1(n_1432), .B2(n_1433), .C1(n_1434), .C2(n_1435), .Y(n_1431) );
BUFx4f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_524), .A2(n_527), .B1(n_847), .B2(n_848), .Y(n_846) );
INVx1_ASAP7_75t_L g906 ( .A(n_524), .Y(n_906) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g828 ( .A(n_526), .Y(n_828) );
INVx3_ASAP7_75t_L g829 ( .A(n_527), .Y(n_829) );
AOI222xp33_ASAP7_75t_L g901 ( .A1(n_527), .A2(n_902), .B1(n_903), .B2(n_904), .C1(n_905), .C2(n_907), .Y(n_901) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND4xp25_ASAP7_75t_SL g894 ( .A(n_529), .B(n_895), .C(n_898), .D(n_901), .Y(n_894) );
NAND4xp25_ASAP7_75t_L g1427 ( .A(n_529), .B(n_1428), .C(n_1431), .D(n_1436), .Y(n_1427) );
INVx5_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI211xp5_ASAP7_75t_L g822 ( .A1(n_530), .A2(n_823), .B(n_824), .C(n_825), .Y(n_822) );
CKINVDCx8_ASAP7_75t_R g849 ( .A(n_530), .Y(n_849) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
OAI21xp33_ASAP7_75t_L g1019 ( .A1(n_531), .A2(n_665), .B(n_1020), .Y(n_1019) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_532), .Y(n_635) );
INVx1_ASAP7_75t_L g653 ( .A(n_532), .Y(n_653) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_532), .Y(n_665) );
INVx2_ASAP7_75t_L g1047 ( .A(n_532), .Y(n_1047) );
BUFx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g854 ( .A(n_538), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g553 ( .A(n_542), .Y(n_553) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_555), .Y(n_554) );
BUFx4f_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AOI33xp33_ASAP7_75t_L g877 ( .A1(n_556), .A2(n_878), .A3(n_879), .B1(n_881), .B2(n_883), .B3(n_885), .Y(n_877) );
BUFx4f_ASAP7_75t_L g942 ( .A(n_556), .Y(n_942) );
AOI33xp33_ASAP7_75t_L g1445 ( .A1(n_556), .A2(n_878), .A3(n_1446), .B1(n_1447), .B2(n_1448), .B3(n_1449), .Y(n_1445) );
INVx1_ASAP7_75t_L g744 ( .A(n_561), .Y(n_744) );
AO22x2_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_676), .B2(n_742), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_624), .Y(n_564) );
NOR3xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_582), .C(n_595), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_575), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_572), .B2(n_573), .Y(n_567) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx2_ASAP7_75t_L g682 ( .A(n_570), .Y(n_682) );
BUFx2_ASAP7_75t_L g950 ( .A(n_570), .Y(n_950) );
BUFx2_ASAP7_75t_L g1397 ( .A(n_570), .Y(n_1397) );
AND2x6_ASAP7_75t_L g573 ( .A(n_571), .B(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g577 ( .A(n_571), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g580 ( .A(n_571), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g955 ( .A(n_571), .B(n_581), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_573), .A2(n_681), .B1(n_682), .B2(n_683), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_573), .A2(n_949), .B1(n_950), .B2(n_951), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1395 ( .A1(n_573), .A2(n_1396), .B1(n_1397), .B2(n_1398), .Y(n_1395) );
NAND2x1p5_ASAP7_75t_L g594 ( .A(n_574), .B(n_588), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B1(n_579), .B2(n_580), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_577), .A2(n_580), .B1(n_685), .B2(n_686), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_577), .A2(n_953), .B1(n_954), .B2(n_955), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_577), .A2(n_580), .B1(n_1400), .B2(n_1401), .Y(n_1399) );
INVx2_ASAP7_75t_SL g929 ( .A(n_581), .Y(n_929) );
INVx2_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2x1_ASAP7_75t_SL g585 ( .A(n_586), .B(n_588), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g1095 ( .A1(n_586), .A2(n_787), .B1(n_1073), .B2(n_1074), .Y(n_1095) );
NAND2x1p5_ASAP7_75t_L g1119 ( .A(n_586), .B(n_1120), .Y(n_1119) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g591 ( .A(n_588), .B(n_592), .Y(n_591) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx4f_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx4f_ASAP7_75t_L g688 ( .A(n_591), .Y(n_688) );
BUFx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx2_ASAP7_75t_L g957 ( .A(n_594), .Y(n_957) );
BUFx3_ASAP7_75t_L g1403 ( .A(n_594), .Y(n_1403) );
OAI33xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .A3(n_603), .B1(n_613), .B2(n_617), .B3(n_621), .Y(n_595) );
OAI33xp33_ASAP7_75t_L g689 ( .A1(n_596), .A2(n_621), .A3(n_690), .B1(n_697), .B2(n_705), .B3(n_711), .Y(n_689) );
INVx1_ASAP7_75t_L g960 ( .A(n_596), .Y(n_960) );
OAI33xp33_ASAP7_75t_L g1404 ( .A1(n_596), .A2(n_621), .A3(n_1405), .B1(n_1408), .B2(n_1412), .B3(n_1415), .Y(n_1404) );
OAI22xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_601), .B2(n_602), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g618 ( .A(n_600), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_610), .B2(n_611), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_605), .A2(n_614), .B1(n_615), .B2(n_616), .Y(n_613) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g699 ( .A(n_608), .Y(n_699) );
BUFx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g970 ( .A(n_609), .Y(n_970) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_614), .A2(n_629), .B1(n_632), .B2(n_638), .C(n_642), .Y(n_628) );
OAI22xp5_ASAP7_75t_SL g1408 ( .A1(n_615), .A2(n_1409), .B1(n_1410), .B2(n_1411), .Y(n_1408) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_616), .A2(n_619), .B1(n_667), .B2(n_669), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_620), .A2(n_649), .B1(n_657), .B2(n_660), .C(n_662), .Y(n_648) );
OAI33xp33_ASAP7_75t_L g958 ( .A1(n_621), .A2(n_959), .A3(n_961), .B1(n_966), .B2(n_974), .B3(n_978), .Y(n_958) );
CKINVDCx8_ASAP7_75t_R g621 ( .A(n_622), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g1039 ( .A(n_622), .B(n_1040), .C(n_1042), .Y(n_1039) );
INVx5_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx6_ASAP7_75t_L g807 ( .A(n_623), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B1(n_671), .B2(n_672), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_625), .A2(n_672), .B1(n_717), .B2(n_741), .Y(n_716) );
AOI31xp33_ASAP7_75t_L g1109 ( .A1(n_625), .A2(n_1110), .A3(n_1121), .B(n_1124), .Y(n_1109) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_648), .C(n_666), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_629), .A2(n_706), .B1(n_719), .B2(n_725), .C(n_729), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g985 ( .A1(n_629), .A2(n_975), .B(n_986), .Y(n_985) );
AOI221xp5_ASAP7_75t_L g1374 ( .A1(n_629), .A2(n_1375), .B1(n_1376), .B2(n_1377), .C(n_1378), .Y(n_1374) );
AND2x4_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
BUFx3_ASAP7_75t_L g639 ( .A(n_630), .Y(n_639) );
INVx1_ASAP7_75t_L g727 ( .A(n_630), .Y(n_727) );
INVx2_ASAP7_75t_SL g734 ( .A(n_630), .Y(n_734) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
HB1xp67_ASAP7_75t_L g1433 ( .A(n_635), .Y(n_1433) );
BUFx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_SL g1379 ( .A(n_644), .Y(n_1379) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
BUFx3_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g1076 ( .A(n_653), .Y(n_1076) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_660), .A2(n_662), .B1(n_715), .B2(n_732), .C(n_737), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_660), .A2(n_662), .B1(n_981), .B2(n_998), .C(n_1001), .Y(n_997) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g1382 ( .A1(n_661), .A2(n_662), .B1(n_1383), .B2(n_1387), .C(n_1388), .Y(n_1382) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g721 ( .A(n_665), .Y(n_721) );
BUFx6f_ASAP7_75t_L g884 ( .A(n_665), .Y(n_884) );
INVx1_ASAP7_75t_L g1385 ( .A(n_665), .Y(n_1385) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_667), .A2(n_669), .B1(n_710), .B2(n_712), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_667), .A2(n_669), .B1(n_977), .B2(n_980), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_667), .A2(n_669), .B1(n_1390), .B2(n_1391), .Y(n_1389) );
INVx6_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx4_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI21xp33_ASAP7_75t_L g982 ( .A1(n_672), .A2(n_983), .B(n_984), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1371 ( .A1(n_672), .A2(n_1372), .B1(n_1373), .B2(n_1392), .Y(n_1371) );
INVx5_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g742 ( .A(n_676), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_716), .Y(n_677) );
NOR3xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_687), .C(n_689), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_684), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B1(n_695), .B2(n_696), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_692), .A2(n_712), .B1(n_713), .B2(n_715), .Y(n_711) );
BUFx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g800 ( .A(n_704), .Y(n_800) );
INVx2_ASAP7_75t_L g803 ( .A(n_704), .Y(n_803) );
HB1xp67_ASAP7_75t_L g1113 ( .A(n_704), .Y(n_1113) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g973 ( .A(n_709), .Y(n_973) );
INVx2_ASAP7_75t_L g1041 ( .A(n_709), .Y(n_1041) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_731), .C(n_740), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g880 ( .A(n_734), .Y(n_880) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
BUFx3_ASAP7_75t_L g939 ( .A(n_739), .Y(n_939) );
XNOR2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_1005), .Y(n_745) );
OA22x2_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_890), .B1(n_891), .B2(n_1004), .Y(n_746) );
INVx1_ASAP7_75t_L g1004 ( .A(n_747), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B1(n_838), .B2(n_889), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
XNOR2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
AOI211xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_756), .B(n_790), .C(n_821), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
AO21x1_ASAP7_75t_SL g857 ( .A1(n_754), .A2(n_858), .B(n_863), .Y(n_857) );
AOI31xp33_ASAP7_75t_L g908 ( .A1(n_754), .A2(n_909), .A3(n_914), .B(n_917), .Y(n_908) );
INVxp67_ASAP7_75t_L g1157 ( .A(n_755), .Y(n_1157) );
NAND4xp25_ASAP7_75t_SL g756 ( .A(n_757), .B(n_764), .C(n_768), .D(n_776), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .B1(n_761), .B2(n_762), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_759), .A2(n_864), .B1(n_865), .B2(n_866), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_759), .A2(n_762), .B1(n_915), .B2(n_916), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_759), .A2(n_762), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1454 ( .A1(n_759), .A2(n_866), .B1(n_1455), .B2(n_1456), .Y(n_1454) );
AND2x4_ASAP7_75t_L g762 ( .A(n_760), .B(n_763), .Y(n_762) );
AND2x4_ASAP7_75t_L g866 ( .A(n_760), .B(n_763), .Y(n_866) );
NAND4xp25_ASAP7_75t_SL g1021 ( .A(n_764), .B(n_1022), .C(n_1025), .D(n_1032), .Y(n_1021) );
CKINVDCx11_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
NOR3xp33_ASAP7_75t_L g858 ( .A(n_765), .B(n_859), .C(n_862), .Y(n_858) );
AOI211xp5_ASAP7_75t_L g909 ( .A1(n_765), .A2(n_869), .B(n_910), .C(n_911), .Y(n_909) );
AOI211xp5_ASAP7_75t_L g1451 ( .A1(n_765), .A2(n_1116), .B(n_1452), .C(n_1453), .Y(n_1451) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVxp67_ASAP7_75t_L g789 ( .A(n_767), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B1(n_773), .B2(n_774), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_770), .A2(n_774), .B1(n_899), .B2(n_918), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_770), .A2(n_774), .B1(n_1015), .B2(n_1033), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_770), .A2(n_1429), .B1(n_1458), .B2(n_1459), .Y(n_1457) );
INVx8_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g1156 ( .A(n_771), .B(n_1157), .Y(n_1156) );
INVx4_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx5_ASAP7_75t_L g1459 ( .A(n_775), .Y(n_1459) );
AOI222xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B1(n_781), .B2(n_782), .C1(n_785), .C2(n_786), .Y(n_776) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_SL g924 ( .A(n_779), .Y(n_924) );
INVx2_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_780), .Y(n_795) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g860 ( .A(n_784), .Y(n_860) );
INVx2_ASAP7_75t_L g912 ( .A(n_784), .Y(n_912) );
AOI222xp33_ASAP7_75t_L g1025 ( .A1(n_784), .A2(n_786), .B1(n_1026), .B2(n_1027), .C1(n_1028), .C2(n_1029), .Y(n_1025) );
AND2x4_ASAP7_75t_L g786 ( .A(n_787), .B(n_789), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g790 ( .A(n_791), .B(n_808), .Y(n_790) );
AOI33xp33_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .A3(n_796), .B1(n_801), .B2(n_804), .B3(n_807), .Y(n_791) );
AOI33xp33_ASAP7_75t_L g867 ( .A1(n_792), .A2(n_807), .A3(n_868), .B1(n_871), .B2(n_874), .B3(n_875), .Y(n_867) );
NAND3xp33_ASAP7_75t_L g1035 ( .A(n_792), .B(n_1036), .C(n_1038), .Y(n_1035) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g873 ( .A(n_800), .Y(n_873) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx2_ASAP7_75t_SL g1037 ( .A(n_803), .Y(n_1037) );
BUFx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_SL g870 ( .A(n_806), .Y(n_870) );
AOI33xp33_ASAP7_75t_L g920 ( .A1(n_807), .A2(n_921), .A3(n_923), .B1(n_925), .B2(n_927), .B3(n_931), .Y(n_920) );
AOI33xp33_ASAP7_75t_L g1440 ( .A1(n_807), .A2(n_921), .A3(n_1441), .B1(n_1442), .B2(n_1443), .B3(n_1444), .Y(n_1440) );
INVx1_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
AOI31xp33_ASAP7_75t_SL g821 ( .A1(n_822), .A2(n_830), .A3(n_833), .B(n_836), .Y(n_821) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g1018 ( .A(n_827), .Y(n_1018) );
INVx1_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
OAI31xp33_ASAP7_75t_L g841 ( .A1(n_837), .A2(n_842), .A3(n_850), .B(n_853), .Y(n_841) );
INVx1_ASAP7_75t_L g889 ( .A(n_838), .Y(n_889) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
AND4x1_ASAP7_75t_L g840 ( .A(n_841), .B(n_857), .C(n_867), .D(n_877), .Y(n_840) );
NAND4xp25_ASAP7_75t_L g888 ( .A(n_841), .B(n_857), .C(n_867), .D(n_877), .Y(n_888) );
NAND3xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_846), .C(n_849), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
AOI33xp33_ASAP7_75t_L g934 ( .A1(n_878), .A2(n_935), .A3(n_938), .B1(n_940), .B2(n_941), .B3(n_942), .Y(n_934) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
XNOR2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_943), .Y(n_891) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_934), .Y(n_919) );
BUFx3_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx3_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g976 ( .A(n_930), .Y(n_976) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
XNOR2x1_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
AND2x2_ASAP7_75t_L g945 ( .A(n_946), .B(n_982), .Y(n_945) );
NOR3xp33_ASAP7_75t_SL g946 ( .A(n_947), .B(n_956), .C(n_958), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_948), .B(n_952), .Y(n_947) );
OAI211xp5_ASAP7_75t_L g989 ( .A1(n_951), .A2(n_990), .B(n_992), .C(n_994), .Y(n_989) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx3_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_967), .A2(n_968), .B1(n_971), .B2(n_972), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_968), .A2(n_975), .B1(n_976), .B2(n_977), .Y(n_974) );
INVx2_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx2_ASAP7_75t_L g1410 ( .A(n_969), .Y(n_1410) );
INVx2_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx1_ASAP7_75t_SL g987 ( .A(n_988), .Y(n_987) );
INVx2_ASAP7_75t_SL g990 ( .A(n_991), .Y(n_990) );
BUFx6f_ASAP7_75t_L g1002 ( .A(n_993), .Y(n_1002) );
INVx1_ASAP7_75t_L g1069 ( .A(n_995), .Y(n_1069) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
INVx3_ASAP7_75t_L g1386 ( .A(n_1000), .Y(n_1386) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_1006), .A2(n_1104), .B1(n_1146), .B2(n_1147), .Y(n_1005) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1006), .Y(n_1146) );
XOR2xp5_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1057), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1009), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1014), .Y(n_1010) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
NAND4xp25_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1039), .C(n_1043), .D(n_1051), .Y(n_1034) );
NAND3xp33_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .C(n_1048), .Y(n_1043) );
INVx3_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
INVx2_ASAP7_75t_L g1133 ( .A(n_1047), .Y(n_1133) );
INVx3_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx2_ASAP7_75t_SL g1058 ( .A(n_1059), .Y(n_1058) );
INVx2_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
NAND4xp75_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1077), .C(n_1099), .D(n_1101), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1071), .Y(n_1062) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
OAI21xp5_ASAP7_75t_L g1077 ( .A1(n_1078), .A2(n_1087), .B(n_1097), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1082), .Y(n_1078) );
BUFx8_ASAP7_75t_SL g1097 ( .A(n_1098), .Y(n_1097) );
INVx2_ASAP7_75t_L g1372 ( .A(n_1098), .Y(n_1372) );
INVx2_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_1105), .Y(n_1147) );
XOR2x2_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1145), .Y(n_1105) );
NOR3xp33_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1109), .C(n_1129), .Y(n_1106) );
NAND4xp25_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1136), .C(n_1139), .D(n_1142), .Y(n_1129) );
BUFx3_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
AND2x4_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1155), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1420 ( .A(n_1150), .B(n_1156), .Y(n_1420) );
NOR2xp33_ASAP7_75t_SL g1150 ( .A(n_1151), .B(n_1153), .Y(n_1150) );
INVx1_ASAP7_75t_SL g1464 ( .A(n_1151), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1151), .B(n_1153), .Y(n_1470) );
HB1xp67_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1153), .B(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
OAI21xp33_ASAP7_75t_L g1158 ( .A1(n_1159), .A2(n_1167), .B(n_1367), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_1161), .A2(n_1221), .B1(n_1222), .B2(n_1223), .Y(n_1220) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1161), .Y(n_1237) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
AND2x4_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1165), .Y(n_1162) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1163), .Y(n_1185) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1164), .B(n_1177), .Y(n_1176) );
AND2x4_ASAP7_75t_L g1184 ( .A(n_1165), .B(n_1185), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1165), .B(n_1185), .Y(n_1191) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1166), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1167 ( .A1(n_1168), .A2(n_1248), .B1(n_1311), .B2(n_1312), .C(n_1340), .Y(n_1167) );
A2O1A1Ixp33_ASAP7_75t_SL g1168 ( .A1(n_1169), .A2(n_1203), .B(n_1230), .C(n_1241), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1186), .Y(n_1169) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1171), .B(n_1261), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1171), .B(n_1228), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1171), .B(n_1269), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1171), .B(n_1321), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1171), .B(n_1290), .Y(n_1355) );
BUFx2_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1207 ( .A(n_1172), .B(n_1208), .Y(n_1207) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1172), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1172), .B(n_1252), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1172), .B(n_1279), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1172), .B(n_1209), .Y(n_1283) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1172), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1172), .B(n_1187), .Y(n_1336) );
AOI211xp5_ASAP7_75t_L g1343 ( .A1(n_1172), .A2(n_1255), .B(n_1344), .C(n_1345), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1172), .B(n_1286), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1183), .Y(n_1172) );
AND2x4_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1178), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1176), .B(n_1179), .Y(n_1200) );
HB1xp67_ASAP7_75t_L g1469 ( .A(n_1177), .Y(n_1469) );
AND2x4_ASAP7_75t_L g1180 ( .A(n_1178), .B(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1179), .B(n_1182), .Y(n_1202) );
BUFx2_ASAP7_75t_L g1235 ( .A(n_1180), .Y(n_1235) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1184), .Y(n_1221) );
BUFx3_ASAP7_75t_L g1242 ( .A(n_1184), .Y(n_1242) );
HB1xp67_ASAP7_75t_L g1467 ( .A(n_1185), .Y(n_1467) );
O2A1O1Ixp33_ASAP7_75t_L g1330 ( .A1(n_1186), .A2(n_1293), .B(n_1331), .C(n_1334), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1192), .Y(n_1186) );
NOR2x1_ASAP7_75t_L g1255 ( .A(n_1187), .B(n_1229), .Y(n_1255) );
AOI21xp5_ASAP7_75t_L g1284 ( .A1(n_1187), .A2(n_1285), .B(n_1288), .Y(n_1284) );
NOR2xp33_ASAP7_75t_L g1290 ( .A(n_1187), .B(n_1193), .Y(n_1290) );
BUFx2_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
BUFx3_ASAP7_75t_L g1208 ( .A(n_1188), .Y(n_1208) );
INVxp67_ASAP7_75t_L g1253 ( .A(n_1188), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1188), .B(n_1297), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1192), .B(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1192), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1197), .Y(n_1192) );
AOI22xp5_ASAP7_75t_L g1313 ( .A1(n_1193), .A2(n_1314), .B1(n_1318), .B2(n_1320), .Y(n_1313) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1194), .B(n_1197), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1194), .B(n_1229), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1194), .B(n_1208), .Y(n_1268) );
OR2x2_ASAP7_75t_L g1298 ( .A(n_1194), .B(n_1197), .Y(n_1298) );
NOR2xp33_ASAP7_75t_L g1362 ( .A(n_1194), .B(n_1208), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1196), .Y(n_1194) );
INVx2_ASAP7_75t_SL g1229 ( .A(n_1197), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1197), .B(n_1208), .Y(n_1279) );
OAI22xp5_ASAP7_75t_L g1198 ( .A1(n_1199), .A2(n_1200), .B1(n_1201), .B2(n_1202), .Y(n_1198) );
BUFx6f_ASAP7_75t_L g1215 ( .A(n_1200), .Y(n_1215) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1202), .Y(n_1218) );
AOI21xp5_ASAP7_75t_L g1203 ( .A1(n_1204), .A2(n_1210), .B(n_1224), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1209), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1207), .B(n_1298), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1208), .B(n_1228), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1208), .B(n_1303), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1208), .B(n_1304), .Y(n_1344) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1209), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1209), .B(n_1336), .Y(n_1335) );
INVx2_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1211), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1276 ( .A1(n_1211), .A2(n_1274), .B1(n_1277), .B2(n_1278), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1211), .B(n_1225), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1211), .B(n_1348), .Y(n_1347) );
INVx2_ASAP7_75t_SL g1211 ( .A(n_1212), .Y(n_1211) );
AND2x4_ASAP7_75t_L g1274 ( .A(n_1212), .B(n_1270), .Y(n_1274) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1212), .Y(n_1281) );
NOR2xp33_ASAP7_75t_L g1295 ( .A(n_1212), .B(n_1296), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1212), .B(n_1265), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1212), .B(n_1238), .Y(n_1321) );
HB1xp67_ASAP7_75t_L g1328 ( .A(n_1212), .Y(n_1328) );
CKINVDCx5p33_ASAP7_75t_R g1212 ( .A(n_1213), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1213), .B(n_1238), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1213), .B(n_1270), .Y(n_1287) );
OR2x2_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1220), .Y(n_1213) );
OAI22xp5_ASAP7_75t_L g1214 ( .A1(n_1215), .A2(n_1216), .B1(n_1217), .B2(n_1219), .Y(n_1214) );
BUFx3_ASAP7_75t_L g1245 ( .A(n_1215), .Y(n_1245) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_1217), .Y(n_1247) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
NOR2xp33_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1226), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1225), .B(n_1268), .Y(n_1267) );
O2A1O1Ixp33_ASAP7_75t_L g1271 ( .A1(n_1225), .A2(n_1229), .B(n_1272), .C(n_1273), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1225), .B(n_1297), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1225), .B(n_1274), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1225), .B(n_1279), .Y(n_1339) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1227), .B(n_1296), .Y(n_1353) );
OAI21xp5_ASAP7_75t_L g1359 ( .A1(n_1227), .A2(n_1287), .B(n_1339), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1228), .B(n_1253), .Y(n_1277) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1228), .Y(n_1316) );
OAI32xp33_ASAP7_75t_L g1262 ( .A1(n_1229), .A2(n_1263), .A3(n_1264), .B1(n_1266), .B2(n_1269), .Y(n_1262) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1238), .Y(n_1231) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1232), .Y(n_1259) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1232), .Y(n_1265) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1233), .Y(n_1286) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1233), .B(n_1238), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1233), .B(n_1270), .Y(n_1333) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1233), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1236), .Y(n_1233) );
INVx3_ASAP7_75t_L g1270 ( .A(n_1238), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1240), .Y(n_1238) );
INVx3_ASAP7_75t_L g1299 ( .A(n_1241), .Y(n_1299) );
OAI21xp5_ASAP7_75t_L g1350 ( .A1(n_1241), .A2(n_1321), .B(n_1351), .Y(n_1350) );
OAI22xp33_ASAP7_75t_L g1243 ( .A1(n_1244), .A2(n_1245), .B1(n_1246), .B2(n_1247), .Y(n_1243) );
NAND5xp2_ASAP7_75t_L g1248 ( .A(n_1249), .B(n_1254), .C(n_1275), .D(n_1284), .E(n_1300), .Y(n_1248) );
OR2x2_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1251), .Y(n_1249) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1252), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1253), .B(n_1283), .Y(n_1282) );
AOI211xp5_ASAP7_75t_L g1254 ( .A1(n_1255), .A2(n_1256), .B(n_1262), .C(n_1271), .Y(n_1254) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
NOR2xp33_ASAP7_75t_L g1366 ( .A(n_1257), .B(n_1302), .Y(n_1366) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1260), .Y(n_1257) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1259), .Y(n_1292) );
O2A1O1Ixp33_ASAP7_75t_L g1346 ( .A1(n_1259), .A2(n_1282), .B(n_1347), .C(n_1349), .Y(n_1346) );
OAI22xp5_ASAP7_75t_SL g1307 ( .A1(n_1260), .A2(n_1308), .B1(n_1309), .B2(n_1310), .Y(n_1307) );
A2O1A1Ixp33_ASAP7_75t_L g1334 ( .A1(n_1260), .A2(n_1335), .B(n_1337), .C(n_1338), .Y(n_1334) );
A2O1A1Ixp33_ASAP7_75t_L g1357 ( .A1(n_1260), .A2(n_1329), .B(n_1358), .C(n_1359), .Y(n_1357) );
CKINVDCx5p33_ASAP7_75t_R g1260 ( .A(n_1261), .Y(n_1260) );
AOI22xp5_ASAP7_75t_L g1275 ( .A1(n_1264), .A2(n_1276), .B1(n_1280), .B2(n_1282), .Y(n_1275) );
OAI211xp5_ASAP7_75t_SL g1312 ( .A1(n_1264), .A2(n_1313), .B(n_1322), .C(n_1330), .Y(n_1312) );
INVx2_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1265), .B(n_1274), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1265), .B(n_1281), .Y(n_1351) );
OAI322xp33_ASAP7_75t_L g1360 ( .A1(n_1266), .A2(n_1273), .A3(n_1309), .B1(n_1310), .B2(n_1361), .C1(n_1363), .C2(n_1365), .Y(n_1360) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1268), .Y(n_1309) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
NAND3xp33_ASAP7_75t_L g1294 ( .A(n_1270), .B(n_1295), .C(n_1297), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1341 ( .A(n_1270), .B(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1277), .Y(n_1324) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1281), .B(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1285), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1287), .Y(n_1285) );
OAI211xp5_ASAP7_75t_L g1288 ( .A1(n_1289), .A2(n_1291), .B(n_1294), .C(n_1299), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1293), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1297), .B(n_1336), .Y(n_1348) );
NOR2xp33_ASAP7_75t_SL g1361 ( .A(n_1297), .B(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1299), .Y(n_1311) );
O2A1O1Ixp33_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1304), .B(n_1305), .C(n_1307), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
OAI21xp5_ASAP7_75t_L g1354 ( .A1(n_1304), .A2(n_1345), .B(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1317), .Y(n_1315) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
O2A1O1Ixp33_ASAP7_75t_L g1322 ( .A1(n_1323), .A2(n_1324), .B(n_1325), .C(n_1327), .Y(n_1322) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1323), .Y(n_1337) );
OAI21xp5_ASAP7_75t_L g1338 ( .A1(n_1324), .A2(n_1333), .B(n_1339), .Y(n_1338) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
NOR2xp33_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1329), .Y(n_1327) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
OAI211xp5_ASAP7_75t_SL g1340 ( .A1(n_1341), .A2(n_1343), .B(n_1346), .C(n_1356), .Y(n_1340) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1348), .Y(n_1358) );
OAI21xp5_ASAP7_75t_L g1349 ( .A1(n_1350), .A2(n_1352), .B(n_1354), .Y(n_1349) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
NOR3xp33_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1360), .C(n_1366), .Y(n_1356) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
BUFx2_ASAP7_75t_SL g1368 ( .A(n_1369), .Y(n_1368) );
XOR2x2_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1416), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1393), .Y(n_1370) );
NAND3xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1382), .C(n_1389), .Y(n_1373) );
OAI22xp5_ASAP7_75t_L g1412 ( .A1(n_1377), .A2(n_1391), .B1(n_1410), .B2(n_1413), .Y(n_1412) );
INVx3_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
NOR3xp33_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1402), .C(n_1404), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1395), .B(n_1399), .Y(n_1394) );
CKINVDCx5p33_ASAP7_75t_R g1413 ( .A(n_1414), .Y(n_1413) );
BUFx2_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
HB1xp67_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1445), .Y(n_1439) );
AOI31xp33_ASAP7_75t_L g1450 ( .A1(n_1451), .A2(n_1454), .A3(n_1457), .B(n_1460), .Y(n_1450) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
CKINVDCx5p33_ASAP7_75t_R g1462 ( .A(n_1463), .Y(n_1462) );
A2O1A1Ixp33_ASAP7_75t_L g1465 ( .A1(n_1464), .A2(n_1466), .B(n_1468), .C(n_1470), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
endmodule